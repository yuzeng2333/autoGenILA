module PID(i_clk, i_rst, i_wb_cyc, i_wb_stb, i_wb_we, i_wb_adr, i_wb_data, o_wb_ack, o_wb_data, o_un, o_valid);
  wire [31:0] _0000_;
  wire _0001_;
  wire [31:0] _0002_;
  wire _0003_;
  wire [15:0] _0004_;
  wire [15:0] _0005_;
  wire [15:0] _0006_;
  wire [15:0] _0007_;
  wire [15:0] _0008_;
  wire [15:0] _0009_;
  wire [1:0] _0010_;
  wire [1:0] _0011_;
  wire [4:0] _0012_;
  wire [31:0] _0013_;
  wire [15:0] _0014_;
  wire _0015_;
  wire _0016_;
  wire [31:0] _0017_;
  wire [15:0] _0018_;
  wire _0019_;
  wire _0020_;
  wire [9:0] _0021_;
  wire [31:0] _0022_;
  wire _0023_;
  wire _0024_;
  wire _0025_;
  wire _0026_;
  wire _0027_;
  wire _0028_;
  wire _0029_;
  wire _0030_;
  wire _0031_;
  wire _0032_;
  wire _0033_;
  wire _0034_;
  wire _0035_;
  wire [31:0] _0036_;
  wire [31:0] _0037_;
  wire _0038_;
  wire _0039_;
  wire _0040_;
  wire _0041_;
  wire _0042_;
  wire _0043_;
  wire _0044_;
  wire _0045_;
  wire _0046_;
  wire _0047_;
  wire _0048_;
  wire _0049_;
  wire _0050_;
  wire _0051_;
  wire _0052_;
  wire _0053_;
  wire _0054_;
  wire _0055_;
  wire _0056_;
  wire _0057_;
  wire _0058_;
  wire _0059_;
  wire _0060_;
  wire _0061_;
  wire _0062_;
  wire _0063_;
  wire _0064_;
  wire _0065_;
  wire _0066_;
  wire _0067_;
  wire _0068_;
  wire _0069_;
  wire _0070_;
  wire _0071_;
  wire _0072_;
  wire [15:0] _0073_;
  wire _0074_;
  wire [15:0] _0075_;
  wire _0076_;
  wire _0077_;
  wire _0078_;
  wire _0079_;
  wire _0080_;
  wire _0081_;
  wire _0082_;
  wire _0083_;
  wire _0084_;
  wire _0085_;
  wire _0086_;
  wire _0087_;
  wire _0088_;
  wire _0089_;
  wire _0090_;
  wire _0091_;
  wire _0092_;
  wire _0093_;
  wire _0094_;
  wire _0095_;
  wire _0096_;
  wire _0097_;
  wire _0098_;
  wire _0099_;
  wire _0100_;
  wire _0101_;
  wire _0102_;
  wire _0103_;
  wire _0104_;
  wire _0105_;
  wire _0106_;
  wire _0107_;
  wire _0108_;
  wire _0109_;
  wire _0110_;
  wire _0111_;
  wire _0112_;
  wire _0113_;
  wire _0114_;
  wire _0115_;
  wire _0116_;
  wire _0117_;
  wire [15:0] _0118_;
  wire [15:0] _0119_;
  wire [15:0] _0120_;
  wire _0121_;
  wire _0122_;
  wire [31:0] _0123_;
  wire [31:0] _0124_;
  wire [31:0] _0125_;
  wire [31:0] _0126_;
  wire [31:0] _0127_;
  wire [31:0] _0128_;
  wire _0129_;
  wire _0130_;
  wire _0131_;
  wire _0132_;
  wire [9:0] _0133_;
  wire [9:0] _0134_;
  wire _0135_;
  wire _0136_;
  wire _0137_;
  wire _0138_;
  wire _0139_;
  wire _0140_;
  wire _0141_;
  wire _0142_;
  wire _0143_;
  wire _0144_;
  wire _0145_;
  wire [15:0] _0146_;
  wire [15:0] _0147_;
  wire [15:0] _0148_;
  wire [15:0] _0149_;
  wire _0150_;
  wire [15:0] _0151_;
  wire [15:0] _0152_;
  wire [15:0] _0153_;
  wire _0154_;
  wire [15:0] _0155_;
  wire [15:0] _0156_;
  wire [15:0] _0157_;
  wire _0158_;
  wire [15:0] _0159_;
  wire [15:0] _0160_;
  wire [15:0] _0161_;
  wire _0162_;
  wire [15:0] _0163_;
  wire [15:0] _0164_;
  wire _0165_;
  wire _0166_;
  wire _0167_;
  wire _0168_;
  wire _0169_;
  wire _0170_;
  wire _0171_;
  wire _0172_;
  wire _0173_;
  wire _0174_;
  wire _0175_;
  wire _0176_;
  wire _0177_;
  wire _0178_;
  wire _0179_;
  wire _0180_;
  wire _0181_;
  wire _0182_;
  wire _0183_;
  wire _0184_;
  wire _0185_;
  wire _0186_;
  wire _0187_;
  wire _0188_;
  wire _0189_;
  wire _0190_;
  wire _0191_;
  wire _0192_;
  wire _0193_;
  wire _0194_;
  wire _0195_;
  wire _0196_;
  wire _0197_;
  wire _0198_;
  wire _0199_;
  wire _0200_;
  wire _0201_;
  wire _0202_;
  wire _0203_;
  wire _0204_;
  wire _0205_;
  wire _0206_;
  wire _0207_;
  wire _0208_;
  wire _0209_;
  wire _0210_;
  wire _0211_;
  wire _0212_;
  wire _0213_;
  wire _0214_;
  wire _0215_;
  wire _0216_;
  wire _0217_;
  wire _0218_;
  wire _0219_;
  wire _0220_;
  wire _0221_;
  wire _0222_;
  wire _0223_;
  wire _0224_;
  wire _0225_;
  wire _0226_;
  wire _0227_;
  wire _0228_;
  wire _0229_;
  wire _0230_;
  wire _0231_;
  wire _0232_;
  wire _0233_;
  wire _0234_;
  wire _0235_;
  wire _0236_;
  wire _0237_;
  wire _0238_;
  wire _0239_;
  wire _0240_;
  wire _0241_;
  wire _0242_;
  wire _0243_;
  wire _0244_;
  wire _0245_;
  wire [15:0] _0246_;
  wire [15:0] _0247_;
  wire [1:0] _0248_;
  wire [1:0] _0249_;
  wire [3:0] _0250_;
  wire [2:0] _0251_;
  wire [2:0] _0252_;
  wire [2:0] _0253_;
  wire [2:0] _0254_;
  wire [3:0] _0255_;
  wire [2:0] _0256_;
  wire [3:0] _0257_;
  wire [2:0] _0258_;
  wire _0259_;
  wire [3:0] _0260_;
  wire [2:0] _0261_;
  wire [1:0] _0262_;
  wire [1:0] _0263_;
  wire [2:0] _0264_;
  wire [1:0] _0265_;
  wire [2:0] _0266_;
  wire [1:0] _0267_;
  wire _0268_;
  wire [2:0] _0269_;
  wire [2:0] _0270_;
  wire _0271_;
  wire _0272_;
  wire [1:0] _0273_;
  wire [1:0] _0274_;
  wire [1:0] _0275_;
  wire [1:0] _0276_;
  wire [1:0] _0277_;
  wire [1:0] _0278_;
  wire [1:0] _0279_;
  wire _0280_;
  wire _0281_;
  wire _0282_;
  wire _0283_;
  wire _0284_;
  wire _0285_;
  wire _0286_;
  wire _0287_;
  wire _0288_;
  wire _0289_;
  wire _0290_;
  wire _0291_;
  wire _0292_;
  wire _0293_;
  wire _0294_;
  wire _0295_;
  wire _0296_;
  wire _0297_;
  wire _0298_;
  wire _0299_;
  wire _0300_;
  wire _0301_;
  wire _0302_;
  wire _0303_;
  wire _0304_;
  wire _0305_;
  wire _0306_;
  wire _0307_;
  wire _0308_;
  wire _0309_;
  wire _0310_;
  wire _0311_;
  wire _0312_;
  wire _0313_;
  wire _0314_;
  wire _0315_;
  wire _0316_;
  wire _0317_;
  wire _0318_;
  wire _0319_;
  wire _0320_;
  wire _0321_;
  wire _0322_;
  wire _0323_;
  wire _0324_;
  wire _0325_;
  wire _0326_;
  wire _0327_;
  wire _0328_;
  wire _0329_;
  wire _0330_;
  wire _0331_;
  wire _0332_;
  wire _0333_;
  wire _0334_;
  wire _0335_;
  wire _0336_;
  wire _0337_;
  wire _0338_;
  wire _0339_;
  wire _0340_;
  wire _0341_;
  wire _0342_;
  wire _0343_;
  wire _0344_;
  wire _0345_;
  wire _0346_;
  wire _0347_;
  wire _0348_;
  wire _0349_;
  wire _0350_;
  wire _0351_;
  wire _0352_;
  wire _0353_;
  wire _0354_;
  wire _0355_;
  wire _0356_;
  wire _0357_;
  wire _0358_;
  wire _0359_;
  wire _0360_;
  wire _0361_;
  wire _0362_;
  wire _0363_;
  wire _0364_;
  wire _0365_;
  wire _0366_;
  wire _0367_;
  wire _0368_;
  wire _0369_;
  wire _0370_;
  wire _0371_;
  wire _0372_;
  wire _0373_;
  wire _0374_;
  wire _0375_;
  wire _0376_;
  wire _0377_;
  wire _0378_;
  wire _0379_;
  wire _0380_;
  wire _0381_;
  wire _0382_;
  wire _0383_;
  wire _0384_;
  wire _0385_;
  wire _0386_;
  wire _0387_;
  wire _0388_;
  wire _0389_;
  wire _0390_;
  wire _0391_;
  wire _0392_;
  wire _0393_;
  wire _0394_;
  wire _0395_;
  wire _0396_;
  wire _0397_;
  wire _0398_;
  wire _0399_;
  wire _0400_;
  wire _0401_;
  wire _0402_;
  wire _0403_;
  wire _0404_;
  wire _0405_;
  wire _0406_;
  wire _0407_;
  wire _0408_;
  wire _0409_;
  wire _0410_;
  wire _0411_;
  wire _0412_;
  wire _0413_;
  wire _0414_;
  wire _0415_;
  wire _0416_;
  wire _0417_;
  wire _0418_;
  wire _0419_;
  wire _0420_;
  wire _0421_;
  wire _0422_;
  wire _0423_;
  wire _0424_;
  wire _0425_;
  wire _0426_;
  wire _0427_;
  wire _0428_;
  wire _0429_;
  wire _0430_;
  wire _0431_;
  wire _0432_;
  wire _0433_;
  wire _0434_;
  wire _0435_;
  wire _0436_;
  wire _0437_;
  wire _0438_;
  wire _0439_;
  wire _0440_;
  wire _0441_;
  wire _0442_;
  wire _0443_;
  wire _0444_;
  wire _0445_;
  wire _0446_;
  wire _0447_;
  wire _0448_;
  wire _0449_;
  wire _0450_;
  wire _0451_;
  wire _0452_;
  wire _0453_;
  wire _0454_;
  wire _0455_;
  wire _0456_;
  wire _0457_;
  wire _0458_;
  wire _0459_;
  wire _0460_;
  wire _0461_;
  wire _0462_;
  wire _0463_;
  wire _0464_;
  wire _0465_;
  wire _0466_;
  wire _0467_;
  wire _0468_;
  wire _0469_;
  wire _0470_;
  wire _0471_;
  wire _0472_;
  wire _0473_;
  wire _0474_;
  wire _0475_;
  wire _0476_;
  wire _0477_;
  wire _0478_;
  wire _0479_;
  wire _0480_;
  wire _0481_;
  wire _0482_;
  wire _0483_;
  wire _0484_;
  wire _0485_;
  wire _0486_;
  wire _0487_;
  wire _0488_;
  wire _0489_;
  wire _0490_;
  wire _0491_;
  wire _0492_;
  wire _0493_;
  wire _0494_;
  wire _0495_;
  wire _0496_;
  wire _0497_;
  wire _0498_;
  wire _0499_;
  wire _0500_;
  wire _0501_;
  wire _0502_;
  wire _0503_;
  wire _0504_;
  wire _0505_;
  wire _0506_;
  wire _0507_;
  wire _0508_;
  wire _0509_;
  wire _0510_;
  wire _0511_;
  wire _0512_;
  wire _0513_;
  wire _0514_;
  wire _0515_;
  wire _0516_;
  wire [15:0] _0517_;
  wire [15:0] _0518_;
  wire [15:0] _0519_;
  reg RS;
  reg [31:0] a;
  wire [31:0] \adder_32bit_0.G0 ;
  wire [15:0] \adder_32bit_0.G1 ;
  wire [15:0] \adder_32bit_0.G2 ;
  wire [15:0] \adder_32bit_0.G3 ;
  wire [15:0] \adder_32bit_0.G4 ;
  wire [15:0] \adder_32bit_0.G5 ;
  wire [31:0] \adder_32bit_0.G6 ;
  wire [31:0] \adder_32bit_0.P0 ;
  wire [15:1] \adder_32bit_0.P1 ;
  wire [15:2] \adder_32bit_0.P2 ;
  wire [15:4] \adder_32bit_0.P3 ;
  wire [15:8] \adder_32bit_0.P4 ;
  wire [31:0] \adder_32bit_0.i_a ;
  wire [31:0] \adder_32bit_0.i_b ;
  wire \adder_32bit_0.i_c ;
  wire [31:0] \adder_32bit_0.o_s ;
  wire \adder_32bit_0.operator_A_0.A ;
  wire \adder_32bit_0.operator_A_0.B ;
  wire \adder_32bit_0.operator_A_0.G ;
  wire \adder_32bit_0.operator_A_0.P ;
  wire \adder_32bit_0.operator_A_1.A ;
  wire \adder_32bit_0.operator_A_1.B ;
  wire \adder_32bit_0.operator_A_1.G ;
  wire \adder_32bit_0.operator_A_1.P ;
  wire \adder_32bit_0.operator_A_10.A ;
  wire \adder_32bit_0.operator_A_10.B ;
  wire \adder_32bit_0.operator_A_10.G ;
  wire \adder_32bit_0.operator_A_10.P ;
  wire \adder_32bit_0.operator_A_11.A ;
  wire \adder_32bit_0.operator_A_11.B ;
  wire \adder_32bit_0.operator_A_11.G ;
  wire \adder_32bit_0.operator_A_11.P ;
  wire \adder_32bit_0.operator_A_12.A ;
  wire \adder_32bit_0.operator_A_12.B ;
  wire \adder_32bit_0.operator_A_12.G ;
  wire \adder_32bit_0.operator_A_12.P ;
  wire \adder_32bit_0.operator_A_13.A ;
  wire \adder_32bit_0.operator_A_13.B ;
  wire \adder_32bit_0.operator_A_13.G ;
  wire \adder_32bit_0.operator_A_13.P ;
  wire \adder_32bit_0.operator_A_14.A ;
  wire \adder_32bit_0.operator_A_14.B ;
  wire \adder_32bit_0.operator_A_14.G ;
  wire \adder_32bit_0.operator_A_14.P ;
  wire \adder_32bit_0.operator_A_15.A ;
  wire \adder_32bit_0.operator_A_15.B ;
  wire \adder_32bit_0.operator_A_15.G ;
  wire \adder_32bit_0.operator_A_15.P ;
  wire \adder_32bit_0.operator_A_16.A ;
  wire \adder_32bit_0.operator_A_16.B ;
  wire \adder_32bit_0.operator_A_16.G ;
  wire \adder_32bit_0.operator_A_16.P ;
  wire \adder_32bit_0.operator_A_17.A ;
  wire \adder_32bit_0.operator_A_17.B ;
  wire \adder_32bit_0.operator_A_17.G ;
  wire \adder_32bit_0.operator_A_17.P ;
  wire \adder_32bit_0.operator_A_18.A ;
  wire \adder_32bit_0.operator_A_18.B ;
  wire \adder_32bit_0.operator_A_18.G ;
  wire \adder_32bit_0.operator_A_18.P ;
  wire \adder_32bit_0.operator_A_19.A ;
  wire \adder_32bit_0.operator_A_19.B ;
  wire \adder_32bit_0.operator_A_19.G ;
  wire \adder_32bit_0.operator_A_19.P ;
  wire \adder_32bit_0.operator_A_2.A ;
  wire \adder_32bit_0.operator_A_2.B ;
  wire \adder_32bit_0.operator_A_2.G ;
  wire \adder_32bit_0.operator_A_2.P ;
  wire \adder_32bit_0.operator_A_20.A ;
  wire \adder_32bit_0.operator_A_20.B ;
  wire \adder_32bit_0.operator_A_20.G ;
  wire \adder_32bit_0.operator_A_20.P ;
  wire \adder_32bit_0.operator_A_21.A ;
  wire \adder_32bit_0.operator_A_21.B ;
  wire \adder_32bit_0.operator_A_21.G ;
  wire \adder_32bit_0.operator_A_21.P ;
  wire \adder_32bit_0.operator_A_22.A ;
  wire \adder_32bit_0.operator_A_22.B ;
  wire \adder_32bit_0.operator_A_22.G ;
  wire \adder_32bit_0.operator_A_22.P ;
  wire \adder_32bit_0.operator_A_23.A ;
  wire \adder_32bit_0.operator_A_23.B ;
  wire \adder_32bit_0.operator_A_23.G ;
  wire \adder_32bit_0.operator_A_23.P ;
  wire \adder_32bit_0.operator_A_24.A ;
  wire \adder_32bit_0.operator_A_24.B ;
  wire \adder_32bit_0.operator_A_24.G ;
  wire \adder_32bit_0.operator_A_24.P ;
  wire \adder_32bit_0.operator_A_25.A ;
  wire \adder_32bit_0.operator_A_25.B ;
  wire \adder_32bit_0.operator_A_25.G ;
  wire \adder_32bit_0.operator_A_25.P ;
  wire \adder_32bit_0.operator_A_26.A ;
  wire \adder_32bit_0.operator_A_26.B ;
  wire \adder_32bit_0.operator_A_26.G ;
  wire \adder_32bit_0.operator_A_26.P ;
  wire \adder_32bit_0.operator_A_27.A ;
  wire \adder_32bit_0.operator_A_27.B ;
  wire \adder_32bit_0.operator_A_27.G ;
  wire \adder_32bit_0.operator_A_27.P ;
  wire \adder_32bit_0.operator_A_28.A ;
  wire \adder_32bit_0.operator_A_28.B ;
  wire \adder_32bit_0.operator_A_28.G ;
  wire \adder_32bit_0.operator_A_28.P ;
  wire \adder_32bit_0.operator_A_29.A ;
  wire \adder_32bit_0.operator_A_29.B ;
  wire \adder_32bit_0.operator_A_29.G ;
  wire \adder_32bit_0.operator_A_29.P ;
  wire \adder_32bit_0.operator_A_3.A ;
  wire \adder_32bit_0.operator_A_3.B ;
  wire \adder_32bit_0.operator_A_3.G ;
  wire \adder_32bit_0.operator_A_3.P ;
  wire \adder_32bit_0.operator_A_30.A ;
  wire \adder_32bit_0.operator_A_30.B ;
  wire \adder_32bit_0.operator_A_30.G ;
  wire \adder_32bit_0.operator_A_30.P ;
  wire \adder_32bit_0.operator_A_31.A ;
  wire \adder_32bit_0.operator_A_31.B ;
  wire \adder_32bit_0.operator_A_31.P ;
  wire \adder_32bit_0.operator_A_4.A ;
  wire \adder_32bit_0.operator_A_4.B ;
  wire \adder_32bit_0.operator_A_4.G ;
  wire \adder_32bit_0.operator_A_4.P ;
  wire \adder_32bit_0.operator_A_5.A ;
  wire \adder_32bit_0.operator_A_5.B ;
  wire \adder_32bit_0.operator_A_5.G ;
  wire \adder_32bit_0.operator_A_5.P ;
  wire \adder_32bit_0.operator_A_6.A ;
  wire \adder_32bit_0.operator_A_6.B ;
  wire \adder_32bit_0.operator_A_6.G ;
  wire \adder_32bit_0.operator_A_6.P ;
  wire \adder_32bit_0.operator_A_7.A ;
  wire \adder_32bit_0.operator_A_7.B ;
  wire \adder_32bit_0.operator_A_7.G ;
  wire \adder_32bit_0.operator_A_7.P ;
  wire \adder_32bit_0.operator_A_8.A ;
  wire \adder_32bit_0.operator_A_8.B ;
  wire \adder_32bit_0.operator_A_8.G ;
  wire \adder_32bit_0.operator_A_8.P ;
  wire \adder_32bit_0.operator_A_9.A ;
  wire \adder_32bit_0.operator_A_9.B ;
  wire \adder_32bit_0.operator_A_9.G ;
  wire \adder_32bit_0.operator_A_9.P ;
  wire \adder_32bit_0.operator_B_stage_1_1.G ;
  wire \adder_32bit_0.operator_B_stage_1_1.G1 ;
  wire \adder_32bit_0.operator_B_stage_1_1.Go ;
  wire \adder_32bit_0.operator_B_stage_1_1.P ;
  wire \adder_32bit_0.operator_B_stage_1_1.P1 ;
  wire \adder_32bit_0.operator_B_stage_1_1.Po ;
  wire \adder_32bit_0.operator_B_stage_1_10.G ;
  wire \adder_32bit_0.operator_B_stage_1_10.G1 ;
  wire \adder_32bit_0.operator_B_stage_1_10.Go ;
  wire \adder_32bit_0.operator_B_stage_1_10.P ;
  wire \adder_32bit_0.operator_B_stage_1_10.P1 ;
  wire \adder_32bit_0.operator_B_stage_1_10.Po ;
  wire \adder_32bit_0.operator_B_stage_1_11.G ;
  wire \adder_32bit_0.operator_B_stage_1_11.G1 ;
  wire \adder_32bit_0.operator_B_stage_1_11.Go ;
  wire \adder_32bit_0.operator_B_stage_1_11.P ;
  wire \adder_32bit_0.operator_B_stage_1_11.P1 ;
  wire \adder_32bit_0.operator_B_stage_1_11.Po ;
  wire \adder_32bit_0.operator_B_stage_1_12.G ;
  wire \adder_32bit_0.operator_B_stage_1_12.G1 ;
  wire \adder_32bit_0.operator_B_stage_1_12.Go ;
  wire \adder_32bit_0.operator_B_stage_1_12.P ;
  wire \adder_32bit_0.operator_B_stage_1_12.P1 ;
  wire \adder_32bit_0.operator_B_stage_1_12.Po ;
  wire \adder_32bit_0.operator_B_stage_1_13.G ;
  wire \adder_32bit_0.operator_B_stage_1_13.G1 ;
  wire \adder_32bit_0.operator_B_stage_1_13.Go ;
  wire \adder_32bit_0.operator_B_stage_1_13.P ;
  wire \adder_32bit_0.operator_B_stage_1_13.P1 ;
  wire \adder_32bit_0.operator_B_stage_1_13.Po ;
  wire \adder_32bit_0.operator_B_stage_1_14.G ;
  wire \adder_32bit_0.operator_B_stage_1_14.G1 ;
  wire \adder_32bit_0.operator_B_stage_1_14.Go ;
  wire \adder_32bit_0.operator_B_stage_1_14.P ;
  wire \adder_32bit_0.operator_B_stage_1_14.P1 ;
  wire \adder_32bit_0.operator_B_stage_1_14.Po ;
  wire \adder_32bit_0.operator_B_stage_1_15.G ;
  wire \adder_32bit_0.operator_B_stage_1_15.G1 ;
  wire \adder_32bit_0.operator_B_stage_1_15.Go ;
  wire \adder_32bit_0.operator_B_stage_1_15.P ;
  wire \adder_32bit_0.operator_B_stage_1_15.P1 ;
  wire \adder_32bit_0.operator_B_stage_1_15.Po ;
  wire \adder_32bit_0.operator_B_stage_1_2.G ;
  wire \adder_32bit_0.operator_B_stage_1_2.G1 ;
  wire \adder_32bit_0.operator_B_stage_1_2.Go ;
  wire \adder_32bit_0.operator_B_stage_1_2.P ;
  wire \adder_32bit_0.operator_B_stage_1_2.P1 ;
  wire \adder_32bit_0.operator_B_stage_1_2.Po ;
  wire \adder_32bit_0.operator_B_stage_1_3.G ;
  wire \adder_32bit_0.operator_B_stage_1_3.G1 ;
  wire \adder_32bit_0.operator_B_stage_1_3.Go ;
  wire \adder_32bit_0.operator_B_stage_1_3.P ;
  wire \adder_32bit_0.operator_B_stage_1_3.P1 ;
  wire \adder_32bit_0.operator_B_stage_1_3.Po ;
  wire \adder_32bit_0.operator_B_stage_1_4.G ;
  wire \adder_32bit_0.operator_B_stage_1_4.G1 ;
  wire \adder_32bit_0.operator_B_stage_1_4.Go ;
  wire \adder_32bit_0.operator_B_stage_1_4.P ;
  wire \adder_32bit_0.operator_B_stage_1_4.P1 ;
  wire \adder_32bit_0.operator_B_stage_1_4.Po ;
  wire \adder_32bit_0.operator_B_stage_1_5.G ;
  wire \adder_32bit_0.operator_B_stage_1_5.G1 ;
  wire \adder_32bit_0.operator_B_stage_1_5.Go ;
  wire \adder_32bit_0.operator_B_stage_1_5.P ;
  wire \adder_32bit_0.operator_B_stage_1_5.P1 ;
  wire \adder_32bit_0.operator_B_stage_1_5.Po ;
  wire \adder_32bit_0.operator_B_stage_1_6.G ;
  wire \adder_32bit_0.operator_B_stage_1_6.G1 ;
  wire \adder_32bit_0.operator_B_stage_1_6.Go ;
  wire \adder_32bit_0.operator_B_stage_1_6.P ;
  wire \adder_32bit_0.operator_B_stage_1_6.P1 ;
  wire \adder_32bit_0.operator_B_stage_1_6.Po ;
  wire \adder_32bit_0.operator_B_stage_1_7.G ;
  wire \adder_32bit_0.operator_B_stage_1_7.G1 ;
  wire \adder_32bit_0.operator_B_stage_1_7.Go ;
  wire \adder_32bit_0.operator_B_stage_1_7.P ;
  wire \adder_32bit_0.operator_B_stage_1_7.P1 ;
  wire \adder_32bit_0.operator_B_stage_1_7.Po ;
  wire \adder_32bit_0.operator_B_stage_1_8.G ;
  wire \adder_32bit_0.operator_B_stage_1_8.G1 ;
  wire \adder_32bit_0.operator_B_stage_1_8.Go ;
  wire \adder_32bit_0.operator_B_stage_1_8.P ;
  wire \adder_32bit_0.operator_B_stage_1_8.P1 ;
  wire \adder_32bit_0.operator_B_stage_1_8.Po ;
  wire \adder_32bit_0.operator_B_stage_1_9.G ;
  wire \adder_32bit_0.operator_B_stage_1_9.G1 ;
  wire \adder_32bit_0.operator_B_stage_1_9.Go ;
  wire \adder_32bit_0.operator_B_stage_1_9.P ;
  wire \adder_32bit_0.operator_B_stage_1_9.P1 ;
  wire \adder_32bit_0.operator_B_stage_1_9.Po ;
  wire \adder_32bit_0.operator_B_stage_2_10.G ;
  wire \adder_32bit_0.operator_B_stage_2_10.G1 ;
  wire \adder_32bit_0.operator_B_stage_2_10.Go ;
  wire \adder_32bit_0.operator_B_stage_2_10.P ;
  wire \adder_32bit_0.operator_B_stage_2_10.P1 ;
  wire \adder_32bit_0.operator_B_stage_2_10.Po ;
  wire \adder_32bit_0.operator_B_stage_2_11.G ;
  wire \adder_32bit_0.operator_B_stage_2_11.G1 ;
  wire \adder_32bit_0.operator_B_stage_2_11.Go ;
  wire \adder_32bit_0.operator_B_stage_2_11.P ;
  wire \adder_32bit_0.operator_B_stage_2_11.P1 ;
  wire \adder_32bit_0.operator_B_stage_2_11.Po ;
  wire \adder_32bit_0.operator_B_stage_2_12.G ;
  wire \adder_32bit_0.operator_B_stage_2_12.G1 ;
  wire \adder_32bit_0.operator_B_stage_2_12.Go ;
  wire \adder_32bit_0.operator_B_stage_2_12.P ;
  wire \adder_32bit_0.operator_B_stage_2_12.P1 ;
  wire \adder_32bit_0.operator_B_stage_2_12.Po ;
  wire \adder_32bit_0.operator_B_stage_2_13.G ;
  wire \adder_32bit_0.operator_B_stage_2_13.G1 ;
  wire \adder_32bit_0.operator_B_stage_2_13.Go ;
  wire \adder_32bit_0.operator_B_stage_2_13.P ;
  wire \adder_32bit_0.operator_B_stage_2_13.P1 ;
  wire \adder_32bit_0.operator_B_stage_2_13.Po ;
  wire \adder_32bit_0.operator_B_stage_2_14.G ;
  wire \adder_32bit_0.operator_B_stage_2_14.G1 ;
  wire \adder_32bit_0.operator_B_stage_2_14.Go ;
  wire \adder_32bit_0.operator_B_stage_2_14.P ;
  wire \adder_32bit_0.operator_B_stage_2_14.P1 ;
  wire \adder_32bit_0.operator_B_stage_2_14.Po ;
  wire \adder_32bit_0.operator_B_stage_2_15.G ;
  wire \adder_32bit_0.operator_B_stage_2_15.G1 ;
  wire \adder_32bit_0.operator_B_stage_2_15.Go ;
  wire \adder_32bit_0.operator_B_stage_2_15.P ;
  wire \adder_32bit_0.operator_B_stage_2_15.P1 ;
  wire \adder_32bit_0.operator_B_stage_2_15.Po ;
  wire \adder_32bit_0.operator_B_stage_2_2.G ;
  wire \adder_32bit_0.operator_B_stage_2_2.G1 ;
  wire \adder_32bit_0.operator_B_stage_2_2.Go ;
  wire \adder_32bit_0.operator_B_stage_2_2.P ;
  wire \adder_32bit_0.operator_B_stage_2_2.P1 ;
  wire \adder_32bit_0.operator_B_stage_2_2.Po ;
  wire \adder_32bit_0.operator_B_stage_2_3.G ;
  wire \adder_32bit_0.operator_B_stage_2_3.G1 ;
  wire \adder_32bit_0.operator_B_stage_2_3.Go ;
  wire \adder_32bit_0.operator_B_stage_2_3.P ;
  wire \adder_32bit_0.operator_B_stage_2_3.P1 ;
  wire \adder_32bit_0.operator_B_stage_2_3.Po ;
  wire \adder_32bit_0.operator_B_stage_2_4.G ;
  wire \adder_32bit_0.operator_B_stage_2_4.G1 ;
  wire \adder_32bit_0.operator_B_stage_2_4.Go ;
  wire \adder_32bit_0.operator_B_stage_2_4.P ;
  wire \adder_32bit_0.operator_B_stage_2_4.P1 ;
  wire \adder_32bit_0.operator_B_stage_2_4.Po ;
  wire \adder_32bit_0.operator_B_stage_2_5.G ;
  wire \adder_32bit_0.operator_B_stage_2_5.G1 ;
  wire \adder_32bit_0.operator_B_stage_2_5.Go ;
  wire \adder_32bit_0.operator_B_stage_2_5.P ;
  wire \adder_32bit_0.operator_B_stage_2_5.P1 ;
  wire \adder_32bit_0.operator_B_stage_2_5.Po ;
  wire \adder_32bit_0.operator_B_stage_2_6.G ;
  wire \adder_32bit_0.operator_B_stage_2_6.G1 ;
  wire \adder_32bit_0.operator_B_stage_2_6.Go ;
  wire \adder_32bit_0.operator_B_stage_2_6.P ;
  wire \adder_32bit_0.operator_B_stage_2_6.P1 ;
  wire \adder_32bit_0.operator_B_stage_2_6.Po ;
  wire \adder_32bit_0.operator_B_stage_2_7.G ;
  wire \adder_32bit_0.operator_B_stage_2_7.G1 ;
  wire \adder_32bit_0.operator_B_stage_2_7.Go ;
  wire \adder_32bit_0.operator_B_stage_2_7.P ;
  wire \adder_32bit_0.operator_B_stage_2_7.P1 ;
  wire \adder_32bit_0.operator_B_stage_2_7.Po ;
  wire \adder_32bit_0.operator_B_stage_2_8.G ;
  wire \adder_32bit_0.operator_B_stage_2_8.G1 ;
  wire \adder_32bit_0.operator_B_stage_2_8.Go ;
  wire \adder_32bit_0.operator_B_stage_2_8.P ;
  wire \adder_32bit_0.operator_B_stage_2_8.P1 ;
  wire \adder_32bit_0.operator_B_stage_2_8.Po ;
  wire \adder_32bit_0.operator_B_stage_2_9.G ;
  wire \adder_32bit_0.operator_B_stage_2_9.G1 ;
  wire \adder_32bit_0.operator_B_stage_2_9.Go ;
  wire \adder_32bit_0.operator_B_stage_2_9.P ;
  wire \adder_32bit_0.operator_B_stage_2_9.P1 ;
  wire \adder_32bit_0.operator_B_stage_2_9.Po ;
  wire \adder_32bit_0.operator_B_stage_3_10.G ;
  wire \adder_32bit_0.operator_B_stage_3_10.G1 ;
  wire \adder_32bit_0.operator_B_stage_3_10.Go ;
  wire \adder_32bit_0.operator_B_stage_3_10.P ;
  wire \adder_32bit_0.operator_B_stage_3_10.P1 ;
  wire \adder_32bit_0.operator_B_stage_3_10.Po ;
  wire \adder_32bit_0.operator_B_stage_3_11.G ;
  wire \adder_32bit_0.operator_B_stage_3_11.G1 ;
  wire \adder_32bit_0.operator_B_stage_3_11.Go ;
  wire \adder_32bit_0.operator_B_stage_3_11.P ;
  wire \adder_32bit_0.operator_B_stage_3_11.P1 ;
  wire \adder_32bit_0.operator_B_stage_3_11.Po ;
  wire \adder_32bit_0.operator_B_stage_3_12.G ;
  wire \adder_32bit_0.operator_B_stage_3_12.G1 ;
  wire \adder_32bit_0.operator_B_stage_3_12.Go ;
  wire \adder_32bit_0.operator_B_stage_3_12.P ;
  wire \adder_32bit_0.operator_B_stage_3_12.P1 ;
  wire \adder_32bit_0.operator_B_stage_3_12.Po ;
  wire \adder_32bit_0.operator_B_stage_3_13.G ;
  wire \adder_32bit_0.operator_B_stage_3_13.G1 ;
  wire \adder_32bit_0.operator_B_stage_3_13.Go ;
  wire \adder_32bit_0.operator_B_stage_3_13.P ;
  wire \adder_32bit_0.operator_B_stage_3_13.P1 ;
  wire \adder_32bit_0.operator_B_stage_3_13.Po ;
  wire \adder_32bit_0.operator_B_stage_3_14.G ;
  wire \adder_32bit_0.operator_B_stage_3_14.G1 ;
  wire \adder_32bit_0.operator_B_stage_3_14.Go ;
  wire \adder_32bit_0.operator_B_stage_3_14.P ;
  wire \adder_32bit_0.operator_B_stage_3_14.P1 ;
  wire \adder_32bit_0.operator_B_stage_3_14.Po ;
  wire \adder_32bit_0.operator_B_stage_3_15.G ;
  wire \adder_32bit_0.operator_B_stage_3_15.G1 ;
  wire \adder_32bit_0.operator_B_stage_3_15.Go ;
  wire \adder_32bit_0.operator_B_stage_3_15.P ;
  wire \adder_32bit_0.operator_B_stage_3_15.P1 ;
  wire \adder_32bit_0.operator_B_stage_3_15.Po ;
  wire \adder_32bit_0.operator_B_stage_3_4.G ;
  wire \adder_32bit_0.operator_B_stage_3_4.G1 ;
  wire \adder_32bit_0.operator_B_stage_3_4.Go ;
  wire \adder_32bit_0.operator_B_stage_3_4.P ;
  wire \adder_32bit_0.operator_B_stage_3_4.P1 ;
  wire \adder_32bit_0.operator_B_stage_3_4.Po ;
  wire \adder_32bit_0.operator_B_stage_3_5.G ;
  wire \adder_32bit_0.operator_B_stage_3_5.G1 ;
  wire \adder_32bit_0.operator_B_stage_3_5.Go ;
  wire \adder_32bit_0.operator_B_stage_3_5.P ;
  wire \adder_32bit_0.operator_B_stage_3_5.P1 ;
  wire \adder_32bit_0.operator_B_stage_3_5.Po ;
  wire \adder_32bit_0.operator_B_stage_3_6.G ;
  wire \adder_32bit_0.operator_B_stage_3_6.G1 ;
  wire \adder_32bit_0.operator_B_stage_3_6.Go ;
  wire \adder_32bit_0.operator_B_stage_3_6.P ;
  wire \adder_32bit_0.operator_B_stage_3_6.P1 ;
  wire \adder_32bit_0.operator_B_stage_3_6.Po ;
  wire \adder_32bit_0.operator_B_stage_3_7.G ;
  wire \adder_32bit_0.operator_B_stage_3_7.G1 ;
  wire \adder_32bit_0.operator_B_stage_3_7.Go ;
  wire \adder_32bit_0.operator_B_stage_3_7.P ;
  wire \adder_32bit_0.operator_B_stage_3_7.P1 ;
  wire \adder_32bit_0.operator_B_stage_3_7.Po ;
  wire \adder_32bit_0.operator_B_stage_3_8.G ;
  wire \adder_32bit_0.operator_B_stage_3_8.G1 ;
  wire \adder_32bit_0.operator_B_stage_3_8.Go ;
  wire \adder_32bit_0.operator_B_stage_3_8.P ;
  wire \adder_32bit_0.operator_B_stage_3_8.P1 ;
  wire \adder_32bit_0.operator_B_stage_3_8.Po ;
  wire \adder_32bit_0.operator_B_stage_3_9.G ;
  wire \adder_32bit_0.operator_B_stage_3_9.G1 ;
  wire \adder_32bit_0.operator_B_stage_3_9.Go ;
  wire \adder_32bit_0.operator_B_stage_3_9.P ;
  wire \adder_32bit_0.operator_B_stage_3_9.P1 ;
  wire \adder_32bit_0.operator_B_stage_3_9.Po ;
  wire \adder_32bit_0.operator_B_stage_4_10.G ;
  wire \adder_32bit_0.operator_B_stage_4_10.G1 ;
  wire \adder_32bit_0.operator_B_stage_4_10.Go ;
  wire \adder_32bit_0.operator_B_stage_4_10.P ;
  wire \adder_32bit_0.operator_B_stage_4_10.P1 ;
  wire \adder_32bit_0.operator_B_stage_4_10.Po ;
  wire \adder_32bit_0.operator_B_stage_4_11.G ;
  wire \adder_32bit_0.operator_B_stage_4_11.G1 ;
  wire \adder_32bit_0.operator_B_stage_4_11.Go ;
  wire \adder_32bit_0.operator_B_stage_4_11.P ;
  wire \adder_32bit_0.operator_B_stage_4_11.P1 ;
  wire \adder_32bit_0.operator_B_stage_4_11.Po ;
  wire \adder_32bit_0.operator_B_stage_4_12.G ;
  wire \adder_32bit_0.operator_B_stage_4_12.G1 ;
  wire \adder_32bit_0.operator_B_stage_4_12.Go ;
  wire \adder_32bit_0.operator_B_stage_4_12.P ;
  wire \adder_32bit_0.operator_B_stage_4_12.P1 ;
  wire \adder_32bit_0.operator_B_stage_4_12.Po ;
  wire \adder_32bit_0.operator_B_stage_4_13.G ;
  wire \adder_32bit_0.operator_B_stage_4_13.G1 ;
  wire \adder_32bit_0.operator_B_stage_4_13.Go ;
  wire \adder_32bit_0.operator_B_stage_4_13.P ;
  wire \adder_32bit_0.operator_B_stage_4_13.P1 ;
  wire \adder_32bit_0.operator_B_stage_4_13.Po ;
  wire \adder_32bit_0.operator_B_stage_4_14.G ;
  wire \adder_32bit_0.operator_B_stage_4_14.G1 ;
  wire \adder_32bit_0.operator_B_stage_4_14.Go ;
  wire \adder_32bit_0.operator_B_stage_4_14.P ;
  wire \adder_32bit_0.operator_B_stage_4_14.P1 ;
  wire \adder_32bit_0.operator_B_stage_4_14.Po ;
  wire \adder_32bit_0.operator_B_stage_4_15.G ;
  wire \adder_32bit_0.operator_B_stage_4_15.G1 ;
  wire \adder_32bit_0.operator_B_stage_4_15.Go ;
  wire \adder_32bit_0.operator_B_stage_4_15.P ;
  wire \adder_32bit_0.operator_B_stage_4_15.P1 ;
  wire \adder_32bit_0.operator_B_stage_4_15.Po ;
  wire \adder_32bit_0.operator_B_stage_4_8.G ;
  wire \adder_32bit_0.operator_B_stage_4_8.G1 ;
  wire \adder_32bit_0.operator_B_stage_4_8.Go ;
  wire \adder_32bit_0.operator_B_stage_4_8.P ;
  wire \adder_32bit_0.operator_B_stage_4_8.P1 ;
  wire \adder_32bit_0.operator_B_stage_4_8.Po ;
  wire \adder_32bit_0.operator_B_stage_4_9.G ;
  wire \adder_32bit_0.operator_B_stage_4_9.G1 ;
  wire \adder_32bit_0.operator_B_stage_4_9.Go ;
  wire \adder_32bit_0.operator_B_stage_4_9.P ;
  wire \adder_32bit_0.operator_B_stage_4_9.P1 ;
  wire \adder_32bit_0.operator_B_stage_4_9.Po ;
  wire \adder_32bit_0.operator_C_stage_1_0.G ;
  wire \adder_32bit_0.operator_C_stage_1_0.G1 ;
  wire \adder_32bit_0.operator_C_stage_1_0.Go ;
  wire \adder_32bit_0.operator_C_stage_1_0.P ;
  wire \adder_32bit_0.operator_C_stage_2_1.G ;
  wire \adder_32bit_0.operator_C_stage_2_1.G1 ;
  wire \adder_32bit_0.operator_C_stage_2_1.Go ;
  wire \adder_32bit_0.operator_C_stage_2_1.P ;
  wire \adder_32bit_0.operator_C_stage_3_2.G ;
  wire \adder_32bit_0.operator_C_stage_3_2.G1 ;
  wire \adder_32bit_0.operator_C_stage_3_2.Go ;
  wire \adder_32bit_0.operator_C_stage_3_2.P ;
  wire \adder_32bit_0.operator_C_stage_3_3.G ;
  wire \adder_32bit_0.operator_C_stage_3_3.G1 ;
  wire \adder_32bit_0.operator_C_stage_3_3.Go ;
  wire \adder_32bit_0.operator_C_stage_3_3.P ;
  wire \adder_32bit_0.operator_C_stage_4_4.G ;
  wire \adder_32bit_0.operator_C_stage_4_4.G1 ;
  wire \adder_32bit_0.operator_C_stage_4_4.Go ;
  wire \adder_32bit_0.operator_C_stage_4_4.P ;
  wire \adder_32bit_0.operator_C_stage_4_5.G ;
  wire \adder_32bit_0.operator_C_stage_4_5.G1 ;
  wire \adder_32bit_0.operator_C_stage_4_5.Go ;
  wire \adder_32bit_0.operator_C_stage_4_5.P ;
  wire \adder_32bit_0.operator_C_stage_4_6.G ;
  wire \adder_32bit_0.operator_C_stage_4_6.G1 ;
  wire \adder_32bit_0.operator_C_stage_4_6.Go ;
  wire \adder_32bit_0.operator_C_stage_4_6.P ;
  wire \adder_32bit_0.operator_C_stage_4_7.G ;
  wire \adder_32bit_0.operator_C_stage_4_7.G1 ;
  wire \adder_32bit_0.operator_C_stage_4_7.Go ;
  wire \adder_32bit_0.operator_C_stage_4_7.P ;
  wire \adder_32bit_0.operator_C_stage_5_10.G ;
  wire \adder_32bit_0.operator_C_stage_5_10.G1 ;
  wire \adder_32bit_0.operator_C_stage_5_10.Go ;
  wire \adder_32bit_0.operator_C_stage_5_10.P ;
  wire \adder_32bit_0.operator_C_stage_5_11.G ;
  wire \adder_32bit_0.operator_C_stage_5_11.G1 ;
  wire \adder_32bit_0.operator_C_stage_5_11.Go ;
  wire \adder_32bit_0.operator_C_stage_5_11.P ;
  wire \adder_32bit_0.operator_C_stage_5_12.G ;
  wire \adder_32bit_0.operator_C_stage_5_12.G1 ;
  wire \adder_32bit_0.operator_C_stage_5_12.Go ;
  wire \adder_32bit_0.operator_C_stage_5_12.P ;
  wire \adder_32bit_0.operator_C_stage_5_13.G ;
  wire \adder_32bit_0.operator_C_stage_5_13.G1 ;
  wire \adder_32bit_0.operator_C_stage_5_13.Go ;
  wire \adder_32bit_0.operator_C_stage_5_13.P ;
  wire \adder_32bit_0.operator_C_stage_5_14.G ;
  wire \adder_32bit_0.operator_C_stage_5_14.G1 ;
  wire \adder_32bit_0.operator_C_stage_5_14.Go ;
  wire \adder_32bit_0.operator_C_stage_5_14.P ;
  wire \adder_32bit_0.operator_C_stage_5_15.G ;
  wire \adder_32bit_0.operator_C_stage_5_15.G1 ;
  wire \adder_32bit_0.operator_C_stage_5_15.Go ;
  wire \adder_32bit_0.operator_C_stage_5_15.P ;
  wire \adder_32bit_0.operator_C_stage_5_8.G ;
  wire \adder_32bit_0.operator_C_stage_5_8.G1 ;
  wire \adder_32bit_0.operator_C_stage_5_8.Go ;
  wire \adder_32bit_0.operator_C_stage_5_8.P ;
  wire \adder_32bit_0.operator_C_stage_5_9.G ;
  wire \adder_32bit_0.operator_C_stage_5_9.G1 ;
  wire \adder_32bit_0.operator_C_stage_5_9.Go ;
  wire \adder_32bit_0.operator_C_stage_5_9.P ;
  wire \adder_32bit_0.operator_C_stage_6_0.G ;
  wire \adder_32bit_0.operator_C_stage_6_0.G1 ;
  wire \adder_32bit_0.operator_C_stage_6_0.Go ;
  wire \adder_32bit_0.operator_C_stage_6_0.P ;
  wire \adder_32bit_0.operator_C_stage_6_1.G ;
  wire \adder_32bit_0.operator_C_stage_6_1.G1 ;
  wire \adder_32bit_0.operator_C_stage_6_1.Go ;
  wire \adder_32bit_0.operator_C_stage_6_1.P ;
  wire \adder_32bit_0.operator_C_stage_6_10.G ;
  wire \adder_32bit_0.operator_C_stage_6_10.G1 ;
  wire \adder_32bit_0.operator_C_stage_6_10.Go ;
  wire \adder_32bit_0.operator_C_stage_6_10.P ;
  wire \adder_32bit_0.operator_C_stage_6_11.G ;
  wire \adder_32bit_0.operator_C_stage_6_11.G1 ;
  wire \adder_32bit_0.operator_C_stage_6_11.Go ;
  wire \adder_32bit_0.operator_C_stage_6_11.P ;
  wire \adder_32bit_0.operator_C_stage_6_12.G ;
  wire \adder_32bit_0.operator_C_stage_6_12.G1 ;
  wire \adder_32bit_0.operator_C_stage_6_12.Go ;
  wire \adder_32bit_0.operator_C_stage_6_12.P ;
  wire \adder_32bit_0.operator_C_stage_6_13.G ;
  wire \adder_32bit_0.operator_C_stage_6_13.G1 ;
  wire \adder_32bit_0.operator_C_stage_6_13.Go ;
  wire \adder_32bit_0.operator_C_stage_6_13.P ;
  wire \adder_32bit_0.operator_C_stage_6_14.G ;
  wire \adder_32bit_0.operator_C_stage_6_14.G1 ;
  wire \adder_32bit_0.operator_C_stage_6_14.Go ;
  wire \adder_32bit_0.operator_C_stage_6_14.P ;
  wire \adder_32bit_0.operator_C_stage_6_15.G1 ;
  wire \adder_32bit_0.operator_C_stage_6_15.P ;
  wire \adder_32bit_0.operator_C_stage_6_2.G ;
  wire \adder_32bit_0.operator_C_stage_6_2.G1 ;
  wire \adder_32bit_0.operator_C_stage_6_2.Go ;
  wire \adder_32bit_0.operator_C_stage_6_2.P ;
  wire \adder_32bit_0.operator_C_stage_6_3.G ;
  wire \adder_32bit_0.operator_C_stage_6_3.G1 ;
  wire \adder_32bit_0.operator_C_stage_6_3.Go ;
  wire \adder_32bit_0.operator_C_stage_6_3.P ;
  wire \adder_32bit_0.operator_C_stage_6_4.G ;
  wire \adder_32bit_0.operator_C_stage_6_4.G1 ;
  wire \adder_32bit_0.operator_C_stage_6_4.Go ;
  wire \adder_32bit_0.operator_C_stage_6_4.P ;
  wire \adder_32bit_0.operator_C_stage_6_5.G ;
  wire \adder_32bit_0.operator_C_stage_6_5.G1 ;
  wire \adder_32bit_0.operator_C_stage_6_5.Go ;
  wire \adder_32bit_0.operator_C_stage_6_5.P ;
  wire \adder_32bit_0.operator_C_stage_6_6.G ;
  wire \adder_32bit_0.operator_C_stage_6_6.G1 ;
  wire \adder_32bit_0.operator_C_stage_6_6.Go ;
  wire \adder_32bit_0.operator_C_stage_6_6.P ;
  wire \adder_32bit_0.operator_C_stage_6_7.G ;
  wire \adder_32bit_0.operator_C_stage_6_7.G1 ;
  wire \adder_32bit_0.operator_C_stage_6_7.Go ;
  wire \adder_32bit_0.operator_C_stage_6_7.P ;
  wire \adder_32bit_0.operator_C_stage_6_8.G ;
  wire \adder_32bit_0.operator_C_stage_6_8.G1 ;
  wire \adder_32bit_0.operator_C_stage_6_8.Go ;
  wire \adder_32bit_0.operator_C_stage_6_8.P ;
  wire \adder_32bit_0.operator_C_stage_6_9.G ;
  wire \adder_32bit_0.operator_C_stage_6_9.G1 ;
  wire \adder_32bit_0.operator_C_stage_6_9.Go ;
  wire \adder_32bit_0.operator_C_stage_6_9.P ;
  wire [2:0] adr;
  wire [3:0] adr_1;
  wire adr_check;
  wire adr_check_1;
  reg cout;
  reg [15:0] \err[0] ;
  reg [15:0] \err[1] ;
  input i_clk;
  input i_rst;
  input [15:0] i_wb_adr;
  input i_wb_cyc;
  input [31:0] i_wb_data;
  input i_wb_stb;
  input i_wb_we;
  reg [15:0] kd;
  reg [15:0] ki;
  reg [15:0] kp;
  reg [15:0] kpd;
  wire [15:0] md;
  reg [1:0] md_index;
  wire [15:0] mr;
  reg [1:0] mr_index;
  wire [31:0] \multiplier_16x16bit_pipelined.A ;
  wire [30:0] \multiplier_16x16bit_pipelined.B ;
  wire [31:0] \multiplier_16x16bit_pipelined.adder_32bit.G0 ;
  wire [15:0] \multiplier_16x16bit_pipelined.adder_32bit.G1 ;
  wire [15:0] \multiplier_16x16bit_pipelined.adder_32bit.G2 ;
  wire [15:0] \multiplier_16x16bit_pipelined.adder_32bit.G3 ;
  wire [15:0] \multiplier_16x16bit_pipelined.adder_32bit.G4 ;
  wire [15:0] \multiplier_16x16bit_pipelined.adder_32bit.G5 ;
  wire [31:0] \multiplier_16x16bit_pipelined.adder_32bit.G6 ;
  wire [31:0] \multiplier_16x16bit_pipelined.adder_32bit.P0 ;
  wire [15:1] \multiplier_16x16bit_pipelined.adder_32bit.P1 ;
  wire [15:2] \multiplier_16x16bit_pipelined.adder_32bit.P2 ;
  wire [15:4] \multiplier_16x16bit_pipelined.adder_32bit.P3 ;
  wire [15:8] \multiplier_16x16bit_pipelined.adder_32bit.P4 ;
  wire [31:0] \multiplier_16x16bit_pipelined.adder_32bit.i_a ;
  wire [31:0] \multiplier_16x16bit_pipelined.adder_32bit.i_b ;
  wire [31:0] \multiplier_16x16bit_pipelined.adder_32bit.o_s ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_A_0.A ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_A_0.B ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_A_0.G ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_A_0.P ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_A_1.A ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_A_1.P ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_A_10.A ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_A_10.B ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_A_10.G ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_A_10.P ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_A_11.A ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_A_11.B ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_A_11.G ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_A_11.P ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_A_12.A ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_A_12.B ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_A_12.G ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_A_12.P ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_A_13.A ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_A_13.B ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_A_13.G ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_A_13.P ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_A_14.A ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_A_14.B ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_A_14.G ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_A_14.P ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_A_15.A ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_A_15.B ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_A_15.G ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_A_15.P ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_A_16.A ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_A_16.B ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_A_16.G ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_A_16.P ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_A_17.A ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_A_17.B ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_A_17.G ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_A_17.P ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_A_18.A ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_A_18.B ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_A_18.G ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_A_18.P ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_A_19.A ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_A_19.B ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_A_19.G ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_A_19.P ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_A_2.A ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_A_2.P ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_A_20.A ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_A_20.B ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_A_20.G ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_A_20.P ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_A_21.A ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_A_21.B ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_A_21.G ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_A_21.P ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_A_22.A ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_A_22.B ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_A_22.G ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_A_22.P ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_A_23.A ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_A_23.B ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_A_23.G ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_A_23.P ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_A_24.A ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_A_24.B ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_A_24.G ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_A_24.P ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_A_25.A ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_A_25.P ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_A_26.A ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_A_26.B ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_A_26.G ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_A_26.P ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_A_27.A ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_A_27.P ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_A_28.A ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_A_28.B ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_A_28.G ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_A_28.P ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_A_29.A ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_A_29.P ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_A_3.A ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_A_3.B ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_A_3.G ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_A_3.P ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_A_30.A ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_A_30.B ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_A_30.G ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_A_30.P ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_A_31.A ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_A_31.P ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_A_4.A ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_A_4.B ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_A_4.G ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_A_4.P ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_A_5.A ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_A_5.B ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_A_5.G ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_A_5.P ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_A_6.A ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_A_6.B ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_A_6.G ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_A_6.P ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_A_7.A ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_A_7.B ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_A_7.G ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_A_7.P ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_A_8.A ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_A_8.B ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_A_8.G ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_A_8.P ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_A_9.A ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_A_9.B ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_A_9.G ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_A_9.P ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_1.P ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_1.P1 ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_1.Po ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_10.G ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_10.G1 ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_10.Go ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_10.P ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_10.P1 ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_10.Po ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_11.G ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_11.G1 ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_11.Go ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_11.P ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_11.P1 ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_11.Po ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_12.G ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_12.G1 ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_12.Go ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_12.P ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_12.P1 ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_12.Po ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_13.G ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_13.Go ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_13.P ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_13.P1 ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_13.Po ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_14.G ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_14.Go ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_14.P ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_14.P1 ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_14.Po ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_15.G ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_15.Go ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_15.P ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_15.P1 ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_15.Po ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_2.G ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_2.G1 ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_2.Go ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_2.P ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_2.P1 ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_2.Po ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_3.G ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_3.G1 ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_3.Go ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_3.P ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_3.P1 ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_3.Po ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_4.G ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_4.G1 ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_4.Go ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_4.P ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_4.P1 ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_4.Po ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_5.G ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_5.G1 ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_5.Go ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_5.P ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_5.P1 ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_5.Po ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_6.G ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_6.G1 ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_6.Go ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_6.P ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_6.P1 ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_6.Po ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_7.G ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_7.G1 ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_7.Go ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_7.P ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_7.P1 ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_7.Po ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_8.G ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_8.G1 ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_8.Go ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_8.P ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_8.P1 ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_8.Po ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_9.G ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_9.G1 ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_9.Go ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_9.P ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_9.P1 ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_9.Po ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_10.G ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_10.G1 ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_10.Go ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_10.P ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_10.P1 ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_10.Po ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_11.G ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_11.G1 ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_11.Go ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_11.P ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_11.P1 ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_11.Po ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_12.G ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_12.G1 ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_12.Go ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_12.P ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_12.P1 ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_12.Po ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_13.G ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_13.G1 ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_13.Go ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_13.P ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_13.P1 ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_13.Po ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_14.G ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_14.G1 ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_14.Go ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_14.P ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_14.P1 ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_14.Po ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_15.G ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_15.G1 ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_15.Go ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_15.P ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_15.P1 ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_15.Po ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_2.G ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_2.Go ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_2.P ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_2.P1 ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_2.Po ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_3.G ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_3.G1 ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_3.Go ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_3.P ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_3.P1 ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_3.Po ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_4.G ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_4.G1 ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_4.Go ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_4.P ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_4.P1 ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_4.Po ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_5.G ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_5.G1 ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_5.Go ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_5.P ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_5.P1 ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_5.Po ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_6.G ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_6.G1 ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_6.Go ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_6.P ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_6.P1 ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_6.Po ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_7.G ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_7.G1 ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_7.Go ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_7.P ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_7.P1 ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_7.Po ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_8.G ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_8.G1 ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_8.Go ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_8.P ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_8.P1 ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_8.Po ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_9.G ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_9.G1 ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_9.Go ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_9.P ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_9.P1 ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_9.Po ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_10.G ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_10.G1 ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_10.Go ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_10.P ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_10.P1 ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_10.Po ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_11.G ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_11.G1 ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_11.Go ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_11.P ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_11.P1 ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_11.Po ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_12.G ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_12.G1 ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_12.Go ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_12.P ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_12.P1 ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_12.Po ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_13.G ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_13.G1 ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_13.Go ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_13.P ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_13.P1 ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_13.Po ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_14.G ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_14.G1 ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_14.Go ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_14.P ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_14.P1 ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_14.Po ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_15.G ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_15.G1 ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_15.Go ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_15.P ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_15.P1 ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_15.Po ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_4.G ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_4.G1 ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_4.Go ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_4.P ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_4.P1 ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_4.Po ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_5.G ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_5.G1 ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_5.Go ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_5.P ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_5.P1 ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_5.Po ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_6.G ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_6.G1 ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_6.Go ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_6.P ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_6.P1 ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_6.Po ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_7.G ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_7.G1 ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_7.Go ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_7.P ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_7.P1 ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_7.Po ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_8.G ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_8.G1 ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_8.Go ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_8.P ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_8.P1 ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_8.Po ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_9.G ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_9.G1 ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_9.Go ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_9.P ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_9.P1 ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_9.Po ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_4_10.G ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_4_10.G1 ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_4_10.Go ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_4_10.P ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_4_10.P1 ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_4_10.Po ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_4_11.G ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_4_11.G1 ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_4_11.Go ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_4_11.P ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_4_11.P1 ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_4_11.Po ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_4_12.G ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_4_12.G1 ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_4_12.Go ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_4_12.P ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_4_12.P1 ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_4_12.Po ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_4_13.G ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_4_13.G1 ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_4_13.Go ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_4_13.P ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_4_13.P1 ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_4_13.Po ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_4_14.G ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_4_14.G1 ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_4_14.Go ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_4_14.P ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_4_14.P1 ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_4_14.Po ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_4_15.G ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_4_15.G1 ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_4_15.Go ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_4_15.P ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_4_15.P1 ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_4_15.Po ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_4_8.G ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_4_8.G1 ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_4_8.Go ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_4_8.P ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_4_8.P1 ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_4_8.Po ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_4_9.G ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_4_9.G1 ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_4_9.Go ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_4_9.P ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_4_9.P1 ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_4_9.Po ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_1_0.G ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_1_0.Go ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_1_0.P ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_2_1.G1 ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_2_1.Go ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_2_1.P ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_3_2.G ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_3_2.G1 ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_3_2.Go ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_3_2.P ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_3_3.G ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_3_3.G1 ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_3_3.Go ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_3_3.P ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_4_4.G ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_4_4.G1 ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_4_4.Go ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_4_4.P ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_4_5.G ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_4_5.G1 ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_4_5.Go ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_4_5.P ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_4_6.G ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_4_6.G1 ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_4_6.Go ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_4_6.P ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_4_7.G ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_4_7.G1 ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_4_7.Go ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_4_7.P ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_5_10.G ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_5_10.G1 ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_5_10.Go ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_5_10.P ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_5_11.G ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_5_11.G1 ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_5_11.Go ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_5_11.P ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_5_12.G ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_5_12.G1 ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_5_12.Go ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_5_12.P ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_5_13.G ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_5_13.G1 ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_5_13.Go ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_5_13.P ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_5_14.G ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_5_14.G1 ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_5_14.Go ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_5_14.P ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_5_15.G ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_5_15.G1 ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_5_15.Go ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_5_15.P ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_5_8.G ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_5_8.G1 ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_5_8.Go ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_5_8.P ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_5_9.G ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_5_9.G1 ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_5_9.Go ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_5_9.P ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_6_0.G1 ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_6_0.Go ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_6_0.P ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_6_1.G ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_6_1.G1 ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_6_1.Go ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_6_1.P ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_6_10.G ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_6_10.G1 ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_6_10.Go ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_6_10.P ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_6_11.G ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_6_11.G1 ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_6_11.Go ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_6_11.P ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_6_12.G1 ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_6_12.Go ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_6_12.P ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_6_13.G1 ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_6_13.Go ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_6_13.P ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_6_14.G1 ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_6_14.Go ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_6_14.P ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_6_15.G1 ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_6_15.P ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_6_2.G ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_6_2.G1 ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_6_2.Go ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_6_2.P ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_6_3.G ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_6_3.G1 ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_6_3.Go ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_6_3.P ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_6_4.G ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_6_4.G1 ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_6_4.Go ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_6_4.P ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_6_5.G ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_6_5.G1 ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_6_5.Go ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_6_5.P ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_6_6.G ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_6_6.G1 ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_6_6.Go ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_6_6.P ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_6_7.G ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_6_7.G1 ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_6_7.Go ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_6_7.P ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_6_8.G ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_6_8.G1 ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_6_8.Go ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_6_8.P ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_6_9.G ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_6_9.G1 ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_6_9.Go ;
  wire \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_6_9.P ;
  wire \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_0.A ;
  wire \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_0.B ;
  wire [2:0] \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_0.codes ;
  wire \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_0.double ;
  wire \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_0.nA ;
  wire \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_0.nB ;
  wire \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_0.nBnC ;
  wire \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_0.negation ;
  wire \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_0.zero ;
  wire \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_1.A ;
  wire \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_1.B ;
  wire \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_1.BC ;
  wire \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_1.C ;
  wire [2:0] \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_1.codes ;
  wire \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_1.double ;
  wire \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_1.nA ;
  wire \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_1.nB ;
  wire \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_1.nBanC ;
  wire \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_1.nBnC ;
  wire \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_1.nC ;
  wire \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_1.negation ;
  wire \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_1.zero ;
  wire \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_2.A ;
  wire \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_2.B ;
  wire \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_2.BC ;
  wire \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_2.C ;
  wire [2:0] \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_2.codes ;
  wire \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_2.double ;
  wire \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_2.nA ;
  wire \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_2.nB ;
  wire \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_2.nBanC ;
  wire \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_2.nBnC ;
  wire \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_2.nC ;
  wire \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_2.negation ;
  wire \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_2.zero ;
  wire \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_3.A ;
  wire \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_3.B ;
  wire \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_3.BC ;
  wire \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_3.C ;
  wire [2:0] \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_3.codes ;
  wire \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_3.double ;
  wire \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_3.nA ;
  wire \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_3.nB ;
  wire \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_3.nBanC ;
  wire \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_3.nBnC ;
  wire \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_3.nC ;
  wire \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_3.negation ;
  wire \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_3.zero ;
  wire \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_4.A ;
  wire \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_4.B ;
  wire \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_4.BC ;
  wire \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_4.C ;
  wire [2:0] \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_4.codes ;
  wire \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_4.double ;
  wire \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_4.nA ;
  wire \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_4.nB ;
  wire \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_4.nBanC ;
  wire \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_4.nBnC ;
  wire \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_4.nC ;
  wire \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_4.negation ;
  wire \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_4.zero ;
  wire \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_5.A ;
  wire \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_5.B ;
  wire \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_5.BC ;
  wire \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_5.C ;
  wire [2:0] \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_5.codes ;
  wire \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_5.double ;
  wire \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_5.nA ;
  wire \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_5.nB ;
  wire \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_5.nBanC ;
  wire \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_5.nBnC ;
  wire \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_5.nC ;
  wire \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_5.negation ;
  wire \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_5.zero ;
  wire \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_6.A ;
  wire \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_6.B ;
  wire \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_6.BC ;
  wire \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_6.C ;
  wire [2:0] \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_6.codes ;
  wire \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_6.double ;
  wire \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_6.nA ;
  wire \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_6.nB ;
  wire \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_6.nBanC ;
  wire \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_6.nBnC ;
  wire \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_6.nC ;
  wire \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_6.negation ;
  wire \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_6.zero ;
  wire \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_7.A ;
  wire \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_7.B ;
  wire \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_7.BC ;
  wire \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_7.C ;
  wire [2:0] \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_7.codes ;
  wire \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_7.double ;
  wire \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_7.nA ;
  wire \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_7.nB ;
  wire \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_7.nBanC ;
  wire \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_7.nBnC ;
  wire \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_7.nC ;
  wire \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_7.negation ;
  wire \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_7.zero ;
  wire [7:0] \multiplier_16x16bit_pipelined.booth_array_0.double ;
  wire [15:0] \multiplier_16x16bit_pipelined.booth_array_0.multiplier ;
  wire [7:0] \multiplier_16x16bit_pipelined.booth_array_0.negation ;
  wire [7:0] \multiplier_16x16bit_pipelined.booth_array_0.zero ;
  wire [7:0] \multiplier_16x16bit_pipelined.double ;
  wire \multiplier_16x16bit_pipelined.i_clk ;
  wire [15:0] \multiplier_16x16bit_pipelined.i_md ;
  wire [15:0] \multiplier_16x16bit_pipelined.i_mr ;
  wire \multiplier_16x16bit_pipelined.i_rst ;
  wire \multiplier_16x16bit_pipelined.i_start ;
  wire \multiplier_16x16bit_pipelined.layer_0_w0[0] ;
  wire \multiplier_16x16bit_pipelined.layer_0_w0[1] ;
  wire \multiplier_16x16bit_pipelined.layer_0_w1 ;
  wire \multiplier_16x16bit_pipelined.layer_0_w10[0] ;
  wire \multiplier_16x16bit_pipelined.layer_0_w10[1] ;
  wire \multiplier_16x16bit_pipelined.layer_0_w10[2] ;
  wire \multiplier_16x16bit_pipelined.layer_0_w10[3] ;
  wire \multiplier_16x16bit_pipelined.layer_0_w10[4] ;
  wire \multiplier_16x16bit_pipelined.layer_0_w10[5] ;
  wire \multiplier_16x16bit_pipelined.layer_0_w10[6] ;
  wire \multiplier_16x16bit_pipelined.layer_0_w11[0] ;
  wire \multiplier_16x16bit_pipelined.layer_0_w11[1] ;
  wire \multiplier_16x16bit_pipelined.layer_0_w11[2] ;
  wire \multiplier_16x16bit_pipelined.layer_0_w11[3] ;
  wire \multiplier_16x16bit_pipelined.layer_0_w11[4] ;
  wire \multiplier_16x16bit_pipelined.layer_0_w11[5] ;
  wire \multiplier_16x16bit_pipelined.layer_0_w12[0] ;
  wire \multiplier_16x16bit_pipelined.layer_0_w12[1] ;
  wire \multiplier_16x16bit_pipelined.layer_0_w12[2] ;
  wire \multiplier_16x16bit_pipelined.layer_0_w12[3] ;
  wire \multiplier_16x16bit_pipelined.layer_0_w12[4] ;
  wire \multiplier_16x16bit_pipelined.layer_0_w12[5] ;
  wire \multiplier_16x16bit_pipelined.layer_0_w12[6] ;
  wire \multiplier_16x16bit_pipelined.layer_0_w12[7] ;
  wire \multiplier_16x16bit_pipelined.layer_0_w13[0] ;
  wire \multiplier_16x16bit_pipelined.layer_0_w13[1] ;
  wire \multiplier_16x16bit_pipelined.layer_0_w13[2] ;
  wire \multiplier_16x16bit_pipelined.layer_0_w13[3] ;
  wire \multiplier_16x16bit_pipelined.layer_0_w13[4] ;
  wire \multiplier_16x16bit_pipelined.layer_0_w13[5] ;
  wire \multiplier_16x16bit_pipelined.layer_0_w13[6] ;
  wire \multiplier_16x16bit_pipelined.layer_0_w14[0] ;
  wire \multiplier_16x16bit_pipelined.layer_0_w14[1] ;
  wire \multiplier_16x16bit_pipelined.layer_0_w14[2] ;
  wire \multiplier_16x16bit_pipelined.layer_0_w14[3] ;
  wire \multiplier_16x16bit_pipelined.layer_0_w14[4] ;
  wire \multiplier_16x16bit_pipelined.layer_0_w14[5] ;
  wire \multiplier_16x16bit_pipelined.layer_0_w14[6] ;
  wire \multiplier_16x16bit_pipelined.layer_0_w14[7] ;
  wire \multiplier_16x16bit_pipelined.layer_0_w14[8] ;
  wire \multiplier_16x16bit_pipelined.layer_0_w15[0] ;
  wire \multiplier_16x16bit_pipelined.layer_0_w15[1] ;
  wire \multiplier_16x16bit_pipelined.layer_0_w15[2] ;
  wire \multiplier_16x16bit_pipelined.layer_0_w15[3] ;
  wire \multiplier_16x16bit_pipelined.layer_0_w15[4] ;
  wire \multiplier_16x16bit_pipelined.layer_0_w15[5] ;
  wire \multiplier_16x16bit_pipelined.layer_0_w15[6] ;
  wire \multiplier_16x16bit_pipelined.layer_0_w15[7] ;
  wire \multiplier_16x16bit_pipelined.layer_0_w16[0] ;
  wire \multiplier_16x16bit_pipelined.layer_0_w16[1] ;
  wire \multiplier_16x16bit_pipelined.layer_0_w16[2] ;
  wire \multiplier_16x16bit_pipelined.layer_0_w16[3] ;
  wire \multiplier_16x16bit_pipelined.layer_0_w16[4] ;
  wire \multiplier_16x16bit_pipelined.layer_0_w16[5] ;
  wire \multiplier_16x16bit_pipelined.layer_0_w16[6] ;
  wire \multiplier_16x16bit_pipelined.layer_0_w16[7] ;
  wire \multiplier_16x16bit_pipelined.layer_0_w17[0] ;
  wire \multiplier_16x16bit_pipelined.layer_0_w17[1] ;
  wire \multiplier_16x16bit_pipelined.layer_0_w17[2] ;
  wire \multiplier_16x16bit_pipelined.layer_0_w17[3] ;
  wire \multiplier_16x16bit_pipelined.layer_0_w17[4] ;
  wire \multiplier_16x16bit_pipelined.layer_0_w17[5] ;
  wire \multiplier_16x16bit_pipelined.layer_0_w17[6] ;
  wire \multiplier_16x16bit_pipelined.layer_0_w18[0] ;
  wire \multiplier_16x16bit_pipelined.layer_0_w18[1] ;
  wire \multiplier_16x16bit_pipelined.layer_0_w18[2] ;
  wire \multiplier_16x16bit_pipelined.layer_0_w18[3] ;
  wire \multiplier_16x16bit_pipelined.layer_0_w18[4] ;
  wire \multiplier_16x16bit_pipelined.layer_0_w18[5] ;
  wire \multiplier_16x16bit_pipelined.layer_0_w18[6] ;
  wire \multiplier_16x16bit_pipelined.layer_0_w19[0] ;
  wire \multiplier_16x16bit_pipelined.layer_0_w19[1] ;
  wire \multiplier_16x16bit_pipelined.layer_0_w19[2] ;
  wire \multiplier_16x16bit_pipelined.layer_0_w19[3] ;
  wire \multiplier_16x16bit_pipelined.layer_0_w19[4] ;
  wire \multiplier_16x16bit_pipelined.layer_0_w19[5] ;
  wire \multiplier_16x16bit_pipelined.layer_0_w20[0] ;
  wire \multiplier_16x16bit_pipelined.layer_0_w20[1] ;
  wire \multiplier_16x16bit_pipelined.layer_0_w20[2] ;
  wire \multiplier_16x16bit_pipelined.layer_0_w20[3] ;
  wire \multiplier_16x16bit_pipelined.layer_0_w20[4] ;
  wire \multiplier_16x16bit_pipelined.layer_0_w20[5] ;
  wire \multiplier_16x16bit_pipelined.layer_0_w21[0] ;
  wire \multiplier_16x16bit_pipelined.layer_0_w21[1] ;
  wire \multiplier_16x16bit_pipelined.layer_0_w21[2] ;
  wire \multiplier_16x16bit_pipelined.layer_0_w21[3] ;
  wire \multiplier_16x16bit_pipelined.layer_0_w21[4] ;
  wire \multiplier_16x16bit_pipelined.layer_0_w22[0] ;
  wire \multiplier_16x16bit_pipelined.layer_0_w22[1] ;
  wire \multiplier_16x16bit_pipelined.layer_0_w22[2] ;
  wire \multiplier_16x16bit_pipelined.layer_0_w22[3] ;
  wire \multiplier_16x16bit_pipelined.layer_0_w22[4] ;
  wire \multiplier_16x16bit_pipelined.layer_0_w23[0] ;
  wire \multiplier_16x16bit_pipelined.layer_0_w23[1] ;
  wire \multiplier_16x16bit_pipelined.layer_0_w23[2] ;
  wire \multiplier_16x16bit_pipelined.layer_0_w23[3] ;
  wire \multiplier_16x16bit_pipelined.layer_0_w24[0] ;
  wire \multiplier_16x16bit_pipelined.layer_0_w24[1] ;
  wire \multiplier_16x16bit_pipelined.layer_0_w24[2] ;
  wire \multiplier_16x16bit_pipelined.layer_0_w24[3] ;
  wire \multiplier_16x16bit_pipelined.layer_0_w25[0] ;
  wire \multiplier_16x16bit_pipelined.layer_0_w25[1] ;
  wire \multiplier_16x16bit_pipelined.layer_0_w25[2] ;
  wire \multiplier_16x16bit_pipelined.layer_0_w26[0] ;
  wire \multiplier_16x16bit_pipelined.layer_0_w26[1] ;
  wire \multiplier_16x16bit_pipelined.layer_0_w26[2] ;
  wire \multiplier_16x16bit_pipelined.layer_0_w27[0] ;
  wire \multiplier_16x16bit_pipelined.layer_0_w27[1] ;
  wire \multiplier_16x16bit_pipelined.layer_0_w28[0] ;
  wire \multiplier_16x16bit_pipelined.layer_0_w28[1] ;
  wire \multiplier_16x16bit_pipelined.layer_0_w29[0] ;
  wire \multiplier_16x16bit_pipelined.layer_0_w2[0] ;
  wire \multiplier_16x16bit_pipelined.layer_0_w2[1] ;
  wire \multiplier_16x16bit_pipelined.layer_0_w2[2] ;
  wire \multiplier_16x16bit_pipelined.layer_0_w30 ;
  wire \multiplier_16x16bit_pipelined.layer_0_w3[0] ;
  wire \multiplier_16x16bit_pipelined.layer_0_w3[1] ;
  wire \multiplier_16x16bit_pipelined.layer_0_w4[0] ;
  wire \multiplier_16x16bit_pipelined.layer_0_w4[1] ;
  wire \multiplier_16x16bit_pipelined.layer_0_w4[2] ;
  wire \multiplier_16x16bit_pipelined.layer_0_w4[3] ;
  wire \multiplier_16x16bit_pipelined.layer_0_w5[0] ;
  wire \multiplier_16x16bit_pipelined.layer_0_w5[1] ;
  wire \multiplier_16x16bit_pipelined.layer_0_w5[2] ;
  wire \multiplier_16x16bit_pipelined.layer_0_w6[0] ;
  wire \multiplier_16x16bit_pipelined.layer_0_w6[1] ;
  wire \multiplier_16x16bit_pipelined.layer_0_w6[2] ;
  wire \multiplier_16x16bit_pipelined.layer_0_w6[3] ;
  wire \multiplier_16x16bit_pipelined.layer_0_w6[4] ;
  wire \multiplier_16x16bit_pipelined.layer_0_w7[0] ;
  wire \multiplier_16x16bit_pipelined.layer_0_w7[1] ;
  wire \multiplier_16x16bit_pipelined.layer_0_w7[2] ;
  wire \multiplier_16x16bit_pipelined.layer_0_w7[3] ;
  wire \multiplier_16x16bit_pipelined.layer_0_w8[0] ;
  wire \multiplier_16x16bit_pipelined.layer_0_w8[1] ;
  wire \multiplier_16x16bit_pipelined.layer_0_w8[2] ;
  wire \multiplier_16x16bit_pipelined.layer_0_w8[3] ;
  wire \multiplier_16x16bit_pipelined.layer_0_w8[4] ;
  wire \multiplier_16x16bit_pipelined.layer_0_w8[5] ;
  wire \multiplier_16x16bit_pipelined.layer_0_w9[0] ;
  wire \multiplier_16x16bit_pipelined.layer_0_w9[1] ;
  wire \multiplier_16x16bit_pipelined.layer_0_w9[2] ;
  wire \multiplier_16x16bit_pipelined.layer_0_w9[3] ;
  wire \multiplier_16x16bit_pipelined.layer_0_w9[4] ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_0.A ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_0.AB ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_0.AxBxCxD ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_0.AxorB ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_0.B ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_0.C ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_0.CD ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_0.CxorD ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_0.D ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_0.S ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_0.carry ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_0.cin ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_0.cout ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_1.A ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_1.AB ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_1.AxBxCxD ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_1.AxorB ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_1.B ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_1.C ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_1.CD ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_1.CxorD ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_1.D ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_1.S ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_1.carry ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_1.cin ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_1.cout ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_10.A ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_10.AB ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_10.AxBxCxD ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_10.AxorB ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_10.B ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_10.C ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_10.CD ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_10.CxorD ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_10.D ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_10.S ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_10.carry ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_10.cin ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_10.cout ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_11.A ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_11.AB ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_11.AxBxCxD ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_11.AxorB ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_11.B ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_11.C ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_11.CD ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_11.CxorD ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_11.D ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_11.S ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_11.carry ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_11.cin ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_11.cout ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_12.A ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_12.AB ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_12.AxBxCxD ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_12.AxorB ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_12.B ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_12.C ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_12.CD ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_12.CxorD ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_12.D ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_12.S ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_12.carry ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_12.cin ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_12.cout ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_13.A ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_13.AB ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_13.AxBxCxD ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_13.AxorB ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_13.B ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_13.C ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_13.CD ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_13.CxorD ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_13.D ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_13.S ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_13.carry ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_13.cin ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_13.cout ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_14.A ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_14.AB ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_14.AxBxCxD ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_14.AxorB ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_14.B ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_14.C ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_14.CD ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_14.CxorD ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_14.D ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_14.S ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_14.carry ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_14.cin ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_14.cout ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_15.A ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_15.AB ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_15.AxBxCxD ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_15.AxorB ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_15.B ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_15.C ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_15.CD ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_15.CxorD ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_15.D ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_15.S ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_15.carry ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_15.cin ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_15.cout ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_16.A ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_16.AB ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_16.AxBxCxD ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_16.AxorB ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_16.B ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_16.C ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_16.CD ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_16.CxorD ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_16.D ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_16.S ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_16.carry ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_16.cout ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_2.A ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_2.AB ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_2.AxBxCxD ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_2.AxorB ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_2.B ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_2.C ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_2.CD ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_2.CxorD ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_2.D ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_2.S ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_2.carry ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_2.cin ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_2.cout ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_3.A ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_3.AB ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_3.AxBxCxD ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_3.AxorB ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_3.B ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_3.C ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_3.CD ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_3.CxorD ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_3.D ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_3.S ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_3.carry ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_3.cin ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_3.cout ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_4.A ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_4.AB ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_4.AxBxCxD ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_4.AxorB ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_4.B ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_4.C ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_4.CD ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_4.CxorD ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_4.D ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_4.S ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_4.carry ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_4.cin ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_4.cout ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_5.A ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_5.AB ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_5.AxBxCxD ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_5.AxorB ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_5.B ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_5.C ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_5.CD ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_5.CxorD ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_5.D ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_5.S ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_5.carry ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_5.cin ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_5.cout ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_6.A ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_6.AB ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_6.AxBxCxD ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_6.AxorB ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_6.B ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_6.C ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_6.CD ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_6.CxorD ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_6.D ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_6.S ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_6.carry ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_6.cin ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_6.cout ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_7.A ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_7.AB ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_7.AxBxCxD ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_7.AxorB ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_7.B ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_7.C ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_7.CD ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_7.CxorD ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_7.D ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_7.S ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_7.carry ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_7.cin ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_7.cout ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_8.A ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_8.AB ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_8.AxBxCxD ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_8.AxorB ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_8.B ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_8.C ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_8.CD ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_8.CxorD ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_8.D ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_8.S ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_8.carry ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_8.cin ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_8.cout ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_9.A ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_9.AB ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_9.AxBxCxD ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_9.AxorB ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_9.B ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_9.C ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_9.CD ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_9.CxorD ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_9.D ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_9.S ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_9.carry ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_9.cin ;
  wire \multiplier_16x16bit_pipelined.layer_1_compressor42_9.cout ;
  wire \multiplier_16x16bit_pipelined.layer_1_full_adder_0.A ;
  wire \multiplier_16x16bit_pipelined.layer_1_full_adder_0.AB ;
  wire \multiplier_16x16bit_pipelined.layer_1_full_adder_0.AxorB ;
  wire \multiplier_16x16bit_pipelined.layer_1_full_adder_0.B ;
  wire \multiplier_16x16bit_pipelined.layer_1_full_adder_0.S ;
  wire \multiplier_16x16bit_pipelined.layer_1_full_adder_0.cin ;
  wire \multiplier_16x16bit_pipelined.layer_1_full_adder_0.cout ;
  wire \multiplier_16x16bit_pipelined.layer_1_full_adder_1.A ;
  wire \multiplier_16x16bit_pipelined.layer_1_full_adder_1.AB ;
  wire \multiplier_16x16bit_pipelined.layer_1_full_adder_1.AxorB ;
  wire \multiplier_16x16bit_pipelined.layer_1_full_adder_1.B ;
  wire \multiplier_16x16bit_pipelined.layer_1_full_adder_1.S ;
  wire \multiplier_16x16bit_pipelined.layer_1_full_adder_1.cin ;
  wire \multiplier_16x16bit_pipelined.layer_1_full_adder_1.cout ;
  wire \multiplier_16x16bit_pipelined.layer_1_full_adder_10.A ;
  wire \multiplier_16x16bit_pipelined.layer_1_full_adder_10.AB ;
  wire \multiplier_16x16bit_pipelined.layer_1_full_adder_10.AxorB ;
  wire \multiplier_16x16bit_pipelined.layer_1_full_adder_10.B ;
  wire \multiplier_16x16bit_pipelined.layer_1_full_adder_10.S ;
  wire \multiplier_16x16bit_pipelined.layer_1_full_adder_10.cin ;
  wire \multiplier_16x16bit_pipelined.layer_1_full_adder_10.cout ;
  wire \multiplier_16x16bit_pipelined.layer_1_full_adder_11.A ;
  wire \multiplier_16x16bit_pipelined.layer_1_full_adder_11.AB ;
  wire \multiplier_16x16bit_pipelined.layer_1_full_adder_11.AxorB ;
  wire \multiplier_16x16bit_pipelined.layer_1_full_adder_11.B ;
  wire \multiplier_16x16bit_pipelined.layer_1_full_adder_11.S ;
  wire \multiplier_16x16bit_pipelined.layer_1_full_adder_11.cout ;
  wire \multiplier_16x16bit_pipelined.layer_1_full_adder_2.A ;
  wire \multiplier_16x16bit_pipelined.layer_1_full_adder_2.AB ;
  wire \multiplier_16x16bit_pipelined.layer_1_full_adder_2.AxorB ;
  wire \multiplier_16x16bit_pipelined.layer_1_full_adder_2.B ;
  wire \multiplier_16x16bit_pipelined.layer_1_full_adder_2.S ;
  wire \multiplier_16x16bit_pipelined.layer_1_full_adder_2.cin ;
  wire \multiplier_16x16bit_pipelined.layer_1_full_adder_2.cout ;
  wire \multiplier_16x16bit_pipelined.layer_1_full_adder_3.A ;
  wire \multiplier_16x16bit_pipelined.layer_1_full_adder_3.AB ;
  wire \multiplier_16x16bit_pipelined.layer_1_full_adder_3.AxorB ;
  wire \multiplier_16x16bit_pipelined.layer_1_full_adder_3.B ;
  wire \multiplier_16x16bit_pipelined.layer_1_full_adder_3.S ;
  wire \multiplier_16x16bit_pipelined.layer_1_full_adder_3.cin ;
  wire \multiplier_16x16bit_pipelined.layer_1_full_adder_3.cout ;
  wire \multiplier_16x16bit_pipelined.layer_1_full_adder_4.A ;
  wire \multiplier_16x16bit_pipelined.layer_1_full_adder_4.AB ;
  wire \multiplier_16x16bit_pipelined.layer_1_full_adder_4.AxorB ;
  wire \multiplier_16x16bit_pipelined.layer_1_full_adder_4.B ;
  wire \multiplier_16x16bit_pipelined.layer_1_full_adder_4.S ;
  wire \multiplier_16x16bit_pipelined.layer_1_full_adder_4.cin ;
  wire \multiplier_16x16bit_pipelined.layer_1_full_adder_4.cout ;
  wire \multiplier_16x16bit_pipelined.layer_1_full_adder_5.A ;
  wire \multiplier_16x16bit_pipelined.layer_1_full_adder_5.AB ;
  wire \multiplier_16x16bit_pipelined.layer_1_full_adder_5.AxorB ;
  wire \multiplier_16x16bit_pipelined.layer_1_full_adder_5.B ;
  wire \multiplier_16x16bit_pipelined.layer_1_full_adder_5.S ;
  wire \multiplier_16x16bit_pipelined.layer_1_full_adder_5.cin ;
  wire \multiplier_16x16bit_pipelined.layer_1_full_adder_5.cout ;
  wire \multiplier_16x16bit_pipelined.layer_1_full_adder_6.A ;
  wire \multiplier_16x16bit_pipelined.layer_1_full_adder_6.AB ;
  wire \multiplier_16x16bit_pipelined.layer_1_full_adder_6.AxorB ;
  wire \multiplier_16x16bit_pipelined.layer_1_full_adder_6.B ;
  wire \multiplier_16x16bit_pipelined.layer_1_full_adder_6.S ;
  wire \multiplier_16x16bit_pipelined.layer_1_full_adder_6.cin ;
  wire \multiplier_16x16bit_pipelined.layer_1_full_adder_6.cout ;
  wire \multiplier_16x16bit_pipelined.layer_1_full_adder_7.A ;
  wire \multiplier_16x16bit_pipelined.layer_1_full_adder_7.AB ;
  wire \multiplier_16x16bit_pipelined.layer_1_full_adder_7.AxorB ;
  wire \multiplier_16x16bit_pipelined.layer_1_full_adder_7.B ;
  wire \multiplier_16x16bit_pipelined.layer_1_full_adder_7.S ;
  wire \multiplier_16x16bit_pipelined.layer_1_full_adder_7.cout ;
  wire \multiplier_16x16bit_pipelined.layer_1_full_adder_8.A ;
  wire \multiplier_16x16bit_pipelined.layer_1_full_adder_8.AB ;
  wire \multiplier_16x16bit_pipelined.layer_1_full_adder_8.AxorB ;
  wire \multiplier_16x16bit_pipelined.layer_1_full_adder_8.B ;
  wire \multiplier_16x16bit_pipelined.layer_1_full_adder_8.S ;
  wire \multiplier_16x16bit_pipelined.layer_1_full_adder_8.cin ;
  wire \multiplier_16x16bit_pipelined.layer_1_full_adder_8.cout ;
  wire \multiplier_16x16bit_pipelined.layer_1_full_adder_9.A ;
  wire \multiplier_16x16bit_pipelined.layer_1_full_adder_9.AB ;
  wire \multiplier_16x16bit_pipelined.layer_1_full_adder_9.AxorB ;
  wire \multiplier_16x16bit_pipelined.layer_1_full_adder_9.B ;
  wire \multiplier_16x16bit_pipelined.layer_1_full_adder_9.S ;
  wire \multiplier_16x16bit_pipelined.layer_1_full_adder_9.cin ;
  wire \multiplier_16x16bit_pipelined.layer_1_full_adder_9.cout ;
  wire \multiplier_16x16bit_pipelined.layer_1_w0[0] ;
  wire \multiplier_16x16bit_pipelined.layer_1_w0[1] ;
  wire \multiplier_16x16bit_pipelined.layer_1_w1 ;
  wire \multiplier_16x16bit_pipelined.layer_1_w10[0] ;
  wire \multiplier_16x16bit_pipelined.layer_1_w10[1] ;
  wire \multiplier_16x16bit_pipelined.layer_1_w10[2] ;
  wire \multiplier_16x16bit_pipelined.layer_1_w10[3] ;
  wire \multiplier_16x16bit_pipelined.layer_1_w10[4] ;
  wire \multiplier_16x16bit_pipelined.layer_1_w11[0] ;
  wire \multiplier_16x16bit_pipelined.layer_1_w11[1] ;
  wire \multiplier_16x16bit_pipelined.layer_1_w11[2] ;
  wire \multiplier_16x16bit_pipelined.layer_1_w11[3] ;
  wire \multiplier_16x16bit_pipelined.layer_1_w12[0] ;
  wire \multiplier_16x16bit_pipelined.layer_1_w12[1] ;
  wire \multiplier_16x16bit_pipelined.layer_1_w12[2] ;
  wire \multiplier_16x16bit_pipelined.layer_1_w12[3] ;
  wire \multiplier_16x16bit_pipelined.layer_1_w13[0] ;
  wire \multiplier_16x16bit_pipelined.layer_1_w13[1] ;
  wire \multiplier_16x16bit_pipelined.layer_1_w13[2] ;
  wire \multiplier_16x16bit_pipelined.layer_1_w13[3] ;
  wire \multiplier_16x16bit_pipelined.layer_1_w13[4] ;
  wire \multiplier_16x16bit_pipelined.layer_1_w13[5] ;
  wire \multiplier_16x16bit_pipelined.layer_1_w14[0] ;
  wire \multiplier_16x16bit_pipelined.layer_1_w14[1] ;
  wire \multiplier_16x16bit_pipelined.layer_1_w14[2] ;
  wire \multiplier_16x16bit_pipelined.layer_1_w14[3] ;
  wire \multiplier_16x16bit_pipelined.layer_1_w14[4] ;
  wire \multiplier_16x16bit_pipelined.layer_1_w15[0] ;
  wire \multiplier_16x16bit_pipelined.layer_1_w15[1] ;
  wire \multiplier_16x16bit_pipelined.layer_1_w15[2] ;
  wire \multiplier_16x16bit_pipelined.layer_1_w15[3] ;
  wire \multiplier_16x16bit_pipelined.layer_1_w15[4] ;
  wire \multiplier_16x16bit_pipelined.layer_1_w16[0] ;
  wire \multiplier_16x16bit_pipelined.layer_1_w16[1] ;
  wire \multiplier_16x16bit_pipelined.layer_1_w16[2] ;
  wire \multiplier_16x16bit_pipelined.layer_1_w16[3] ;
  wire \multiplier_16x16bit_pipelined.layer_1_w16[4] ;
  wire \multiplier_16x16bit_pipelined.layer_1_w17[0] ;
  wire \multiplier_16x16bit_pipelined.layer_1_w17[1] ;
  wire \multiplier_16x16bit_pipelined.layer_1_w17[2] ;
  wire \multiplier_16x16bit_pipelined.layer_1_w17[3] ;
  wire \multiplier_16x16bit_pipelined.layer_1_w17[4] ;
  wire \multiplier_16x16bit_pipelined.layer_1_w18[0] ;
  wire \multiplier_16x16bit_pipelined.layer_1_w18[1] ;
  wire \multiplier_16x16bit_pipelined.layer_1_w18[2] ;
  wire \multiplier_16x16bit_pipelined.layer_1_w18[3] ;
  wire \multiplier_16x16bit_pipelined.layer_1_w18[4] ;
  wire \multiplier_16x16bit_pipelined.layer_1_w18[5] ;
  wire \multiplier_16x16bit_pipelined.layer_1_w19[0] ;
  wire \multiplier_16x16bit_pipelined.layer_1_w19[1] ;
  wire \multiplier_16x16bit_pipelined.layer_1_w19[2] ;
  wire \multiplier_16x16bit_pipelined.layer_1_w19[3] ;
  wire \multiplier_16x16bit_pipelined.layer_1_w20[0] ;
  wire \multiplier_16x16bit_pipelined.layer_1_w20[1] ;
  wire \multiplier_16x16bit_pipelined.layer_1_w20[2] ;
  wire \multiplier_16x16bit_pipelined.layer_1_w20[3] ;
  wire \multiplier_16x16bit_pipelined.layer_1_w21[0] ;
  wire \multiplier_16x16bit_pipelined.layer_1_w21[1] ;
  wire \multiplier_16x16bit_pipelined.layer_1_w21[2] ;
  wire \multiplier_16x16bit_pipelined.layer_1_w22[0] ;
  wire \multiplier_16x16bit_pipelined.layer_1_w22[1] ;
  wire \multiplier_16x16bit_pipelined.layer_1_w22[2] ;
  wire \multiplier_16x16bit_pipelined.layer_1_w23[0] ;
  wire \multiplier_16x16bit_pipelined.layer_1_w23[1] ;
  wire \multiplier_16x16bit_pipelined.layer_1_w23[2] ;
  wire \multiplier_16x16bit_pipelined.layer_1_w24[0] ;
  wire \multiplier_16x16bit_pipelined.layer_1_w24[1] ;
  wire \multiplier_16x16bit_pipelined.layer_1_w24[2] ;
  wire \multiplier_16x16bit_pipelined.layer_1_w24[3] ;
  wire \multiplier_16x16bit_pipelined.layer_1_w25[0] ;
  wire \multiplier_16x16bit_pipelined.layer_1_w25[1] ;
  wire \multiplier_16x16bit_pipelined.layer_1_w26[0] ;
  wire \multiplier_16x16bit_pipelined.layer_1_w26[1] ;
  wire \multiplier_16x16bit_pipelined.layer_1_w27[0] ;
  wire \multiplier_16x16bit_pipelined.layer_1_w27[1] ;
  wire \multiplier_16x16bit_pipelined.layer_1_w28[0] ;
  wire \multiplier_16x16bit_pipelined.layer_1_w28[1] ;
  wire \multiplier_16x16bit_pipelined.layer_1_w28[2] ;
  wire \multiplier_16x16bit_pipelined.layer_1_w29[0] ;
  wire \multiplier_16x16bit_pipelined.layer_1_w2[0] ;
  wire \multiplier_16x16bit_pipelined.layer_1_w2[1] ;
  wire \multiplier_16x16bit_pipelined.layer_1_w2[2] ;
  wire \multiplier_16x16bit_pipelined.layer_1_w30 ;
  wire \multiplier_16x16bit_pipelined.layer_1_w3[0] ;
  wire \multiplier_16x16bit_pipelined.layer_1_w3[1] ;
  wire \multiplier_16x16bit_pipelined.layer_1_w4[0] ;
  wire \multiplier_16x16bit_pipelined.layer_1_w4[1] ;
  wire \multiplier_16x16bit_pipelined.layer_1_w5[0] ;
  wire \multiplier_16x16bit_pipelined.layer_1_w5[1] ;
  wire \multiplier_16x16bit_pipelined.layer_1_w6[0] ;
  wire \multiplier_16x16bit_pipelined.layer_1_w6[1] ;
  wire \multiplier_16x16bit_pipelined.layer_1_w7[0] ;
  wire \multiplier_16x16bit_pipelined.layer_1_w7[1] ;
  wire \multiplier_16x16bit_pipelined.layer_1_w7[2] ;
  wire \multiplier_16x16bit_pipelined.layer_1_w7[3] ;
  wire \multiplier_16x16bit_pipelined.layer_1_w8[0] ;
  wire \multiplier_16x16bit_pipelined.layer_1_w8[1] ;
  wire \multiplier_16x16bit_pipelined.layer_1_w8[2] ;
  wire \multiplier_16x16bit_pipelined.layer_1_w9[0] ;
  wire \multiplier_16x16bit_pipelined.layer_1_w9[1] ;
  wire \multiplier_16x16bit_pipelined.layer_1_w9[2] ;
  wire \multiplier_16x16bit_pipelined.layer_2_compressor42_0.A ;
  wire \multiplier_16x16bit_pipelined.layer_2_compressor42_0.AB ;
  wire \multiplier_16x16bit_pipelined.layer_2_compressor42_0.AxBxCxD ;
  wire \multiplier_16x16bit_pipelined.layer_2_compressor42_0.AxorB ;
  wire \multiplier_16x16bit_pipelined.layer_2_compressor42_0.B ;
  wire \multiplier_16x16bit_pipelined.layer_2_compressor42_0.C ;
  wire \multiplier_16x16bit_pipelined.layer_2_compressor42_0.CD ;
  wire \multiplier_16x16bit_pipelined.layer_2_compressor42_0.CxorD ;
  wire \multiplier_16x16bit_pipelined.layer_2_compressor42_0.D ;
  wire \multiplier_16x16bit_pipelined.layer_2_compressor42_0.S ;
  wire \multiplier_16x16bit_pipelined.layer_2_compressor42_0.carry ;
  wire \multiplier_16x16bit_pipelined.layer_2_compressor42_0.cin ;
  wire \multiplier_16x16bit_pipelined.layer_2_compressor42_0.cout ;
  wire \multiplier_16x16bit_pipelined.layer_2_compressor42_1.A ;
  wire \multiplier_16x16bit_pipelined.layer_2_compressor42_1.AB ;
  wire \multiplier_16x16bit_pipelined.layer_2_compressor42_1.AxBxCxD ;
  wire \multiplier_16x16bit_pipelined.layer_2_compressor42_1.AxorB ;
  wire \multiplier_16x16bit_pipelined.layer_2_compressor42_1.B ;
  wire \multiplier_16x16bit_pipelined.layer_2_compressor42_1.C ;
  wire \multiplier_16x16bit_pipelined.layer_2_compressor42_1.CD ;
  wire \multiplier_16x16bit_pipelined.layer_2_compressor42_1.CxorD ;
  wire \multiplier_16x16bit_pipelined.layer_2_compressor42_1.D ;
  wire \multiplier_16x16bit_pipelined.layer_2_compressor42_1.S ;
  wire \multiplier_16x16bit_pipelined.layer_2_compressor42_1.carry ;
  wire \multiplier_16x16bit_pipelined.layer_2_compressor42_1.cin ;
  wire \multiplier_16x16bit_pipelined.layer_2_compressor42_1.cout ;
  wire \multiplier_16x16bit_pipelined.layer_2_compressor42_2.A ;
  wire \multiplier_16x16bit_pipelined.layer_2_compressor42_2.AB ;
  wire \multiplier_16x16bit_pipelined.layer_2_compressor42_2.AxBxCxD ;
  wire \multiplier_16x16bit_pipelined.layer_2_compressor42_2.AxorB ;
  wire \multiplier_16x16bit_pipelined.layer_2_compressor42_2.B ;
  wire \multiplier_16x16bit_pipelined.layer_2_compressor42_2.C ;
  wire \multiplier_16x16bit_pipelined.layer_2_compressor42_2.CD ;
  wire \multiplier_16x16bit_pipelined.layer_2_compressor42_2.CxorD ;
  wire \multiplier_16x16bit_pipelined.layer_2_compressor42_2.D ;
  wire \multiplier_16x16bit_pipelined.layer_2_compressor42_2.S ;
  wire \multiplier_16x16bit_pipelined.layer_2_compressor42_2.carry ;
  wire \multiplier_16x16bit_pipelined.layer_2_compressor42_2.cin ;
  wire \multiplier_16x16bit_pipelined.layer_2_compressor42_2.cout ;
  wire \multiplier_16x16bit_pipelined.layer_2_compressor42_3.A ;
  wire \multiplier_16x16bit_pipelined.layer_2_compressor42_3.AB ;
  wire \multiplier_16x16bit_pipelined.layer_2_compressor42_3.AxBxCxD ;
  wire \multiplier_16x16bit_pipelined.layer_2_compressor42_3.AxorB ;
  wire \multiplier_16x16bit_pipelined.layer_2_compressor42_3.B ;
  wire \multiplier_16x16bit_pipelined.layer_2_compressor42_3.C ;
  wire \multiplier_16x16bit_pipelined.layer_2_compressor42_3.CD ;
  wire \multiplier_16x16bit_pipelined.layer_2_compressor42_3.CxorD ;
  wire \multiplier_16x16bit_pipelined.layer_2_compressor42_3.D ;
  wire \multiplier_16x16bit_pipelined.layer_2_compressor42_3.S ;
  wire \multiplier_16x16bit_pipelined.layer_2_compressor42_3.carry ;
  wire \multiplier_16x16bit_pipelined.layer_2_compressor42_3.cin ;
  wire \multiplier_16x16bit_pipelined.layer_2_compressor42_3.cout ;
  wire \multiplier_16x16bit_pipelined.layer_2_compressor42_4.A ;
  wire \multiplier_16x16bit_pipelined.layer_2_compressor42_4.AB ;
  wire \multiplier_16x16bit_pipelined.layer_2_compressor42_4.AxBxCxD ;
  wire \multiplier_16x16bit_pipelined.layer_2_compressor42_4.AxorB ;
  wire \multiplier_16x16bit_pipelined.layer_2_compressor42_4.B ;
  wire \multiplier_16x16bit_pipelined.layer_2_compressor42_4.C ;
  wire \multiplier_16x16bit_pipelined.layer_2_compressor42_4.CD ;
  wire \multiplier_16x16bit_pipelined.layer_2_compressor42_4.CxorD ;
  wire \multiplier_16x16bit_pipelined.layer_2_compressor42_4.D ;
  wire \multiplier_16x16bit_pipelined.layer_2_compressor42_4.S ;
  wire \multiplier_16x16bit_pipelined.layer_2_compressor42_4.carry ;
  wire \multiplier_16x16bit_pipelined.layer_2_compressor42_4.cin ;
  wire \multiplier_16x16bit_pipelined.layer_2_compressor42_4.cout ;
  wire \multiplier_16x16bit_pipelined.layer_2_compressor42_5.A ;
  wire \multiplier_16x16bit_pipelined.layer_2_compressor42_5.AB ;
  wire \multiplier_16x16bit_pipelined.layer_2_compressor42_5.AxBxCxD ;
  wire \multiplier_16x16bit_pipelined.layer_2_compressor42_5.AxorB ;
  wire \multiplier_16x16bit_pipelined.layer_2_compressor42_5.B ;
  wire \multiplier_16x16bit_pipelined.layer_2_compressor42_5.C ;
  wire \multiplier_16x16bit_pipelined.layer_2_compressor42_5.CD ;
  wire \multiplier_16x16bit_pipelined.layer_2_compressor42_5.CxorD ;
  wire \multiplier_16x16bit_pipelined.layer_2_compressor42_5.D ;
  wire \multiplier_16x16bit_pipelined.layer_2_compressor42_5.S ;
  wire \multiplier_16x16bit_pipelined.layer_2_compressor42_5.carry ;
  wire \multiplier_16x16bit_pipelined.layer_2_compressor42_5.cin ;
  wire \multiplier_16x16bit_pipelined.layer_2_compressor42_5.cout ;
  wire \multiplier_16x16bit_pipelined.layer_2_compressor42_6.A ;
  wire \multiplier_16x16bit_pipelined.layer_2_compressor42_6.AB ;
  wire \multiplier_16x16bit_pipelined.layer_2_compressor42_6.AxBxCxD ;
  wire \multiplier_16x16bit_pipelined.layer_2_compressor42_6.AxorB ;
  wire \multiplier_16x16bit_pipelined.layer_2_compressor42_6.B ;
  wire \multiplier_16x16bit_pipelined.layer_2_compressor42_6.C ;
  wire \multiplier_16x16bit_pipelined.layer_2_compressor42_6.CD ;
  wire \multiplier_16x16bit_pipelined.layer_2_compressor42_6.CxorD ;
  wire \multiplier_16x16bit_pipelined.layer_2_compressor42_6.D ;
  wire \multiplier_16x16bit_pipelined.layer_2_compressor42_6.S ;
  wire \multiplier_16x16bit_pipelined.layer_2_compressor42_6.carry ;
  wire \multiplier_16x16bit_pipelined.layer_2_compressor42_6.cin ;
  wire \multiplier_16x16bit_pipelined.layer_2_compressor42_6.cout ;
  wire \multiplier_16x16bit_pipelined.layer_2_compressor42_7.A ;
  wire \multiplier_16x16bit_pipelined.layer_2_compressor42_7.AB ;
  wire \multiplier_16x16bit_pipelined.layer_2_compressor42_7.AxBxCxD ;
  wire \multiplier_16x16bit_pipelined.layer_2_compressor42_7.AxorB ;
  wire \multiplier_16x16bit_pipelined.layer_2_compressor42_7.B ;
  wire \multiplier_16x16bit_pipelined.layer_2_compressor42_7.C ;
  wire \multiplier_16x16bit_pipelined.layer_2_compressor42_7.CD ;
  wire \multiplier_16x16bit_pipelined.layer_2_compressor42_7.CxorD ;
  wire \multiplier_16x16bit_pipelined.layer_2_compressor42_7.D ;
  wire \multiplier_16x16bit_pipelined.layer_2_compressor42_7.S ;
  wire \multiplier_16x16bit_pipelined.layer_2_compressor42_7.carry ;
  wire \multiplier_16x16bit_pipelined.layer_2_compressor42_7.cout ;
  wire \multiplier_16x16bit_pipelined.layer_2_full_adder_0.A ;
  wire \multiplier_16x16bit_pipelined.layer_2_full_adder_0.AB ;
  wire \multiplier_16x16bit_pipelined.layer_2_full_adder_0.AxorB ;
  wire \multiplier_16x16bit_pipelined.layer_2_full_adder_0.B ;
  wire \multiplier_16x16bit_pipelined.layer_2_full_adder_0.S ;
  wire \multiplier_16x16bit_pipelined.layer_2_full_adder_0.cin ;
  wire \multiplier_16x16bit_pipelined.layer_2_full_adder_0.cout ;
  wire \multiplier_16x16bit_pipelined.layer_2_full_adder_1.A ;
  wire \multiplier_16x16bit_pipelined.layer_2_full_adder_1.AB ;
  wire \multiplier_16x16bit_pipelined.layer_2_full_adder_1.AxorB ;
  wire \multiplier_16x16bit_pipelined.layer_2_full_adder_1.B ;
  wire \multiplier_16x16bit_pipelined.layer_2_full_adder_1.S ;
  wire \multiplier_16x16bit_pipelined.layer_2_full_adder_1.cin ;
  wire \multiplier_16x16bit_pipelined.layer_2_full_adder_1.cout ;
  wire \multiplier_16x16bit_pipelined.layer_2_full_adder_10.A ;
  wire \multiplier_16x16bit_pipelined.layer_2_full_adder_10.AB ;
  wire \multiplier_16x16bit_pipelined.layer_2_full_adder_10.AxorB ;
  wire \multiplier_16x16bit_pipelined.layer_2_full_adder_10.B ;
  wire \multiplier_16x16bit_pipelined.layer_2_full_adder_10.S ;
  wire \multiplier_16x16bit_pipelined.layer_2_full_adder_10.cout ;
  wire \multiplier_16x16bit_pipelined.layer_2_full_adder_11.A ;
  wire \multiplier_16x16bit_pipelined.layer_2_full_adder_11.AB ;
  wire \multiplier_16x16bit_pipelined.layer_2_full_adder_11.AxorB ;
  wire \multiplier_16x16bit_pipelined.layer_2_full_adder_11.B ;
  wire \multiplier_16x16bit_pipelined.layer_2_full_adder_11.S ;
  wire \multiplier_16x16bit_pipelined.layer_2_full_adder_11.cin ;
  wire \multiplier_16x16bit_pipelined.layer_2_full_adder_11.cout ;
  wire \multiplier_16x16bit_pipelined.layer_2_full_adder_2.A ;
  wire \multiplier_16x16bit_pipelined.layer_2_full_adder_2.AB ;
  wire \multiplier_16x16bit_pipelined.layer_2_full_adder_2.AxorB ;
  wire \multiplier_16x16bit_pipelined.layer_2_full_adder_2.B ;
  wire \multiplier_16x16bit_pipelined.layer_2_full_adder_2.S ;
  wire \multiplier_16x16bit_pipelined.layer_2_full_adder_2.cin ;
  wire \multiplier_16x16bit_pipelined.layer_2_full_adder_2.cout ;
  wire \multiplier_16x16bit_pipelined.layer_2_full_adder_3.A ;
  wire \multiplier_16x16bit_pipelined.layer_2_full_adder_3.AB ;
  wire \multiplier_16x16bit_pipelined.layer_2_full_adder_3.AxorB ;
  wire \multiplier_16x16bit_pipelined.layer_2_full_adder_3.B ;
  wire \multiplier_16x16bit_pipelined.layer_2_full_adder_3.S ;
  wire \multiplier_16x16bit_pipelined.layer_2_full_adder_3.cin ;
  wire \multiplier_16x16bit_pipelined.layer_2_full_adder_3.cout ;
  wire \multiplier_16x16bit_pipelined.layer_2_full_adder_4.A ;
  wire \multiplier_16x16bit_pipelined.layer_2_full_adder_4.AB ;
  wire \multiplier_16x16bit_pipelined.layer_2_full_adder_4.AxorB ;
  wire \multiplier_16x16bit_pipelined.layer_2_full_adder_4.B ;
  wire \multiplier_16x16bit_pipelined.layer_2_full_adder_4.S ;
  wire \multiplier_16x16bit_pipelined.layer_2_full_adder_4.cin ;
  wire \multiplier_16x16bit_pipelined.layer_2_full_adder_4.cout ;
  wire \multiplier_16x16bit_pipelined.layer_2_full_adder_5.A ;
  wire \multiplier_16x16bit_pipelined.layer_2_full_adder_5.AB ;
  wire \multiplier_16x16bit_pipelined.layer_2_full_adder_5.AxorB ;
  wire \multiplier_16x16bit_pipelined.layer_2_full_adder_5.B ;
  wire \multiplier_16x16bit_pipelined.layer_2_full_adder_5.S ;
  wire \multiplier_16x16bit_pipelined.layer_2_full_adder_5.cin ;
  wire \multiplier_16x16bit_pipelined.layer_2_full_adder_5.cout ;
  wire \multiplier_16x16bit_pipelined.layer_2_full_adder_6.A ;
  wire \multiplier_16x16bit_pipelined.layer_2_full_adder_6.AB ;
  wire \multiplier_16x16bit_pipelined.layer_2_full_adder_6.AxorB ;
  wire \multiplier_16x16bit_pipelined.layer_2_full_adder_6.B ;
  wire \multiplier_16x16bit_pipelined.layer_2_full_adder_6.S ;
  wire \multiplier_16x16bit_pipelined.layer_2_full_adder_6.cin ;
  wire \multiplier_16x16bit_pipelined.layer_2_full_adder_6.cout ;
  wire \multiplier_16x16bit_pipelined.layer_2_full_adder_7.A ;
  wire \multiplier_16x16bit_pipelined.layer_2_full_adder_7.AB ;
  wire \multiplier_16x16bit_pipelined.layer_2_full_adder_7.AxorB ;
  wire \multiplier_16x16bit_pipelined.layer_2_full_adder_7.B ;
  wire \multiplier_16x16bit_pipelined.layer_2_full_adder_7.S ;
  wire \multiplier_16x16bit_pipelined.layer_2_full_adder_7.cin ;
  wire \multiplier_16x16bit_pipelined.layer_2_full_adder_7.cout ;
  wire \multiplier_16x16bit_pipelined.layer_2_full_adder_8.A ;
  wire \multiplier_16x16bit_pipelined.layer_2_full_adder_8.AB ;
  wire \multiplier_16x16bit_pipelined.layer_2_full_adder_8.AxorB ;
  wire \multiplier_16x16bit_pipelined.layer_2_full_adder_8.B ;
  wire \multiplier_16x16bit_pipelined.layer_2_full_adder_8.S ;
  wire \multiplier_16x16bit_pipelined.layer_2_full_adder_8.cin ;
  wire \multiplier_16x16bit_pipelined.layer_2_full_adder_8.cout ;
  wire \multiplier_16x16bit_pipelined.layer_2_full_adder_9.A ;
  wire \multiplier_16x16bit_pipelined.layer_2_full_adder_9.AB ;
  wire \multiplier_16x16bit_pipelined.layer_2_full_adder_9.AxorB ;
  wire \multiplier_16x16bit_pipelined.layer_2_full_adder_9.B ;
  wire \multiplier_16x16bit_pipelined.layer_2_full_adder_9.S ;
  wire \multiplier_16x16bit_pipelined.layer_2_full_adder_9.cin ;
  wire \multiplier_16x16bit_pipelined.layer_2_full_adder_9.cout ;
  wire [1:0] \multiplier_16x16bit_pipelined.layer_2_w0 ;
  wire \multiplier_16x16bit_pipelined.layer_2_w1 ;
  wire [1:0] \multiplier_16x16bit_pipelined.layer_2_w10 ;
  wire [3:0] \multiplier_16x16bit_pipelined.layer_2_w11 ;
  wire [2:0] \multiplier_16x16bit_pipelined.layer_2_w12 ;
  wire [2:0] \multiplier_16x16bit_pipelined.layer_2_w13 ;
  wire [2:0] \multiplier_16x16bit_pipelined.layer_2_w14 ;
  wire [2:0] \multiplier_16x16bit_pipelined.layer_2_w15 ;
  wire [2:0] \multiplier_16x16bit_pipelined.layer_2_w16 ;
  wire [2:0] \multiplier_16x16bit_pipelined.layer_2_w17 ;
  wire [3:0] \multiplier_16x16bit_pipelined.layer_2_w18 ;
  wire [2:0] \multiplier_16x16bit_pipelined.layer_2_w19 ;
  wire [2:0] \multiplier_16x16bit_pipelined.layer_2_w2 ;
  wire [3:0] \multiplier_16x16bit_pipelined.layer_2_w20 ;
  wire [1:0] \multiplier_16x16bit_pipelined.layer_2_w21 ;
  wire [1:0] \multiplier_16x16bit_pipelined.layer_2_w22 ;
  wire [1:0] \multiplier_16x16bit_pipelined.layer_2_w23 ;
  wire [2:0] \multiplier_16x16bit_pipelined.layer_2_w24 ;
  wire [1:0] \multiplier_16x16bit_pipelined.layer_2_w25 ;
  wire [2:0] \multiplier_16x16bit_pipelined.layer_2_w26 ;
  wire [1:0] \multiplier_16x16bit_pipelined.layer_2_w27 ;
  wire \multiplier_16x16bit_pipelined.layer_2_w28 ;
  wire [1:0] \multiplier_16x16bit_pipelined.layer_2_w29 ;
  wire [1:0] \multiplier_16x16bit_pipelined.layer_2_w3 ;
  wire \multiplier_16x16bit_pipelined.layer_2_w30 ;
  wire [1:0] \multiplier_16x16bit_pipelined.layer_2_w4 ;
  wire [1:0] \multiplier_16x16bit_pipelined.layer_2_w5 ;
  wire [1:0] \multiplier_16x16bit_pipelined.layer_2_w6 ;
  wire [1:0] \multiplier_16x16bit_pipelined.layer_2_w7 ;
  wire [1:0] \multiplier_16x16bit_pipelined.layer_2_w8 ;
  wire [1:0] \multiplier_16x16bit_pipelined.layer_2_w9 ;
  wire \multiplier_16x16bit_pipelined.layer_3_full_adder_0.A ;
  wire \multiplier_16x16bit_pipelined.layer_3_full_adder_0.AB ;
  wire \multiplier_16x16bit_pipelined.layer_3_full_adder_0.AxorB ;
  wire \multiplier_16x16bit_pipelined.layer_3_full_adder_0.B ;
  wire \multiplier_16x16bit_pipelined.layer_3_full_adder_0.S ;
  wire \multiplier_16x16bit_pipelined.layer_3_full_adder_0.cin ;
  wire \multiplier_16x16bit_pipelined.layer_3_full_adder_0.cout ;
  wire \multiplier_16x16bit_pipelined.layer_3_full_adder_1.A ;
  wire \multiplier_16x16bit_pipelined.layer_3_full_adder_1.AB ;
  wire \multiplier_16x16bit_pipelined.layer_3_full_adder_1.AxorB ;
  wire \multiplier_16x16bit_pipelined.layer_3_full_adder_1.B ;
  wire \multiplier_16x16bit_pipelined.layer_3_full_adder_1.S ;
  wire \multiplier_16x16bit_pipelined.layer_3_full_adder_1.cin ;
  wire \multiplier_16x16bit_pipelined.layer_3_full_adder_1.cout ;
  wire \multiplier_16x16bit_pipelined.layer_3_full_adder_10.A ;
  wire \multiplier_16x16bit_pipelined.layer_3_full_adder_10.AB ;
  wire \multiplier_16x16bit_pipelined.layer_3_full_adder_10.AxorB ;
  wire \multiplier_16x16bit_pipelined.layer_3_full_adder_10.B ;
  wire \multiplier_16x16bit_pipelined.layer_3_full_adder_10.S ;
  wire \multiplier_16x16bit_pipelined.layer_3_full_adder_10.cin ;
  wire \multiplier_16x16bit_pipelined.layer_3_full_adder_10.cout ;
  wire \multiplier_16x16bit_pipelined.layer_3_full_adder_11.A ;
  wire \multiplier_16x16bit_pipelined.layer_3_full_adder_11.AB ;
  wire \multiplier_16x16bit_pipelined.layer_3_full_adder_11.AxorB ;
  wire \multiplier_16x16bit_pipelined.layer_3_full_adder_11.B ;
  wire \multiplier_16x16bit_pipelined.layer_3_full_adder_11.S ;
  wire \multiplier_16x16bit_pipelined.layer_3_full_adder_11.cin ;
  wire \multiplier_16x16bit_pipelined.layer_3_full_adder_11.cout ;
  wire \multiplier_16x16bit_pipelined.layer_3_full_adder_12.A ;
  wire \multiplier_16x16bit_pipelined.layer_3_full_adder_12.AB ;
  wire \multiplier_16x16bit_pipelined.layer_3_full_adder_12.AxorB ;
  wire \multiplier_16x16bit_pipelined.layer_3_full_adder_12.B ;
  wire \multiplier_16x16bit_pipelined.layer_3_full_adder_12.S ;
  wire \multiplier_16x16bit_pipelined.layer_3_full_adder_12.cin ;
  wire \multiplier_16x16bit_pipelined.layer_3_full_adder_12.cout ;
  wire \multiplier_16x16bit_pipelined.layer_3_full_adder_13.A ;
  wire \multiplier_16x16bit_pipelined.layer_3_full_adder_13.AB ;
  wire \multiplier_16x16bit_pipelined.layer_3_full_adder_13.AxorB ;
  wire \multiplier_16x16bit_pipelined.layer_3_full_adder_13.B ;
  wire \multiplier_16x16bit_pipelined.layer_3_full_adder_13.S ;
  wire \multiplier_16x16bit_pipelined.layer_3_full_adder_13.cin ;
  wire \multiplier_16x16bit_pipelined.layer_3_full_adder_13.cout ;
  wire \multiplier_16x16bit_pipelined.layer_3_full_adder_2.A ;
  wire \multiplier_16x16bit_pipelined.layer_3_full_adder_2.AB ;
  wire \multiplier_16x16bit_pipelined.layer_3_full_adder_2.AxorB ;
  wire \multiplier_16x16bit_pipelined.layer_3_full_adder_2.B ;
  wire \multiplier_16x16bit_pipelined.layer_3_full_adder_2.S ;
  wire \multiplier_16x16bit_pipelined.layer_3_full_adder_2.cin ;
  wire \multiplier_16x16bit_pipelined.layer_3_full_adder_2.cout ;
  wire \multiplier_16x16bit_pipelined.layer_3_full_adder_3.A ;
  wire \multiplier_16x16bit_pipelined.layer_3_full_adder_3.AB ;
  wire \multiplier_16x16bit_pipelined.layer_3_full_adder_3.AxorB ;
  wire \multiplier_16x16bit_pipelined.layer_3_full_adder_3.B ;
  wire \multiplier_16x16bit_pipelined.layer_3_full_adder_3.S ;
  wire \multiplier_16x16bit_pipelined.layer_3_full_adder_3.cin ;
  wire \multiplier_16x16bit_pipelined.layer_3_full_adder_3.cout ;
  wire \multiplier_16x16bit_pipelined.layer_3_full_adder_4.A ;
  wire \multiplier_16x16bit_pipelined.layer_3_full_adder_4.AB ;
  wire \multiplier_16x16bit_pipelined.layer_3_full_adder_4.AxorB ;
  wire \multiplier_16x16bit_pipelined.layer_3_full_adder_4.B ;
  wire \multiplier_16x16bit_pipelined.layer_3_full_adder_4.S ;
  wire \multiplier_16x16bit_pipelined.layer_3_full_adder_4.cin ;
  wire \multiplier_16x16bit_pipelined.layer_3_full_adder_4.cout ;
  wire \multiplier_16x16bit_pipelined.layer_3_full_adder_5.A ;
  wire \multiplier_16x16bit_pipelined.layer_3_full_adder_5.AB ;
  wire \multiplier_16x16bit_pipelined.layer_3_full_adder_5.AxorB ;
  wire \multiplier_16x16bit_pipelined.layer_3_full_adder_5.B ;
  wire \multiplier_16x16bit_pipelined.layer_3_full_adder_5.S ;
  wire \multiplier_16x16bit_pipelined.layer_3_full_adder_5.cin ;
  wire \multiplier_16x16bit_pipelined.layer_3_full_adder_5.cout ;
  wire \multiplier_16x16bit_pipelined.layer_3_full_adder_6.A ;
  wire \multiplier_16x16bit_pipelined.layer_3_full_adder_6.AB ;
  wire \multiplier_16x16bit_pipelined.layer_3_full_adder_6.AxorB ;
  wire \multiplier_16x16bit_pipelined.layer_3_full_adder_6.B ;
  wire \multiplier_16x16bit_pipelined.layer_3_full_adder_6.S ;
  wire \multiplier_16x16bit_pipelined.layer_3_full_adder_6.cin ;
  wire \multiplier_16x16bit_pipelined.layer_3_full_adder_6.cout ;
  wire \multiplier_16x16bit_pipelined.layer_3_full_adder_7.A ;
  wire \multiplier_16x16bit_pipelined.layer_3_full_adder_7.AB ;
  wire \multiplier_16x16bit_pipelined.layer_3_full_adder_7.AxorB ;
  wire \multiplier_16x16bit_pipelined.layer_3_full_adder_7.B ;
  wire \multiplier_16x16bit_pipelined.layer_3_full_adder_7.S ;
  wire \multiplier_16x16bit_pipelined.layer_3_full_adder_7.cin ;
  wire \multiplier_16x16bit_pipelined.layer_3_full_adder_7.cout ;
  wire \multiplier_16x16bit_pipelined.layer_3_full_adder_8.A ;
  wire \multiplier_16x16bit_pipelined.layer_3_full_adder_8.AB ;
  wire \multiplier_16x16bit_pipelined.layer_3_full_adder_8.AxorB ;
  wire \multiplier_16x16bit_pipelined.layer_3_full_adder_8.B ;
  wire \multiplier_16x16bit_pipelined.layer_3_full_adder_8.S ;
  wire \multiplier_16x16bit_pipelined.layer_3_full_adder_8.cin ;
  wire \multiplier_16x16bit_pipelined.layer_3_full_adder_8.cout ;
  wire \multiplier_16x16bit_pipelined.layer_3_full_adder_9.A ;
  wire \multiplier_16x16bit_pipelined.layer_3_full_adder_9.AB ;
  wire \multiplier_16x16bit_pipelined.layer_3_full_adder_9.AxorB ;
  wire \multiplier_16x16bit_pipelined.layer_3_full_adder_9.B ;
  wire \multiplier_16x16bit_pipelined.layer_3_full_adder_9.S ;
  wire \multiplier_16x16bit_pipelined.layer_3_full_adder_9.cin ;
  wire \multiplier_16x16bit_pipelined.layer_3_full_adder_9.cout ;
  wire \multiplier_16x16bit_pipelined.layer_3_w0[0] ;
  wire \multiplier_16x16bit_pipelined.layer_3_w0[1] ;
  wire \multiplier_16x16bit_pipelined.layer_3_w1 ;
  wire \multiplier_16x16bit_pipelined.layer_3_w10[0] ;
  wire \multiplier_16x16bit_pipelined.layer_3_w10[1] ;
  wire \multiplier_16x16bit_pipelined.layer_3_w11[0] ;
  wire \multiplier_16x16bit_pipelined.layer_3_w11[1] ;
  wire \multiplier_16x16bit_pipelined.layer_3_w12[0] ;
  wire \multiplier_16x16bit_pipelined.layer_3_w12[1] ;
  wire \multiplier_16x16bit_pipelined.layer_3_w13[0] ;
  wire \multiplier_16x16bit_pipelined.layer_3_w13[1] ;
  wire \multiplier_16x16bit_pipelined.layer_3_w14[0] ;
  wire \multiplier_16x16bit_pipelined.layer_3_w14[1] ;
  wire \multiplier_16x16bit_pipelined.layer_3_w15[0] ;
  wire \multiplier_16x16bit_pipelined.layer_3_w15[1] ;
  wire \multiplier_16x16bit_pipelined.layer_3_w16[0] ;
  wire \multiplier_16x16bit_pipelined.layer_3_w16[1] ;
  wire \multiplier_16x16bit_pipelined.layer_3_w16[2] ;
  wire \multiplier_16x16bit_pipelined.layer_3_w17[0] ;
  wire \multiplier_16x16bit_pipelined.layer_3_w17[1] ;
  wire \multiplier_16x16bit_pipelined.layer_3_w18[0] ;
  wire \multiplier_16x16bit_pipelined.layer_3_w18[1] ;
  wire \multiplier_16x16bit_pipelined.layer_3_w18[2] ;
  wire \multiplier_16x16bit_pipelined.layer_3_w19[0] ;
  wire \multiplier_16x16bit_pipelined.layer_3_w19[1] ;
  wire \multiplier_16x16bit_pipelined.layer_3_w20[0] ;
  wire \multiplier_16x16bit_pipelined.layer_3_w20[1] ;
  wire \multiplier_16x16bit_pipelined.layer_3_w20[2] ;
  wire \multiplier_16x16bit_pipelined.layer_3_w21[0] ;
  wire \multiplier_16x16bit_pipelined.layer_3_w21[1] ;
  wire \multiplier_16x16bit_pipelined.layer_3_w22[0] ;
  wire \multiplier_16x16bit_pipelined.layer_3_w22[1] ;
  wire \multiplier_16x16bit_pipelined.layer_3_w22[2] ;
  wire \multiplier_16x16bit_pipelined.layer_3_w23[0] ;
  wire \multiplier_16x16bit_pipelined.layer_3_w23[1] ;
  wire \multiplier_16x16bit_pipelined.layer_3_w24 ;
  wire \multiplier_16x16bit_pipelined.layer_3_w25[0] ;
  wire \multiplier_16x16bit_pipelined.layer_3_w25[1] ;
  wire \multiplier_16x16bit_pipelined.layer_3_w25[2] ;
  wire \multiplier_16x16bit_pipelined.layer_3_w26 ;
  wire \multiplier_16x16bit_pipelined.layer_3_w27[0] ;
  wire \multiplier_16x16bit_pipelined.layer_3_w27[1] ;
  wire \multiplier_16x16bit_pipelined.layer_3_w27[2] ;
  wire \multiplier_16x16bit_pipelined.layer_3_w28 ;
  wire \multiplier_16x16bit_pipelined.layer_3_w29 ;
  wire \multiplier_16x16bit_pipelined.layer_3_w2[0] ;
  wire \multiplier_16x16bit_pipelined.layer_3_w2[1] ;
  wire \multiplier_16x16bit_pipelined.layer_3_w2[2] ;
  wire \multiplier_16x16bit_pipelined.layer_3_w30[0] ;
  wire \multiplier_16x16bit_pipelined.layer_3_w30[1] ;
  wire \multiplier_16x16bit_pipelined.layer_3_w31 ;
  wire \multiplier_16x16bit_pipelined.layer_3_w3[0] ;
  wire \multiplier_16x16bit_pipelined.layer_3_w3[1] ;
  wire \multiplier_16x16bit_pipelined.layer_3_w4[0] ;
  wire \multiplier_16x16bit_pipelined.layer_3_w4[1] ;
  wire \multiplier_16x16bit_pipelined.layer_3_w5[0] ;
  wire \multiplier_16x16bit_pipelined.layer_3_w5[1] ;
  wire \multiplier_16x16bit_pipelined.layer_3_w6[0] ;
  wire \multiplier_16x16bit_pipelined.layer_3_w6[1] ;
  wire \multiplier_16x16bit_pipelined.layer_3_w7[0] ;
  wire \multiplier_16x16bit_pipelined.layer_3_w7[1] ;
  wire \multiplier_16x16bit_pipelined.layer_3_w8[0] ;
  wire \multiplier_16x16bit_pipelined.layer_3_w8[1] ;
  wire \multiplier_16x16bit_pipelined.layer_3_w9[0] ;
  wire \multiplier_16x16bit_pipelined.layer_3_w9[1] ;
  wire \multiplier_16x16bit_pipelined.layer_4_full_adder_0.A ;
  wire \multiplier_16x16bit_pipelined.layer_4_full_adder_0.AB ;
  wire \multiplier_16x16bit_pipelined.layer_4_full_adder_0.AxorB ;
  wire \multiplier_16x16bit_pipelined.layer_4_full_adder_0.B ;
  wire \multiplier_16x16bit_pipelined.layer_4_full_adder_0.S ;
  wire \multiplier_16x16bit_pipelined.layer_4_full_adder_0.cin ;
  wire \multiplier_16x16bit_pipelined.layer_4_full_adder_0.cout ;
  wire \multiplier_16x16bit_pipelined.layer_4_full_adder_1.A ;
  wire \multiplier_16x16bit_pipelined.layer_4_full_adder_1.AB ;
  wire \multiplier_16x16bit_pipelined.layer_4_full_adder_1.AxorB ;
  wire \multiplier_16x16bit_pipelined.layer_4_full_adder_1.B ;
  wire \multiplier_16x16bit_pipelined.layer_4_full_adder_1.S ;
  wire \multiplier_16x16bit_pipelined.layer_4_full_adder_1.cin ;
  wire \multiplier_16x16bit_pipelined.layer_4_full_adder_1.cout ;
  wire \multiplier_16x16bit_pipelined.layer_4_full_adder_2.A ;
  wire \multiplier_16x16bit_pipelined.layer_4_full_adder_2.AB ;
  wire \multiplier_16x16bit_pipelined.layer_4_full_adder_2.AxorB ;
  wire \multiplier_16x16bit_pipelined.layer_4_full_adder_2.B ;
  wire \multiplier_16x16bit_pipelined.layer_4_full_adder_2.S ;
  wire \multiplier_16x16bit_pipelined.layer_4_full_adder_2.cin ;
  wire \multiplier_16x16bit_pipelined.layer_4_full_adder_2.cout ;
  wire \multiplier_16x16bit_pipelined.layer_4_full_adder_3.A ;
  wire \multiplier_16x16bit_pipelined.layer_4_full_adder_3.AB ;
  wire \multiplier_16x16bit_pipelined.layer_4_full_adder_3.AxorB ;
  wire \multiplier_16x16bit_pipelined.layer_4_full_adder_3.B ;
  wire \multiplier_16x16bit_pipelined.layer_4_full_adder_3.S ;
  wire \multiplier_16x16bit_pipelined.layer_4_full_adder_3.cin ;
  wire \multiplier_16x16bit_pipelined.layer_4_full_adder_3.cout ;
  wire \multiplier_16x16bit_pipelined.layer_4_full_adder_4.A ;
  wire \multiplier_16x16bit_pipelined.layer_4_full_adder_4.AB ;
  wire \multiplier_16x16bit_pipelined.layer_4_full_adder_4.AxorB ;
  wire \multiplier_16x16bit_pipelined.layer_4_full_adder_4.B ;
  wire \multiplier_16x16bit_pipelined.layer_4_full_adder_4.S ;
  wire \multiplier_16x16bit_pipelined.layer_4_full_adder_4.cin ;
  wire \multiplier_16x16bit_pipelined.layer_4_full_adder_4.cout ;
  wire \multiplier_16x16bit_pipelined.layer_4_full_adder_5.A ;
  wire \multiplier_16x16bit_pipelined.layer_4_full_adder_5.AB ;
  wire \multiplier_16x16bit_pipelined.layer_4_full_adder_5.AxorB ;
  wire \multiplier_16x16bit_pipelined.layer_4_full_adder_5.B ;
  wire \multiplier_16x16bit_pipelined.layer_4_full_adder_5.S ;
  wire \multiplier_16x16bit_pipelined.layer_4_full_adder_5.cin ;
  wire \multiplier_16x16bit_pipelined.layer_4_full_adder_5.cout ;
  wire \multiplier_16x16bit_pipelined.layer_4_full_adder_6.A ;
  wire \multiplier_16x16bit_pipelined.layer_4_full_adder_6.AB ;
  wire \multiplier_16x16bit_pipelined.layer_4_full_adder_6.AxorB ;
  wire \multiplier_16x16bit_pipelined.layer_4_full_adder_6.B ;
  wire \multiplier_16x16bit_pipelined.layer_4_full_adder_6.S ;
  wire \multiplier_16x16bit_pipelined.layer_4_full_adder_6.cin ;
  wire \multiplier_16x16bit_pipelined.layer_4_full_adder_6.cout ;
  wire \multiplier_16x16bit_pipelined.layer_4_half_adder_0.A ;
  wire \multiplier_16x16bit_pipelined.layer_4_half_adder_0.B ;
  wire \multiplier_16x16bit_pipelined.layer_4_half_adder_0.S ;
  wire \multiplier_16x16bit_pipelined.layer_4_half_adder_0.carry ;
  wire \multiplier_16x16bit_pipelined.layer_4_half_adder_1.A ;
  wire \multiplier_16x16bit_pipelined.layer_4_half_adder_1.B ;
  wire \multiplier_16x16bit_pipelined.layer_4_half_adder_1.S ;
  wire \multiplier_16x16bit_pipelined.layer_4_half_adder_1.carry ;
  wire \multiplier_16x16bit_pipelined.layer_4_half_adder_10.A ;
  wire \multiplier_16x16bit_pipelined.layer_4_half_adder_10.B ;
  wire \multiplier_16x16bit_pipelined.layer_4_half_adder_10.S ;
  wire \multiplier_16x16bit_pipelined.layer_4_half_adder_10.carry ;
  wire \multiplier_16x16bit_pipelined.layer_4_half_adder_11.A ;
  wire \multiplier_16x16bit_pipelined.layer_4_half_adder_11.B ;
  wire \multiplier_16x16bit_pipelined.layer_4_half_adder_11.S ;
  wire \multiplier_16x16bit_pipelined.layer_4_half_adder_11.carry ;
  wire \multiplier_16x16bit_pipelined.layer_4_half_adder_12.A ;
  wire \multiplier_16x16bit_pipelined.layer_4_half_adder_12.B ;
  wire \multiplier_16x16bit_pipelined.layer_4_half_adder_12.S ;
  wire \multiplier_16x16bit_pipelined.layer_4_half_adder_12.carry ;
  wire \multiplier_16x16bit_pipelined.layer_4_half_adder_13.A ;
  wire \multiplier_16x16bit_pipelined.layer_4_half_adder_13.B ;
  wire \multiplier_16x16bit_pipelined.layer_4_half_adder_13.S ;
  wire \multiplier_16x16bit_pipelined.layer_4_half_adder_13.carry ;
  wire \multiplier_16x16bit_pipelined.layer_4_half_adder_14.A ;
  wire \multiplier_16x16bit_pipelined.layer_4_half_adder_14.B ;
  wire \multiplier_16x16bit_pipelined.layer_4_half_adder_14.S ;
  wire \multiplier_16x16bit_pipelined.layer_4_half_adder_14.carry ;
  wire \multiplier_16x16bit_pipelined.layer_4_half_adder_15.A ;
  wire \multiplier_16x16bit_pipelined.layer_4_half_adder_15.B ;
  wire \multiplier_16x16bit_pipelined.layer_4_half_adder_15.S ;
  wire \multiplier_16x16bit_pipelined.layer_4_half_adder_15.carry ;
  wire \multiplier_16x16bit_pipelined.layer_4_half_adder_16.A ;
  wire \multiplier_16x16bit_pipelined.layer_4_half_adder_16.B ;
  wire \multiplier_16x16bit_pipelined.layer_4_half_adder_16.S ;
  wire \multiplier_16x16bit_pipelined.layer_4_half_adder_16.carry ;
  wire \multiplier_16x16bit_pipelined.layer_4_half_adder_2.A ;
  wire \multiplier_16x16bit_pipelined.layer_4_half_adder_2.B ;
  wire \multiplier_16x16bit_pipelined.layer_4_half_adder_2.S ;
  wire \multiplier_16x16bit_pipelined.layer_4_half_adder_2.carry ;
  wire \multiplier_16x16bit_pipelined.layer_4_half_adder_3.A ;
  wire \multiplier_16x16bit_pipelined.layer_4_half_adder_3.B ;
  wire \multiplier_16x16bit_pipelined.layer_4_half_adder_3.S ;
  wire \multiplier_16x16bit_pipelined.layer_4_half_adder_3.carry ;
  wire \multiplier_16x16bit_pipelined.layer_4_half_adder_4.A ;
  wire \multiplier_16x16bit_pipelined.layer_4_half_adder_4.B ;
  wire \multiplier_16x16bit_pipelined.layer_4_half_adder_4.S ;
  wire \multiplier_16x16bit_pipelined.layer_4_half_adder_4.carry ;
  wire \multiplier_16x16bit_pipelined.layer_4_half_adder_5.A ;
  wire \multiplier_16x16bit_pipelined.layer_4_half_adder_5.B ;
  wire \multiplier_16x16bit_pipelined.layer_4_half_adder_5.S ;
  wire \multiplier_16x16bit_pipelined.layer_4_half_adder_5.carry ;
  wire \multiplier_16x16bit_pipelined.layer_4_half_adder_6.A ;
  wire \multiplier_16x16bit_pipelined.layer_4_half_adder_6.B ;
  wire \multiplier_16x16bit_pipelined.layer_4_half_adder_6.S ;
  wire \multiplier_16x16bit_pipelined.layer_4_half_adder_6.carry ;
  wire \multiplier_16x16bit_pipelined.layer_4_half_adder_7.A ;
  wire \multiplier_16x16bit_pipelined.layer_4_half_adder_7.B ;
  wire \multiplier_16x16bit_pipelined.layer_4_half_adder_7.S ;
  wire \multiplier_16x16bit_pipelined.layer_4_half_adder_7.carry ;
  wire \multiplier_16x16bit_pipelined.layer_4_half_adder_8.A ;
  wire \multiplier_16x16bit_pipelined.layer_4_half_adder_8.B ;
  wire \multiplier_16x16bit_pipelined.layer_4_half_adder_8.S ;
  wire \multiplier_16x16bit_pipelined.layer_4_half_adder_8.carry ;
  wire \multiplier_16x16bit_pipelined.layer_4_half_adder_9.A ;
  wire \multiplier_16x16bit_pipelined.layer_4_half_adder_9.B ;
  wire \multiplier_16x16bit_pipelined.layer_4_half_adder_9.S ;
  wire \multiplier_16x16bit_pipelined.layer_4_half_adder_9.carry ;
  wire \multiplier_16x16bit_pipelined.layer_4_w0[0] ;
  wire \multiplier_16x16bit_pipelined.layer_4_w0[1] ;
  wire \multiplier_16x16bit_pipelined.layer_4_w1 ;
  wire \multiplier_16x16bit_pipelined.layer_4_w10[0] ;
  wire \multiplier_16x16bit_pipelined.layer_4_w10[1] ;
  wire \multiplier_16x16bit_pipelined.layer_4_w11[0] ;
  wire \multiplier_16x16bit_pipelined.layer_4_w11[1] ;
  wire \multiplier_16x16bit_pipelined.layer_4_w12[0] ;
  wire \multiplier_16x16bit_pipelined.layer_4_w12[1] ;
  wire \multiplier_16x16bit_pipelined.layer_4_w13[0] ;
  wire \multiplier_16x16bit_pipelined.layer_4_w13[1] ;
  wire \multiplier_16x16bit_pipelined.layer_4_w14[0] ;
  wire \multiplier_16x16bit_pipelined.layer_4_w14[1] ;
  wire \multiplier_16x16bit_pipelined.layer_4_w15[0] ;
  wire \multiplier_16x16bit_pipelined.layer_4_w15[1] ;
  wire \multiplier_16x16bit_pipelined.layer_4_w16[0] ;
  wire \multiplier_16x16bit_pipelined.layer_4_w16[1] ;
  wire \multiplier_16x16bit_pipelined.layer_4_w17[0] ;
  wire \multiplier_16x16bit_pipelined.layer_4_w17[1] ;
  wire \multiplier_16x16bit_pipelined.layer_4_w18[0] ;
  wire \multiplier_16x16bit_pipelined.layer_4_w18[1] ;
  wire \multiplier_16x16bit_pipelined.layer_4_w19[0] ;
  wire \multiplier_16x16bit_pipelined.layer_4_w19[1] ;
  wire \multiplier_16x16bit_pipelined.layer_4_w2 ;
  wire \multiplier_16x16bit_pipelined.layer_4_w20[0] ;
  wire \multiplier_16x16bit_pipelined.layer_4_w20[1] ;
  wire \multiplier_16x16bit_pipelined.layer_4_w21[0] ;
  wire \multiplier_16x16bit_pipelined.layer_4_w21[1] ;
  wire \multiplier_16x16bit_pipelined.layer_4_w22[0] ;
  wire \multiplier_16x16bit_pipelined.layer_4_w22[1] ;
  wire \multiplier_16x16bit_pipelined.layer_4_w23[0] ;
  wire \multiplier_16x16bit_pipelined.layer_4_w23[1] ;
  wire \multiplier_16x16bit_pipelined.layer_4_w24[0] ;
  wire \multiplier_16x16bit_pipelined.layer_4_w24[1] ;
  wire \multiplier_16x16bit_pipelined.layer_4_w25 ;
  wire \multiplier_16x16bit_pipelined.layer_4_w26[0] ;
  wire \multiplier_16x16bit_pipelined.layer_4_w26[1] ;
  wire \multiplier_16x16bit_pipelined.layer_4_w27 ;
  wire \multiplier_16x16bit_pipelined.layer_4_w28[0] ;
  wire \multiplier_16x16bit_pipelined.layer_4_w28[1] ;
  wire \multiplier_16x16bit_pipelined.layer_4_w29 ;
  wire \multiplier_16x16bit_pipelined.layer_4_w30[0] ;
  wire \multiplier_16x16bit_pipelined.layer_4_w30[1] ;
  wire \multiplier_16x16bit_pipelined.layer_4_w31 ;
  wire \multiplier_16x16bit_pipelined.layer_4_w3[0] ;
  wire \multiplier_16x16bit_pipelined.layer_4_w3[1] ;
  wire \multiplier_16x16bit_pipelined.layer_4_w4[0] ;
  wire \multiplier_16x16bit_pipelined.layer_4_w4[1] ;
  wire \multiplier_16x16bit_pipelined.layer_4_w5[0] ;
  wire \multiplier_16x16bit_pipelined.layer_4_w5[1] ;
  wire \multiplier_16x16bit_pipelined.layer_4_w6[0] ;
  wire \multiplier_16x16bit_pipelined.layer_4_w6[1] ;
  wire \multiplier_16x16bit_pipelined.layer_4_w7[0] ;
  wire \multiplier_16x16bit_pipelined.layer_4_w7[1] ;
  wire \multiplier_16x16bit_pipelined.layer_4_w8[0] ;
  wire \multiplier_16x16bit_pipelined.layer_4_w8[1] ;
  wire \multiplier_16x16bit_pipelined.layer_4_w9[0] ;
  wire \multiplier_16x16bit_pipelined.layer_4_w9[1] ;
  reg [15:0] \multiplier_16x16bit_pipelined.md ;
  reg [15:0] \multiplier_16x16bit_pipelined.mr ;
  wire [7:0] \multiplier_16x16bit_pipelined.negation ;
  wire [31:0] \multiplier_16x16bit_pipelined.o_product ;
  wire \multiplier_16x16bit_pipelined.partial_product_gen_0.double ;
  wire [15:0] \multiplier_16x16bit_pipelined.partial_product_gen_0.md ;
  wire \multiplier_16x16bit_pipelined.partial_product_gen_0.negation ;
  wire [15:0] \multiplier_16x16bit_pipelined.partial_product_gen_0.nmd ;
  wire [16:0] \multiplier_16x16bit_pipelined.partial_product_gen_0.pp ;
  wire \multiplier_16x16bit_pipelined.partial_product_gen_0.zero ;
  wire [15:0] \multiplier_16x16bit_pipelined.partial_product_gen_0.zmd ;
  wire \multiplier_16x16bit_pipelined.partial_product_gen_1.double ;
  wire [15:0] \multiplier_16x16bit_pipelined.partial_product_gen_1.md ;
  wire \multiplier_16x16bit_pipelined.partial_product_gen_1.negation ;
  wire [15:0] \multiplier_16x16bit_pipelined.partial_product_gen_1.nmd ;
  wire [16:0] \multiplier_16x16bit_pipelined.partial_product_gen_1.pp ;
  wire \multiplier_16x16bit_pipelined.partial_product_gen_1.zero ;
  wire [15:0] \multiplier_16x16bit_pipelined.partial_product_gen_1.zmd ;
  wire \multiplier_16x16bit_pipelined.partial_product_gen_2.double ;
  wire [15:0] \multiplier_16x16bit_pipelined.partial_product_gen_2.md ;
  wire \multiplier_16x16bit_pipelined.partial_product_gen_2.negation ;
  wire [15:0] \multiplier_16x16bit_pipelined.partial_product_gen_2.nmd ;
  wire [16:0] \multiplier_16x16bit_pipelined.partial_product_gen_2.pp ;
  wire \multiplier_16x16bit_pipelined.partial_product_gen_2.zero ;
  wire [15:0] \multiplier_16x16bit_pipelined.partial_product_gen_2.zmd ;
  wire \multiplier_16x16bit_pipelined.partial_product_gen_3.double ;
  wire [15:0] \multiplier_16x16bit_pipelined.partial_product_gen_3.md ;
  wire \multiplier_16x16bit_pipelined.partial_product_gen_3.negation ;
  wire [15:0] \multiplier_16x16bit_pipelined.partial_product_gen_3.nmd ;
  wire [16:0] \multiplier_16x16bit_pipelined.partial_product_gen_3.pp ;
  wire \multiplier_16x16bit_pipelined.partial_product_gen_3.zero ;
  wire [15:0] \multiplier_16x16bit_pipelined.partial_product_gen_3.zmd ;
  wire \multiplier_16x16bit_pipelined.partial_product_gen_4.double ;
  wire [15:0] \multiplier_16x16bit_pipelined.partial_product_gen_4.md ;
  wire \multiplier_16x16bit_pipelined.partial_product_gen_4.negation ;
  wire [15:0] \multiplier_16x16bit_pipelined.partial_product_gen_4.nmd ;
  wire [16:0] \multiplier_16x16bit_pipelined.partial_product_gen_4.pp ;
  wire \multiplier_16x16bit_pipelined.partial_product_gen_4.zero ;
  wire [15:0] \multiplier_16x16bit_pipelined.partial_product_gen_4.zmd ;
  wire \multiplier_16x16bit_pipelined.partial_product_gen_5.double ;
  wire [15:0] \multiplier_16x16bit_pipelined.partial_product_gen_5.md ;
  wire \multiplier_16x16bit_pipelined.partial_product_gen_5.negation ;
  wire [15:0] \multiplier_16x16bit_pipelined.partial_product_gen_5.nmd ;
  wire [16:0] \multiplier_16x16bit_pipelined.partial_product_gen_5.pp ;
  wire \multiplier_16x16bit_pipelined.partial_product_gen_5.zero ;
  wire [15:0] \multiplier_16x16bit_pipelined.partial_product_gen_5.zmd ;
  wire \multiplier_16x16bit_pipelined.partial_product_gen_6.double ;
  wire [15:0] \multiplier_16x16bit_pipelined.partial_product_gen_6.md ;
  wire \multiplier_16x16bit_pipelined.partial_product_gen_6.negation ;
  wire [15:0] \multiplier_16x16bit_pipelined.partial_product_gen_6.nmd ;
  wire [16:0] \multiplier_16x16bit_pipelined.partial_product_gen_6.pp ;
  wire \multiplier_16x16bit_pipelined.partial_product_gen_6.zero ;
  wire [15:0] \multiplier_16x16bit_pipelined.partial_product_gen_6.zmd ;
  wire \multiplier_16x16bit_pipelined.partial_product_gen_7.double ;
  wire [15:0] \multiplier_16x16bit_pipelined.partial_product_gen_7.md ;
  wire \multiplier_16x16bit_pipelined.partial_product_gen_7.negation ;
  wire [15:0] \multiplier_16x16bit_pipelined.partial_product_gen_7.nmd ;
  wire [16:0] \multiplier_16x16bit_pipelined.partial_product_gen_7.pp ;
  wire \multiplier_16x16bit_pipelined.partial_product_gen_7.zero ;
  wire [15:0] \multiplier_16x16bit_pipelined.partial_product_gen_7.zmd ;
  reg [1:0] \multiplier_16x16bit_pipelined.reg_layer_2_w0 ;
  reg \multiplier_16x16bit_pipelined.reg_layer_2_w1 ;
  reg [1:0] \multiplier_16x16bit_pipelined.reg_layer_2_w10 ;
  reg [3:0] \multiplier_16x16bit_pipelined.reg_layer_2_w11 ;
  reg [2:0] \multiplier_16x16bit_pipelined.reg_layer_2_w12 ;
  reg [2:0] \multiplier_16x16bit_pipelined.reg_layer_2_w13 ;
  reg [2:0] \multiplier_16x16bit_pipelined.reg_layer_2_w14 ;
  reg [2:0] \multiplier_16x16bit_pipelined.reg_layer_2_w15 ;
  reg [3:0] \multiplier_16x16bit_pipelined.reg_layer_2_w16 ;
  reg [2:0] \multiplier_16x16bit_pipelined.reg_layer_2_w17 ;
  reg [3:0] \multiplier_16x16bit_pipelined.reg_layer_2_w18 ;
  reg [2:0] \multiplier_16x16bit_pipelined.reg_layer_2_w19 ;
  reg [2:0] \multiplier_16x16bit_pipelined.reg_layer_2_w2 ;
  reg [3:0] \multiplier_16x16bit_pipelined.reg_layer_2_w20 ;
  reg [2:0] \multiplier_16x16bit_pipelined.reg_layer_2_w21 ;
  reg [1:0] \multiplier_16x16bit_pipelined.reg_layer_2_w22 ;
  reg [1:0] \multiplier_16x16bit_pipelined.reg_layer_2_w23 ;
  reg [2:0] \multiplier_16x16bit_pipelined.reg_layer_2_w24 ;
  reg [1:0] \multiplier_16x16bit_pipelined.reg_layer_2_w25 ;
  reg [2:0] \multiplier_16x16bit_pipelined.reg_layer_2_w26 ;
  reg [1:0] \multiplier_16x16bit_pipelined.reg_layer_2_w27 ;
  reg \multiplier_16x16bit_pipelined.reg_layer_2_w28 ;
  reg [2:0] \multiplier_16x16bit_pipelined.reg_layer_2_w29 ;
  reg [1:0] \multiplier_16x16bit_pipelined.reg_layer_2_w3 ;
  reg \multiplier_16x16bit_pipelined.reg_layer_2_w30 ;
  reg \multiplier_16x16bit_pipelined.reg_layer_2_w31 ;
  reg [1:0] \multiplier_16x16bit_pipelined.reg_layer_2_w4 ;
  reg [1:0] \multiplier_16x16bit_pipelined.reg_layer_2_w5 ;
  reg [1:0] \multiplier_16x16bit_pipelined.reg_layer_2_w6 ;
  reg [1:0] \multiplier_16x16bit_pipelined.reg_layer_2_w7 ;
  reg [1:0] \multiplier_16x16bit_pipelined.reg_layer_2_w8 ;
  reg [1:0] \multiplier_16x16bit_pipelined.reg_layer_2_w9 ;
  reg \multiplier_16x16bit_pipelined.stage_0_ready ;
  wire [7:0] \multiplier_16x16bit_pipelined.zero ;
  output [31:0] o_un;
  output o_valid;
  output o_wb_ack;
  output [31:0] o_wb_data;
  reg [4:0] of;
  wire \of_addition[0] ;
  wire \of_addition[1] ;
  reg [31:0] p;
  wire [31:0] product;
  reg [15:0] pv;
  wire rack;
  wire [31:0] \rdata[0] ;
  wire [31:0] \rdata[10] ;
  wire [31:0] \rdata[1] ;
  wire [31:0] \rdata[2] ;
  wire [31:0] \rdata[3] ;
  wire [31:0] \rdata[4] ;
  wire [31:0] \rdata[5] ;
  wire [31:0] \rdata[6] ;
  wire [31:0] \rdata[7] ;
  wire [31:0] \rdata[8] ;
  wire [31:0] \rdata[9] ;
  wire re;
  wire [10:0] rl;
  reg rla;
  reg rlb;
  reg [31:0] sigma;
  reg [15:0] sp;
  reg start;
  reg state_0;
  reg [9:0] state_1;
  wire [31:0] sum;
  reg [31:0] un;
  wire update_esu;
  wire update_kpd;
  reg wack;
  wire we;
  wire [0:7] wl;
  wire wlRS;
  reg wla;
  reg wlb;
  assign _0026_ = i_wb_cyc & i_wb_we;
  assign we = _0026_ & i_wb_stb;
  assign _0027_ = i_wb_cyc & _0070_;
  assign re = _0027_ & i_wb_stb;
  assign _0028_ = re & adr_check_1;
  assign _0029_ = _0028_ & _0077_;
  assign _0030_ = re & _0078_;
  assign o_wb_ack = _0081_ & i_wb_stb;
  assign _0036_ = 3'b111 - i_wb_adr[4:2];
  assign _0037_ = 4'b1111 - i_wb_adr[5:2];
  wire [4:0] fangyuan0;
  assign fangyuan0 = { _0082_, _0083_, _0084_, _0039_, _0085_ };

  assign _0031_ = | fangyuan0;
  wire [1:0] fangyuan1;
  assign fangyuan1 = { _0101_, _0102_ };

  assign _0032_ = | fangyuan1;
  wire [1:0] fangyuan2;
  assign fangyuan2 = { _0096_, _0102_ };

  assign _0033_ = | fangyuan2;
  wire [2:0] fangyuan3;
  assign fangyuan3 = { _0096_, _0102_, _0121_ };

  assign _0034_ = | fangyuan3;
  wire [1:0] fangyuan4;
  assign fangyuan4 = { _0101_, _0113_ };

  assign _0035_ = | fangyuan4;
  assign adr_check_1 = ! i_wb_adr[15:6];
  assign _0038_ = ~ i_wb_adr[5];
  assign _0039_ = i_wb_adr[5:2] == 4'b1011;
  assign _0040_ = ! i_wb_data;
  assign _0041_ = i_wb_adr[4:2] == 3'b100;
  assign _0042_ = mr_index == 1'b1;
  assign _0043_ = mr_index == 2'b10;
  assign _0044_ = md_index == 2'b10;
  assign _0045_ = md_index == 1'b1;
  assign adr_check = _0038_ && adr_check_1;
  assign _0046_ = wack && _0061_;
  assign _0047_ = we && _0062_;
  assign _0048_ = _0039_ && _0063_;
  assign _0049_ = _0048_ && _0040_;
  assign _0050_ = wack && _0071_;
  assign _0051_ = _0050_ && _0072_;
  assign update_kpd = _0051_ && adr_check;
  assign _0052_ = wack && _0041_;
  assign update_esu = _0052_ && adr_check;
  assign _0053_ = p[15] && a[15];
  assign _0054_ = _0053_ && _0064_;
  assign _0055_ = _0065_ && _0066_;
  assign _0056_ = _0055_ && \adder_32bit_0.o_s [15];
  assign _0057_ = p[31] && a[31];
  assign _0058_ = _0057_ && _0067_;
  assign _0059_ = _0068_ && _0069_;
  assign _0060_ = _0059_ && \adder_32bit_0.o_s [31];
  assign _0061_ = ! i_wb_stb;
  assign _0062_ = ! wack;
  assign _0063_ = ! wlRS;
  assign _0064_ = ! \adder_32bit_0.o_s [15];
  assign _0065_ = ! p[15];
  assign _0066_ = ! a[15];
  assign _0067_ = ! \adder_32bit_0.o_s [31];
  assign _0068_ = ! p[31];
  assign _0069_ = ! a[31];
  assign \of_addition[0] = _0054_ || _0056_;
  assign \of_addition[1] = _0058_ || _0060_;
  assign _0070_ = ~ i_wb_we;
  assign _0071_ = ~ i_wb_adr[4];
  assign _0072_ = ~ i_wb_adr[2];
  assign _0073_ = ~ pv;
  assign _0074_ = ~ pv[15];
  assign _0075_ = ~ \err[0] ;
  assign _0076_ = ~ \err[0] [15];
  assign \multiplier_16x16bit_pipelined.i_rst = ~ i_rst;
  assign _0077_ = ~ _0165_;
  assign _0078_ = ~ adr_check_1;
  assign o_valid = ~ rlb;
  assign _0079_ = of[4] | \of_addition[1] ;
  assign _0080_ = of[3] | \of_addition[1] ;
  assign rl[5] = rla | rlb;
  assign rack = _0029_ | _0030_;
  assign _0081_ = wack | rack;
  assign wlRS = wla | wlb;
  always @(posedge i_clk)
    if (i_rst)
      cout <= 1'b0;
    else
      cout <= _0003_;
  always @(posedge i_clk)
    if (i_rst)
      wla <= 1'b0;
    else
      wla <= _0024_;
  always @(posedge i_clk)
    if (i_rst)
      wlb <= 1'b0;
    else
      wlb <= _0025_;
  always @(posedge i_clk)
    if (i_rst)
      state_1 <= 10'b0000000001;
    else
      state_1 <= _0021_;
  always @(posedge i_clk)
    if (i_rst)
      rla <= 1'b0;
    else
      rla <= _0015_;
  always @(posedge i_clk)
    if (i_rst)
      rlb <= 1'b0;
    else
      rlb <= _0016_;
  always @(posedge i_clk)
    if (i_rst)
      of <= 5'b00000;
    else
      of <= _0012_;
  always @(posedge i_clk)
    if (i_rst)
      kpd <= 16'b0000000000000000;
    else
      kpd <= _0009_;
  always @(posedge i_clk)
    if (i_rst)
      p <= 32'd0;
    else
      p <= _0013_;
  always @(posedge i_clk)
    if (i_rst)
      a <= 32'd0;
    else
      a <= _0002_;
  always @(posedge i_clk)
    if (i_rst)
      sigma <= 32'd0;
    else
      sigma <= _0017_;
  always @(posedge i_clk)
    if (i_rst)
      un <= 32'd0;
    else
      un <= _0022_;
  always @(posedge i_clk)
    if (i_rst)
      start <= 1'b0;
    else
      start <= _0019_;
  always @(posedge i_clk)
    if (i_rst)
      mr_index <= 2'b00;
    else
      mr_index <= _0011_;
  always @(posedge i_clk)
    if (i_rst)
      md_index <= 2'b00;
    else
      md_index <= _0010_;
  always @(posedge i_clk)
    if (i_rst)
      \err[0] <= 16'b0000000000000000;
    else
      \err[0] <= _0004_;
  always @(posedge i_clk)
    if (i_rst)
      \err[1] <= 16'b0000000000000000;
    else
      \err[1] <= _0005_;
  always @(posedge i_clk)
    if (i_rst)
      kp <= 16'b0000000000000000;
    else
      kp <= _0008_;
  always @(posedge i_clk)
    if (i_rst)
      ki <= 16'b0000000000000000;
    else
      ki <= _0007_;
  always @(posedge i_clk)
    if (i_rst)
      kd <= 16'b0000000000000000;
    else
      kd <= _0006_;
  always @(posedge i_clk)
    if (i_rst)
      sp <= 16'b0000000000000000;
    else
      sp <= _0018_;
  always @(posedge i_clk)
    if (i_rst)
      pv <= 16'b0000000000000000;
    else
      pv <= _0014_;
  always @(posedge i_clk)
    if (i_rst)
      wack <= 1'b0;
    else
      wack <= _0023_;
  always @(posedge i_clk)
    if (i_rst)
      state_0 <= 1'b0;
    else
      state_0 <= _0020_;
  always @(posedge i_clk)
    if (i_rst)
      RS <= 1'b0;
    else
      RS <= _0001_;
  wire [31:0] fangyuan5;
  assign fangyuan5 = { kp[15], kp[15], kp[15], kp[15], kp[15], kp[15], kp[15], kp[15], kp[15], kp[15], kp[15], kp[15], kp[15], kp[15], kp[15], kp[15], kp };
  wire [351:0] fangyuan6;
  assign fangyuan6 = { ki[15], ki[15], ki[15], ki[15], ki[15], ki[15], ki[15], ki[15], ki[15], ki[15], ki[15], ki[15], ki[15], ki[15], ki[15], ki[15], ki, kd[15], kd[15], kd[15], kd[15], kd[15], kd[15], kd[15], kd[15], kd[15], kd[15], kd[15], kd[15], kd[15], kd[15], kd[15], kd[15], kd, sp[15], sp[15], sp[15], sp[15], sp[15], sp[15], sp[15], sp[15], sp[15], sp[15], sp[15], sp[15], sp[15], sp[15], sp[15], sp[15], sp, pv[15], pv[15], pv[15], pv[15], pv[15], pv[15], pv[15], pv[15], pv[15], pv[15], pv[15], pv[15], pv[15], pv[15], pv[15], pv[15], pv, kpd[15], kpd[15], kpd[15], kpd[15], kpd[15], kpd[15], kpd[15], kpd[15], kpd[15], kpd[15], kpd[15], kpd[15], kpd[15], kpd[15], kpd[15], kpd[15], kpd, \err[0] [15], \err[0] [15], \err[0] [15], \err[0] [15], \err[0] [15], \err[0] [15], \err[0] [15], \err[0] [15], \err[0] [15], \err[0] [15], \err[0] [15], \err[0] [15], \err[0] [15], \err[0] [15], \err[0] [15], \err[0] [15], \err[0] , \err[1] [15], \err[1] [15], \err[1] [15], \err[1] [15], \err[1] [15], \err[1] [15], \err[1] [15], \err[1] [15], \err[1] [15], \err[1] [15], \err[1] [15], \err[1] [15], \err[1] [15], \err[1] [15], \err[1] [15], \err[1] [15], \err[1] , un, sigma, 27'b000000000000000000000000000, of, 16'b0000000000000000, 16'b0000000000000000 };
  wire [10:0] fangyuan7;
  assign fangyuan7 = { _0095_, _0094_, _0093_, _0092_, _0091_, _0090_, _0089_, _0088_, _0087_, _0086_, _0031_ };

  always @(fangyuan5 or fangyuan6 or fangyuan7) begin
    casez (fangyuan7)
      11'b??????????1 :
        _0000_ = fangyuan6 [31:0] ;
      11'b?????????1? :
        _0000_ = fangyuan6 [63:32] ;
      11'b????????1?? :
        _0000_ = fangyuan6 [95:64] ;
      11'b???????1??? :
        _0000_ = fangyuan6 [127:96] ;
      11'b??????1???? :
        _0000_ = fangyuan6 [159:128] ;
      11'b?????1????? :
        _0000_ = fangyuan6 [191:160] ;
      11'b????1?????? :
        _0000_ = fangyuan6 [223:192] ;
      11'b???1??????? :
        _0000_ = fangyuan6 [255:224] ;
      11'b??1???????? :
        _0000_ = fangyuan6 [287:256] ;
      11'b?1????????? :
        _0000_ = fangyuan6 [319:288] ;
      11'b1?????????? :
        _0000_ = fangyuan6 [351:320] ;
      default:
        _0000_ = fangyuan5 ;
    endcase
  end
  assign _0082_ = i_wb_adr[5:2] == 4'b1111;
  assign _0083_ = i_wb_adr[5:2] == 4'b1110;
  assign _0084_ = i_wb_adr[5:2] == 4'b1101;
  assign _0085_ = i_wb_adr[5:2] == 4'b1100;
  assign _0086_ = i_wb_adr[5:2] == 4'b1010;
  assign _0087_ = i_wb_adr[5:2] == 4'b1001;
  assign _0088_ = i_wb_adr[5:2] == 4'b1000;
  assign _0089_ = i_wb_adr[5:2] == 3'b111;
  assign _0090_ = i_wb_adr[5:2] == 3'b110;
  assign _0091_ = i_wb_adr[5:2] == 3'b101;
  assign _0092_ = i_wb_adr[5:2] == 3'b100;
  assign _0093_ = i_wb_adr[5:2] == 2'b11;
  assign _0094_ = i_wb_adr[5:2] == 2'b10;
  assign _0095_ = i_wb_adr[5:2] == 1'b1;
  wire [1:0] fangyuan8;
  assign fangyuan8 = { _0099_, _0079_ };
  wire [1:0] fangyuan9;
  assign fangyuan9 = { _0100_, _0096_ };

  always @(of[4] or fangyuan8 or fangyuan9) begin
    casez (fangyuan9)
      2'b?1 :
        _0012_[4] = fangyuan8 [0:0] ;
      2'b1? :
        _0012_[4] = fangyuan8 [1:1] ;
      default:
        _0012_[4] = of[4] ;
    endcase
  end
  assign _0096_ = state_1 == 8'b10000000;
  assign _0097_ = RS ? 1'b0 : of[4];
  assign _0098_ = update_esu ? of[4] : _0097_;
  assign _0099_ = update_kpd ? of[4] : _0098_;
  assign _0100_ = state_1 == 1'b1;
  wire [2:0] fangyuan10;
  assign fangyuan10 = { _0105_, _0079_, _0080_ };
  wire [2:0] fangyuan11;
  assign fangyuan11 = { _0100_, _0096_, _0032_ };

  always @(of[3] or fangyuan10 or fangyuan11) begin
    casez (fangyuan11)
      3'b??1 :
        _0012_[3] = fangyuan10 [0:0] ;
      3'b?1? :
        _0012_[3] = fangyuan10 [1:1] ;
      3'b1?? :
        _0012_[3] = fangyuan10 [2:2] ;
      default:
        _0012_[3] = of[3] ;
    endcase
  end
  assign _0101_ = state_1 == 10'b1000000000;
  assign _0102_ = state_1 == 9'b100000000;
  assign _0103_ = RS ? 1'b0 : of[3];
  assign _0104_ = update_esu ? of[3] : _0103_;
  assign _0105_ = update_kpd ? of[3] : _0104_;
  wire [1:0] fangyuan12;
  assign fangyuan12 = { _0109_, of[1] };
  wire [1:0] fangyuan13;
  assign fangyuan13 = { _0100_, _0106_ };

  always @(of[2] or fangyuan12 or fangyuan13) begin
    casez (fangyuan13)
      2'b?1 :
        _0012_[2] = fangyuan12 [0:0] ;
      2'b1? :
        _0012_[2] = fangyuan12 [1:1] ;
      default:
        _0012_[2] = of[2] ;
    endcase
  end
  assign _0106_ = state_1 == 5'b10000;
  assign _0107_ = RS ? 1'b0 : of[2];
  assign _0108_ = update_esu ? of[2] : _0107_;
  assign _0109_ = update_kpd ? of[2] : _0108_;
  wire [1:0] fangyuan14;
  assign fangyuan14 = { _0112_, \of_addition[0] };
  wire [1:0] fangyuan15;
  assign fangyuan15 = { _0100_, _0106_ };

  always @(of[1] or fangyuan14 or fangyuan15) begin
    casez (fangyuan15)
      2'b?1 :
        _0012_[1] = fangyuan14 [0:0] ;
      2'b1? :
        _0012_[1] = fangyuan14 [1:1] ;
      default:
        _0012_[1] = of[1] ;
    endcase
  end
  assign _0110_ = RS ? 1'b0 : of[1];
  assign _0111_ = update_esu ? of[1] : _0110_;
  assign _0112_ = update_kpd ? of[1] : _0111_;
  wire [1:0] fangyuan16;
  assign fangyuan16 = { _0116_, \of_addition[0] };
  wire [1:0] fangyuan17;
  assign fangyuan17 = { _0100_, _0113_ };

  always @(of[0] or fangyuan16 or fangyuan17) begin
    casez (fangyuan17)
      2'b?1 :
        _0012_[0] = fangyuan16 [0:0] ;
      2'b1? :
        _0012_[0] = fangyuan16 [1:1] ;
      default:
        _0012_[0] = of[0] ;
    endcase
  end
  assign _0113_ = state_1 == 3'b100;
  assign _0114_ = RS ? 1'b0 : of[0];
  assign _0115_ = update_esu ? of[0] : _0114_;
  assign _0116_ = update_kpd ? of[0] : _0115_;
  assign _0005_ = _0117_ ? \adder_32bit_0.o_s [15:0] : \err[1] ;
  assign _0117_ = state_1 == 6'b100000;
  wire [31:0] fangyuan18;
  assign fangyuan18 = { _0120_, \adder_32bit_0.o_s [15:0] };
  wire [1:0] fangyuan19;
  assign fangyuan19 = { _0100_, _0106_ };

  always @(\err[0] or fangyuan18 or fangyuan19) begin
    casez (fangyuan19)
      2'b?1 :
        _0004_ = fangyuan18 [15:0] ;
      2'b1? :
        _0004_ = fangyuan18 [31:16] ;
      default:
        _0004_ = \err[0] ;
    endcase
  end
  assign _0118_ = RS ? 16'b0000000000000000 : \err[0] ;
  assign _0119_ = update_esu ? \err[0] : _0118_;
  assign _0120_ = update_kpd ? \err[0] : _0119_;
  wire [2:0] fangyuan20;
  assign fangyuan20 = { _0106_, _0117_, _0121_ };

  always @(md_index or fangyuan20) begin
    casez (fangyuan20)
      3'b??1 :
        _0010_ = 2'b00 ;
      3'b?1? :
        _0010_ = 2'b10 ;
      3'b1?? :
        _0010_ = 2'b01 ;
      default:
        _0010_ = md_index ;
    endcase
  end
  assign _0121_ = state_1 == 7'b1000000;
  wire [2:0] fangyuan21;
  assign fangyuan21 = { _0106_, _0117_, _0121_ };

  always @(mr_index or fangyuan21) begin
    casez (fangyuan21)
      3'b??1 :
        _0011_ = 2'b00 ;
      3'b?1? :
        _0011_ = 2'b10 ;
      3'b1?? :
        _0011_ = 2'b01 ;
      default:
        _0011_ = mr_index ;
    endcase
  end
  wire [1:0] fangyuan22;
  assign fangyuan22 = { _0122_, _0121_ };

  always @(start or fangyuan22) begin
    casez (fangyuan22)
      2'b?1 :
        _0019_ = 1'b0 ;
      2'b1? :
        _0019_ = 1'b1 ;
      default:
        _0019_ = start ;
    endcase
  end
  assign _0122_ = state_1 == 4'b1000;
  wire [63:0] fangyuan23;
  assign fangyuan23 = { _0125_, \adder_32bit_0.o_s };
  wire [1:0] fangyuan24;
  assign fangyuan24 = { _0100_, _0101_ };

  always @(un or fangyuan23 or fangyuan24) begin
    casez (fangyuan24)
      2'b?1 :
        _0022_ = fangyuan23 [31:0] ;
      2'b1? :
        _0022_ = fangyuan23 [63:32] ;
      default:
        _0022_ = un ;
    endcase
  end
  assign _0123_ = RS ? 32'd0 : un;
  assign _0124_ = update_esu ? un : _0123_;
  assign _0125_ = update_kpd ? un : _0124_;
  wire [63:0] fangyuan25;
  assign fangyuan25 = { _0128_, \adder_32bit_0.o_s };
  wire [1:0] fangyuan26;
  assign fangyuan26 = { _0100_, _0096_ };

  always @(sigma or fangyuan25 or fangyuan26) begin
    casez (fangyuan26)
      2'b?1 :
        _0017_ = fangyuan25 [31:0] ;
      2'b1? :
        _0017_ = fangyuan25 [63:32] ;
      default:
        _0017_ = sigma ;
    endcase
  end
  assign _0126_ = RS ? 32'd0 : sigma;
  assign _0127_ = update_esu ? sigma : _0126_;
  assign _0128_ = update_kpd ? sigma : _0127_;
  wire [159:0] fangyuan27;
  assign fangyuan27 = { kd[15], kd[15], kd[15], kd[15], kd[15], kd[15], kd[15], kd[15], kd[15], kd[15], kd[15], kd[15], kd[15], kd[15], kd[15], kd[15], kd, _0074_, _0074_, _0074_, _0074_, _0074_, _0074_, _0074_, _0074_, _0074_, _0074_, _0074_, _0074_, _0074_, _0074_, _0074_, _0074_, _0073_, 16'b0000000000000000, 16'b0000000000000001, sigma, \adder_32bit_0.o_s };
  wire [4:0] fangyuan28;
  assign fangyuan28 = { _0129_, _0122_, _0106_, _0121_, _0033_ };

  always @(a or fangyuan27 or fangyuan28) begin
    casez (fangyuan28)
      5'b????1 :
        _0002_ = fangyuan27 [31:0] ;
      5'b???1? :
        _0002_ = fangyuan27 [63:32] ;
      5'b??1?? :
        _0002_ = fangyuan27 [95:64] ;
      5'b?1??? :
        _0002_ = fangyuan27 [127:96] ;
      5'b1???? :
        _0002_ = fangyuan27 [159:128] ;
      default:
        _0002_ = a ;
    endcase
  end
  assign _0129_ = state_1 == 2'b10;
  wire [127:0] fangyuan29;
  assign fangyuan29 = { kp[15], kp[15], kp[15], kp[15], kp[15], kp[15], kp[15], kp[15], kp[15], kp[15], kp[15], kp[15], kp[15], kp[15], kp[15], kp[15], kp, sp[15], sp[15], sp[15], sp[15], sp[15], sp[15], sp[15], sp[15], sp[15], sp[15], sp[15], sp[15], sp[15], sp[15], sp[15], sp[15], sp, _0076_, _0076_, _0076_, _0076_, _0076_, _0076_, _0076_, _0076_, _0076_, _0076_, _0076_, _0076_, _0076_, _0076_, _0076_, _0076_, _0075_, \multiplier_16x16bit_pipelined.adder_32bit.o_s [31:1], \multiplier_16x16bit_pipelined.adder_32bit.operator_A_0.P };
  wire [3:0] fangyuan30;
  assign fangyuan30 = { _0129_, _0122_, _0106_, _0034_ };

  always @(p or fangyuan29 or fangyuan30) begin
    casez (fangyuan30)
      4'b???1 :
        _0013_ = fangyuan29 [31:0] ;
      4'b??1? :
        _0013_ = fangyuan29 [63:32] ;
      4'b?1?? :
        _0013_ = fangyuan29 [95:64] ;
      4'b1??? :
        _0013_ = fangyuan29 [127:96] ;
      default:
        _0013_ = p ;
    endcase
  end
  assign _0009_ = _0113_ ? \adder_32bit_0.o_s [15:0] : kpd;
  wire [1:0] fangyuan31;
  assign fangyuan31 = { _0131_, 1'b0 };
  wire [1:0] fangyuan32;
  assign fangyuan32 = { _0100_, _0101_ };

  always @(rlb or fangyuan31 or fangyuan32) begin
    casez (fangyuan32)
      2'b?1 :
        _0016_ = fangyuan31 [0:0] ;
      2'b1? :
        _0016_ = fangyuan31 [1:1] ;
      default:
        _0016_ = rlb ;
    endcase
  end
  assign _0130_ = update_esu ? 1'b1 : rlb;
  assign _0131_ = update_kpd ? rlb : _0130_;
  wire [1:0] fangyuan33;
  assign fangyuan33 = { _0132_, 1'b0 };
  wire [1:0] fangyuan34;
  assign fangyuan34 = { _0100_, _0113_ };

  always @(rla or fangyuan33 or fangyuan34) begin
    casez (fangyuan34)
      2'b?1 :
        _0015_ = fangyuan33 [0:0] ;
      2'b1? :
        _0015_ = fangyuan33 [1:1] ;
      default:
        _0015_ = rla ;
    endcase
  end
  assign _0132_ = update_kpd ? 1'b1 : rla;
  wire [89:0] fangyuan35;
  assign fangyuan35 = { _0134_, 16'b0000000100000001, 16'b0000000010000000, 16'b0100000000100000, 16'b0001000000001000, 16'b0000000000000001 };
  wire [8:0] fangyuan36;
  assign fangyuan36 = { _0100_, _0129_, _0122_, _0106_, _0117_, _0121_, _0096_, _0102_, _0035_ };

  always @(state_1 or fangyuan35 or fangyuan36) begin
    casez (fangyuan36)
      9'b????????1 :
        _0021_ = fangyuan35 [9:0] ;
      9'b???????1? :
        _0021_ = fangyuan35 [19:10] ;
      9'b??????1?? :
        _0021_ = fangyuan35 [29:20] ;
      9'b?????1??? :
        _0021_ = fangyuan35 [39:30] ;
      9'b????1???? :
        _0021_ = fangyuan35 [49:40] ;
      9'b???1????? :
        _0021_ = fangyuan35 [59:50] ;
      9'b??1?????? :
        _0021_ = fangyuan35 [69:60] ;
      9'b?1??????? :
        _0021_ = fangyuan35 [79:70] ;
      9'b1???????? :
        _0021_ = fangyuan35 [89:80] ;
      default:
        _0021_ = state_1 ;
    endcase
  end
  assign _0133_ = update_esu ? 10'b0000001000 : state_1;
  assign _0134_ = update_kpd ? 10'b0000000010 : _0133_;
  wire [1:0] fangyuan37;
  assign fangyuan37 = { _0136_, 1'b0 };
  wire [1:0] fangyuan38;
  assign fangyuan38 = { _0100_, _0101_ };

  always @(wlb or fangyuan37 or fangyuan38) begin
    casez (fangyuan38)
      2'b?1 :
        _0025_ = fangyuan37 [0:0] ;
      2'b1? :
        _0025_ = fangyuan37 [1:1] ;
      default:
        _0025_ = wlb ;
    endcase
  end
  assign _0135_ = update_esu ? 1'b1 : wlb;
  assign _0136_ = update_kpd ? wlb : _0135_;
  wire [1:0] fangyuan39;
  assign fangyuan39 = { _0138_, 1'b0 };
  wire [1:0] fangyuan40;
  assign fangyuan40 = { _0100_, _0035_ };

  always @(wla or fangyuan39 or fangyuan40) begin
    casez (fangyuan40)
      2'b?1 :
        _0024_ = fangyuan39 [0:0] ;
      2'b1? :
        _0024_ = fangyuan39 [1:1] ;
      default:
        _0024_ = wla ;
    endcase
  end
  assign _0137_ = update_esu ? 1'b1 : wla;
  assign _0138_ = update_kpd ? 1'b1 : _0137_;
  wire [1:0] fangyuan41;
  assign fangyuan41 = { _0122_, _0106_ };

  always @(cout or fangyuan41) begin
    casez (fangyuan41)
      2'b?1 :
        _0003_ = 1'b0 ;
      2'b1? :
        _0003_ = 1'b1 ;
      default:
        _0003_ = cout ;
    endcase
  end
  assign _0139_ = adr_check ? 1'b0 : _0049_;
  assign _0001_ = state_0 ? _0139_ : 1'b0;
  assign _0141_ = adr_check ? _0140_ : 1'b0;
  wire [1:0] fangyuan42;
  assign fangyuan42 = { _0047_, _0141_ };
  wire [1:0] fangyuan43;
  assign fangyuan43 = { _0142_, state_0 };

  always @(1'b0 or fangyuan42 or fangyuan43) begin
    casez (fangyuan43)
      2'b?1 :
        _0020_ = fangyuan42 [0:0] ;
      2'b1? :
        _0020_ = fangyuan42 [1:1] ;
      default:
        _0020_ = 1'b0 ;
    endcase
  end
  assign _0142_ = ~ state_0;
  assign _0143_ = _0046_ ? 1'b0 : wack;
  assign _0144_ = _0140_ ? _0143_ : 1'b1;
  assign _0145_ = adr_check ? _0144_ : 1'b1;
  assign _0023_ = state_0 ? _0145_ : _0143_;
  assign _0146_ = _0041_ ? i_wb_data[15:0] : pv;
  assign _0147_ = _0140_ ? pv : _0146_;
  assign _0148_ = adr_check ? _0147_ : pv;
  assign _0014_ = state_0 ? _0148_ : pv;
  assign _0149_ = _0150_ ? i_wb_data[15:0] : sp;
  assign _0150_ = i_wb_adr[4:2] == 2'b11;
  assign _0151_ = _0140_ ? sp : _0149_;
  assign _0152_ = adr_check ? _0151_ : sp;
  assign _0018_ = state_0 ? _0152_ : sp;
  assign _0153_ = _0154_ ? i_wb_data[15:0] : kd;
  assign _0154_ = i_wb_adr[4:2] == 2'b10;
  assign _0155_ = _0140_ ? kd : _0153_;
  assign _0156_ = adr_check ? _0155_ : kd;
  assign _0006_ = state_0 ? _0156_ : kd;
  assign _0157_ = _0158_ ? i_wb_data[15:0] : ki;
  assign _0158_ = i_wb_adr[4:2] == 1'b1;
  assign _0159_ = _0140_ ? ki : _0157_;
  assign _0160_ = adr_check ? _0159_ : ki;
  assign _0007_ = state_0 ? _0160_ : ki;
  assign _0161_ = _0162_ ? i_wb_data[15:0] : kp;
  assign _0162_ = ! i_wb_adr[4:2];
  assign _0163_ = _0140_ ? kp : _0161_;
  assign _0164_ = adr_check ? _0163_ : kp;
  assign _0008_ = state_0 ? _0164_ : kp;
  wire [7:0] fangyuan44;
  assign fangyuan44 = { wla, wla, wla, wlb, wlb, 3'b000 };

  assign _0140_ = fangyuan44[$signed(_0036_) +: 1];
  wire [15:0] fangyuan45;
  assign fangyuan45 = { 5'b00000, rla, rlb, rlb, rlb, rlb, rl[5], 5'b00000 };

  assign _0165_ = fangyuan45[$signed(_0037_) +: 1];
  assign \adder_32bit_0.o_s [0] = \adder_32bit_0.operator_A_0.P ^ cout;
  assign \adder_32bit_0.o_s [1] = \adder_32bit_0.operator_A_1.P ^ \adder_32bit_0.operator_C_stage_1_0.Go ;
  assign \adder_32bit_0.o_s [2] = \adder_32bit_0.operator_A_2.P ^ \adder_32bit_0.operator_C_stage_6_0.Go ;
  assign \adder_32bit_0.o_s [3] = \adder_32bit_0.operator_A_3.P ^ \adder_32bit_0.operator_C_stage_2_1.Go ;
  assign \adder_32bit_0.o_s [4] = \adder_32bit_0.operator_A_4.P ^ \adder_32bit_0.operator_C_stage_6_1.Go ;
  assign \adder_32bit_0.o_s [5] = \adder_32bit_0.operator_A_5.P ^ \adder_32bit_0.operator_C_stage_3_2.Go ;
  assign \adder_32bit_0.o_s [6] = \adder_32bit_0.operator_A_6.P ^ \adder_32bit_0.operator_C_stage_6_2.Go ;
  assign \adder_32bit_0.o_s [7] = \adder_32bit_0.operator_A_7.P ^ \adder_32bit_0.operator_C_stage_3_3.Go ;
  assign \adder_32bit_0.o_s [8] = \adder_32bit_0.operator_A_8.P ^ \adder_32bit_0.operator_C_stage_6_3.Go ;
  assign \adder_32bit_0.o_s [9] = \adder_32bit_0.operator_A_9.P ^ \adder_32bit_0.operator_C_stage_4_4.Go ;
  assign \adder_32bit_0.o_s [10] = \adder_32bit_0.operator_A_10.P ^ \adder_32bit_0.operator_C_stage_6_4.Go ;
  assign \adder_32bit_0.o_s [11] = \adder_32bit_0.operator_A_11.P ^ \adder_32bit_0.operator_C_stage_4_5.Go ;
  assign \adder_32bit_0.o_s [12] = \adder_32bit_0.operator_A_12.P ^ \adder_32bit_0.operator_C_stage_6_5.Go ;
  assign \adder_32bit_0.o_s [13] = \adder_32bit_0.operator_A_13.P ^ \adder_32bit_0.operator_C_stage_4_6.Go ;
  assign \adder_32bit_0.o_s [14] = \adder_32bit_0.operator_A_14.P ^ \adder_32bit_0.operator_C_stage_6_6.Go ;
  assign \adder_32bit_0.o_s [15] = \adder_32bit_0.operator_A_15.P ^ \adder_32bit_0.operator_C_stage_4_7.Go ;
  assign \adder_32bit_0.o_s [16] = \adder_32bit_0.operator_A_16.P ^ \adder_32bit_0.operator_C_stage_6_7.Go ;
  assign \adder_32bit_0.o_s [17] = \adder_32bit_0.operator_A_17.P ^ \adder_32bit_0.operator_C_stage_5_8.Go ;
  assign \adder_32bit_0.o_s [18] = \adder_32bit_0.operator_A_18.P ^ \adder_32bit_0.operator_C_stage_6_8.Go ;
  assign \adder_32bit_0.o_s [19] = \adder_32bit_0.operator_A_19.P ^ \adder_32bit_0.operator_C_stage_5_9.Go ;
  assign \adder_32bit_0.o_s [20] = \adder_32bit_0.operator_A_20.P ^ \adder_32bit_0.operator_C_stage_6_9.Go ;
  assign \adder_32bit_0.o_s [21] = \adder_32bit_0.operator_A_21.P ^ \adder_32bit_0.operator_C_stage_5_10.Go ;
  assign \adder_32bit_0.o_s [22] = \adder_32bit_0.operator_A_22.P ^ \adder_32bit_0.operator_C_stage_6_10.Go ;
  assign \adder_32bit_0.o_s [23] = \adder_32bit_0.operator_A_23.P ^ \adder_32bit_0.operator_C_stage_5_11.Go ;
  assign \adder_32bit_0.o_s [24] = \adder_32bit_0.operator_A_24.P ^ \adder_32bit_0.operator_C_stage_6_11.Go ;
  assign \adder_32bit_0.o_s [25] = \adder_32bit_0.operator_A_25.P ^ \adder_32bit_0.operator_C_stage_5_12.Go ;
  assign \adder_32bit_0.o_s [26] = \adder_32bit_0.operator_A_26.P ^ \adder_32bit_0.operator_C_stage_6_12.Go ;
  assign \adder_32bit_0.o_s [27] = \adder_32bit_0.operator_A_27.P ^ \adder_32bit_0.operator_C_stage_5_13.Go ;
  assign \adder_32bit_0.o_s [28] = \adder_32bit_0.operator_A_28.P ^ \adder_32bit_0.operator_C_stage_6_13.Go ;
  assign \adder_32bit_0.o_s [29] = \adder_32bit_0.operator_A_29.P ^ \adder_32bit_0.operator_C_stage_5_14.Go ;
  assign \adder_32bit_0.o_s [30] = \adder_32bit_0.operator_A_30.P ^ \adder_32bit_0.operator_C_stage_6_14.Go ;
  assign \adder_32bit_0.o_s [31] = \adder_32bit_0.operator_A_31.P ^ \adder_32bit_0.operator_C_stage_5_15.Go ;
  assign \adder_32bit_0.operator_A_0.G = a[0] & p[0];
  assign \adder_32bit_0.operator_A_0.P = a[0] ^ p[0];
  assign \adder_32bit_0.operator_A_1.G = a[1] & p[1];
  assign \adder_32bit_0.operator_A_1.P = a[1] ^ p[1];
  assign \adder_32bit_0.operator_A_10.G = a[10] & p[10];
  assign \adder_32bit_0.operator_A_10.P = a[10] ^ p[10];
  assign \adder_32bit_0.operator_A_11.G = a[11] & p[11];
  assign \adder_32bit_0.operator_A_11.P = a[11] ^ p[11];
  assign \adder_32bit_0.operator_A_12.G = a[12] & p[12];
  assign \adder_32bit_0.operator_A_12.P = a[12] ^ p[12];
  assign \adder_32bit_0.operator_A_13.G = a[13] & p[13];
  assign \adder_32bit_0.operator_A_13.P = a[13] ^ p[13];
  assign \adder_32bit_0.operator_A_14.G = a[14] & p[14];
  assign \adder_32bit_0.operator_A_14.P = a[14] ^ p[14];
  assign \adder_32bit_0.operator_A_15.G = a[15] & p[15];
  assign \adder_32bit_0.operator_A_15.P = a[15] ^ p[15];
  assign \adder_32bit_0.operator_A_16.G = a[16] & p[16];
  assign \adder_32bit_0.operator_A_16.P = a[16] ^ p[16];
  assign \adder_32bit_0.operator_A_17.G = a[17] & p[17];
  assign \adder_32bit_0.operator_A_17.P = a[17] ^ p[17];
  assign \adder_32bit_0.operator_A_18.G = a[18] & p[18];
  assign \adder_32bit_0.operator_A_18.P = a[18] ^ p[18];
  assign \adder_32bit_0.operator_A_19.G = a[19] & p[19];
  assign \adder_32bit_0.operator_A_19.P = a[19] ^ p[19];
  assign \adder_32bit_0.operator_A_2.G = a[2] & p[2];
  assign \adder_32bit_0.operator_A_2.P = a[2] ^ p[2];
  assign \adder_32bit_0.operator_A_20.G = a[20] & p[20];
  assign \adder_32bit_0.operator_A_20.P = a[20] ^ p[20];
  assign \adder_32bit_0.operator_A_21.G = a[21] & p[21];
  assign \adder_32bit_0.operator_A_21.P = a[21] ^ p[21];
  assign \adder_32bit_0.operator_A_22.G = a[22] & p[22];
  assign \adder_32bit_0.operator_A_22.P = a[22] ^ p[22];
  assign \adder_32bit_0.operator_A_23.G = a[23] & p[23];
  assign \adder_32bit_0.operator_A_23.P = a[23] ^ p[23];
  assign \adder_32bit_0.operator_A_24.G = a[24] & p[24];
  assign \adder_32bit_0.operator_A_24.P = a[24] ^ p[24];
  assign \adder_32bit_0.operator_A_25.G = a[25] & p[25];
  assign \adder_32bit_0.operator_A_25.P = a[25] ^ p[25];
  assign \adder_32bit_0.operator_A_26.G = a[26] & p[26];
  assign \adder_32bit_0.operator_A_26.P = a[26] ^ p[26];
  assign \adder_32bit_0.operator_A_27.G = a[27] & p[27];
  assign \adder_32bit_0.operator_A_27.P = a[27] ^ p[27];
  assign \adder_32bit_0.operator_A_28.G = a[28] & p[28];
  assign \adder_32bit_0.operator_A_28.P = a[28] ^ p[28];
  assign \adder_32bit_0.operator_A_29.G = a[29] & p[29];
  assign \adder_32bit_0.operator_A_29.P = a[29] ^ p[29];
  assign \adder_32bit_0.operator_A_3.G = a[3] & p[3];
  assign \adder_32bit_0.operator_A_3.P = a[3] ^ p[3];
  assign \adder_32bit_0.operator_A_30.G = a[30] & p[30];
  assign \adder_32bit_0.operator_A_30.P = a[30] ^ p[30];
  assign \adder_32bit_0.operator_A_31.P = a[31] ^ p[31];
  assign \adder_32bit_0.operator_A_4.G = a[4] & p[4];
  assign \adder_32bit_0.operator_A_4.P = a[4] ^ p[4];
  assign \adder_32bit_0.operator_A_5.G = a[5] & p[5];
  assign \adder_32bit_0.operator_A_5.P = a[5] ^ p[5];
  assign \adder_32bit_0.operator_A_6.G = a[6] & p[6];
  assign \adder_32bit_0.operator_A_6.P = a[6] ^ p[6];
  assign \adder_32bit_0.operator_A_7.G = a[7] & p[7];
  assign \adder_32bit_0.operator_A_7.P = a[7] ^ p[7];
  assign \adder_32bit_0.operator_A_8.G = a[8] & p[8];
  assign \adder_32bit_0.operator_A_8.P = a[8] ^ p[8];
  assign \adder_32bit_0.operator_A_9.G = a[9] & p[9];
  assign \adder_32bit_0.operator_A_9.P = a[9] ^ p[9];
  assign \adder_32bit_0.operator_B_stage_1_1.Po = \adder_32bit_0.operator_A_2.P & \adder_32bit_0.operator_A_1.P ;
  assign _0166_ = \adder_32bit_0.operator_A_2.P & \adder_32bit_0.operator_A_1.G ;
  assign \adder_32bit_0.operator_B_stage_1_1.Go = \adder_32bit_0.operator_A_2.G | _0166_;
  assign \adder_32bit_0.operator_B_stage_1_10.Po = \adder_32bit_0.operator_A_20.P & \adder_32bit_0.operator_A_19.P ;
  assign _0167_ = \adder_32bit_0.operator_A_20.P & \adder_32bit_0.operator_A_19.G ;
  assign \adder_32bit_0.operator_B_stage_1_10.Go = \adder_32bit_0.operator_A_20.G | _0167_;
  assign \adder_32bit_0.operator_B_stage_1_11.Po = \adder_32bit_0.operator_A_22.P & \adder_32bit_0.operator_A_21.P ;
  assign _0168_ = \adder_32bit_0.operator_A_22.P & \adder_32bit_0.operator_A_21.G ;
  assign \adder_32bit_0.operator_B_stage_1_11.Go = \adder_32bit_0.operator_A_22.G | _0168_;
  assign \adder_32bit_0.operator_B_stage_1_12.Po = \adder_32bit_0.operator_A_24.P & \adder_32bit_0.operator_A_23.P ;
  assign _0169_ = \adder_32bit_0.operator_A_24.P & \adder_32bit_0.operator_A_23.G ;
  assign \adder_32bit_0.operator_B_stage_1_12.Go = \adder_32bit_0.operator_A_24.G | _0169_;
  assign \adder_32bit_0.operator_B_stage_1_13.Po = \adder_32bit_0.operator_A_26.P & \adder_32bit_0.operator_A_25.P ;
  assign _0170_ = \adder_32bit_0.operator_A_26.P & \adder_32bit_0.operator_A_25.G ;
  assign \adder_32bit_0.operator_B_stage_1_13.Go = \adder_32bit_0.operator_A_26.G | _0170_;
  assign \adder_32bit_0.operator_B_stage_1_14.Po = \adder_32bit_0.operator_A_28.P & \adder_32bit_0.operator_A_27.P ;
  assign _0171_ = \adder_32bit_0.operator_A_28.P & \adder_32bit_0.operator_A_27.G ;
  assign \adder_32bit_0.operator_B_stage_1_14.Go = \adder_32bit_0.operator_A_28.G | _0171_;
  assign \adder_32bit_0.operator_B_stage_1_15.Po = \adder_32bit_0.operator_A_30.P & \adder_32bit_0.operator_A_29.P ;
  assign _0172_ = \adder_32bit_0.operator_A_30.P & \adder_32bit_0.operator_A_29.G ;
  assign \adder_32bit_0.operator_B_stage_1_15.Go = \adder_32bit_0.operator_A_30.G | _0172_;
  assign \adder_32bit_0.operator_B_stage_1_2.Po = \adder_32bit_0.operator_A_4.P & \adder_32bit_0.operator_A_3.P ;
  assign _0173_ = \adder_32bit_0.operator_A_4.P & \adder_32bit_0.operator_A_3.G ;
  assign \adder_32bit_0.operator_B_stage_1_2.Go = \adder_32bit_0.operator_A_4.G | _0173_;
  assign \adder_32bit_0.operator_B_stage_1_3.Po = \adder_32bit_0.operator_A_6.P & \adder_32bit_0.operator_A_5.P ;
  assign _0174_ = \adder_32bit_0.operator_A_6.P & \adder_32bit_0.operator_A_5.G ;
  assign \adder_32bit_0.operator_B_stage_1_3.Go = \adder_32bit_0.operator_A_6.G | _0174_;
  assign \adder_32bit_0.operator_B_stage_1_4.Po = \adder_32bit_0.operator_A_8.P & \adder_32bit_0.operator_A_7.P ;
  assign _0175_ = \adder_32bit_0.operator_A_8.P & \adder_32bit_0.operator_A_7.G ;
  assign \adder_32bit_0.operator_B_stage_1_4.Go = \adder_32bit_0.operator_A_8.G | _0175_;
  assign \adder_32bit_0.operator_B_stage_1_5.Po = \adder_32bit_0.operator_A_10.P & \adder_32bit_0.operator_A_9.P ;
  assign _0176_ = \adder_32bit_0.operator_A_10.P & \adder_32bit_0.operator_A_9.G ;
  assign \adder_32bit_0.operator_B_stage_1_5.Go = \adder_32bit_0.operator_A_10.G | _0176_;
  assign \adder_32bit_0.operator_B_stage_1_6.Po = \adder_32bit_0.operator_A_12.P & \adder_32bit_0.operator_A_11.P ;
  assign _0177_ = \adder_32bit_0.operator_A_12.P & \adder_32bit_0.operator_A_11.G ;
  assign \adder_32bit_0.operator_B_stage_1_6.Go = \adder_32bit_0.operator_A_12.G | _0177_;
  assign \adder_32bit_0.operator_B_stage_1_7.Po = \adder_32bit_0.operator_A_14.P & \adder_32bit_0.operator_A_13.P ;
  assign _0178_ = \adder_32bit_0.operator_A_14.P & \adder_32bit_0.operator_A_13.G ;
  assign \adder_32bit_0.operator_B_stage_1_7.Go = \adder_32bit_0.operator_A_14.G | _0178_;
  assign \adder_32bit_0.operator_B_stage_1_8.Po = \adder_32bit_0.operator_A_16.P & \adder_32bit_0.operator_A_15.P ;
  assign _0179_ = \adder_32bit_0.operator_A_16.P & \adder_32bit_0.operator_A_15.G ;
  assign \adder_32bit_0.operator_B_stage_1_8.Go = \adder_32bit_0.operator_A_16.G | _0179_;
  assign \adder_32bit_0.operator_B_stage_1_9.Po = \adder_32bit_0.operator_A_18.P & \adder_32bit_0.operator_A_17.P ;
  assign _0180_ = \adder_32bit_0.operator_A_18.P & \adder_32bit_0.operator_A_17.G ;
  assign \adder_32bit_0.operator_B_stage_1_9.Go = \adder_32bit_0.operator_A_18.G | _0180_;
  assign \adder_32bit_0.operator_B_stage_2_10.Po = \adder_32bit_0.operator_B_stage_1_10.Po & \adder_32bit_0.operator_B_stage_1_9.Po ;
  assign _0181_ = \adder_32bit_0.operator_B_stage_1_10.Po & \adder_32bit_0.operator_B_stage_1_9.Go ;
  assign \adder_32bit_0.operator_B_stage_2_10.Go = \adder_32bit_0.operator_B_stage_1_10.Go | _0181_;
  assign \adder_32bit_0.operator_B_stage_2_11.Po = \adder_32bit_0.operator_B_stage_1_11.Po & \adder_32bit_0.operator_B_stage_1_10.Po ;
  assign _0182_ = \adder_32bit_0.operator_B_stage_1_11.Po & \adder_32bit_0.operator_B_stage_1_10.Go ;
  assign \adder_32bit_0.operator_B_stage_2_11.Go = \adder_32bit_0.operator_B_stage_1_11.Go | _0182_;
  assign \adder_32bit_0.operator_B_stage_2_12.Po = \adder_32bit_0.operator_B_stage_1_12.Po & \adder_32bit_0.operator_B_stage_1_11.Po ;
  assign _0183_ = \adder_32bit_0.operator_B_stage_1_12.Po & \adder_32bit_0.operator_B_stage_1_11.Go ;
  assign \adder_32bit_0.operator_B_stage_2_12.Go = \adder_32bit_0.operator_B_stage_1_12.Go | _0183_;
  assign \adder_32bit_0.operator_B_stage_2_13.Po = \adder_32bit_0.operator_B_stage_1_13.Po & \adder_32bit_0.operator_B_stage_1_12.Po ;
  assign _0184_ = \adder_32bit_0.operator_B_stage_1_13.Po & \adder_32bit_0.operator_B_stage_1_12.Go ;
  assign \adder_32bit_0.operator_B_stage_2_13.Go = \adder_32bit_0.operator_B_stage_1_13.Go | _0184_;
  assign \adder_32bit_0.operator_B_stage_2_14.Po = \adder_32bit_0.operator_B_stage_1_14.Po & \adder_32bit_0.operator_B_stage_1_13.Po ;
  assign _0185_ = \adder_32bit_0.operator_B_stage_1_14.Po & \adder_32bit_0.operator_B_stage_1_13.Go ;
  assign \adder_32bit_0.operator_B_stage_2_14.Go = \adder_32bit_0.operator_B_stage_1_14.Go | _0185_;
  assign \adder_32bit_0.operator_B_stage_2_15.Po = \adder_32bit_0.operator_B_stage_1_15.Po & \adder_32bit_0.operator_B_stage_1_14.Po ;
  assign _0186_ = \adder_32bit_0.operator_B_stage_1_15.Po & \adder_32bit_0.operator_B_stage_1_14.Go ;
  assign \adder_32bit_0.operator_B_stage_2_15.Go = \adder_32bit_0.operator_B_stage_1_15.Go | _0186_;
  assign \adder_32bit_0.operator_B_stage_2_2.Po = \adder_32bit_0.operator_B_stage_1_2.Po & \adder_32bit_0.operator_B_stage_1_1.Po ;
  assign _0187_ = \adder_32bit_0.operator_B_stage_1_2.Po & \adder_32bit_0.operator_B_stage_1_1.Go ;
  assign \adder_32bit_0.operator_B_stage_2_2.Go = \adder_32bit_0.operator_B_stage_1_2.Go | _0187_;
  assign \adder_32bit_0.operator_B_stage_2_3.Po = \adder_32bit_0.operator_B_stage_1_3.Po & \adder_32bit_0.operator_B_stage_1_2.Po ;
  assign _0188_ = \adder_32bit_0.operator_B_stage_1_3.Po & \adder_32bit_0.operator_B_stage_1_2.Go ;
  assign \adder_32bit_0.operator_B_stage_2_3.Go = \adder_32bit_0.operator_B_stage_1_3.Go | _0188_;
  assign \adder_32bit_0.operator_B_stage_2_4.Po = \adder_32bit_0.operator_B_stage_1_4.Po & \adder_32bit_0.operator_B_stage_1_3.Po ;
  assign _0189_ = \adder_32bit_0.operator_B_stage_1_4.Po & \adder_32bit_0.operator_B_stage_1_3.Go ;
  assign \adder_32bit_0.operator_B_stage_2_4.Go = \adder_32bit_0.operator_B_stage_1_4.Go | _0189_;
  assign \adder_32bit_0.operator_B_stage_2_5.Po = \adder_32bit_0.operator_B_stage_1_5.Po & \adder_32bit_0.operator_B_stage_1_4.Po ;
  assign _0190_ = \adder_32bit_0.operator_B_stage_1_5.Po & \adder_32bit_0.operator_B_stage_1_4.Go ;
  assign \adder_32bit_0.operator_B_stage_2_5.Go = \adder_32bit_0.operator_B_stage_1_5.Go | _0190_;
  assign \adder_32bit_0.operator_B_stage_2_6.Po = \adder_32bit_0.operator_B_stage_1_6.Po & \adder_32bit_0.operator_B_stage_1_5.Po ;
  assign _0191_ = \adder_32bit_0.operator_B_stage_1_6.Po & \adder_32bit_0.operator_B_stage_1_5.Go ;
  assign \adder_32bit_0.operator_B_stage_2_6.Go = \adder_32bit_0.operator_B_stage_1_6.Go | _0191_;
  assign \adder_32bit_0.operator_B_stage_2_7.Po = \adder_32bit_0.operator_B_stage_1_7.Po & \adder_32bit_0.operator_B_stage_1_6.Po ;
  assign _0192_ = \adder_32bit_0.operator_B_stage_1_7.Po & \adder_32bit_0.operator_B_stage_1_6.Go ;
  assign \adder_32bit_0.operator_B_stage_2_7.Go = \adder_32bit_0.operator_B_stage_1_7.Go | _0192_;
  assign \adder_32bit_0.operator_B_stage_2_8.Po = \adder_32bit_0.operator_B_stage_1_8.Po & \adder_32bit_0.operator_B_stage_1_7.Po ;
  assign _0193_ = \adder_32bit_0.operator_B_stage_1_8.Po & \adder_32bit_0.operator_B_stage_1_7.Go ;
  assign \adder_32bit_0.operator_B_stage_2_8.Go = \adder_32bit_0.operator_B_stage_1_8.Go | _0193_;
  assign \adder_32bit_0.operator_B_stage_2_9.Po = \adder_32bit_0.operator_B_stage_1_9.Po & \adder_32bit_0.operator_B_stage_1_8.Po ;
  assign _0194_ = \adder_32bit_0.operator_B_stage_1_9.Po & \adder_32bit_0.operator_B_stage_1_8.Go ;
  assign \adder_32bit_0.operator_B_stage_2_9.Go = \adder_32bit_0.operator_B_stage_1_9.Go | _0194_;
  assign \adder_32bit_0.operator_B_stage_3_10.Po = \adder_32bit_0.operator_B_stage_2_10.Po & \adder_32bit_0.operator_B_stage_2_8.Po ;
  assign _0195_ = \adder_32bit_0.operator_B_stage_2_10.Po & \adder_32bit_0.operator_B_stage_2_8.Go ;
  assign \adder_32bit_0.operator_B_stage_3_10.Go = \adder_32bit_0.operator_B_stage_2_10.Go | _0195_;
  assign \adder_32bit_0.operator_B_stage_3_11.Po = \adder_32bit_0.operator_B_stage_2_11.Po & \adder_32bit_0.operator_B_stage_2_9.Po ;
  assign _0196_ = \adder_32bit_0.operator_B_stage_2_11.Po & \adder_32bit_0.operator_B_stage_2_9.Go ;
  assign \adder_32bit_0.operator_B_stage_3_11.Go = \adder_32bit_0.operator_B_stage_2_11.Go | _0196_;
  assign \adder_32bit_0.operator_B_stage_3_12.Po = \adder_32bit_0.operator_B_stage_2_12.Po & \adder_32bit_0.operator_B_stage_2_10.Po ;
  assign _0197_ = \adder_32bit_0.operator_B_stage_2_12.Po & \adder_32bit_0.operator_B_stage_2_10.Go ;
  assign \adder_32bit_0.operator_B_stage_3_12.Go = \adder_32bit_0.operator_B_stage_2_12.Go | _0197_;
  assign \adder_32bit_0.operator_B_stage_3_13.Po = \adder_32bit_0.operator_B_stage_2_13.Po & \adder_32bit_0.operator_B_stage_2_11.Po ;
  assign _0198_ = \adder_32bit_0.operator_B_stage_2_13.Po & \adder_32bit_0.operator_B_stage_2_11.Go ;
  assign \adder_32bit_0.operator_B_stage_3_13.Go = \adder_32bit_0.operator_B_stage_2_13.Go | _0198_;
  assign \adder_32bit_0.operator_B_stage_3_14.Po = \adder_32bit_0.operator_B_stage_2_14.Po & \adder_32bit_0.operator_B_stage_2_12.Po ;
  assign _0199_ = \adder_32bit_0.operator_B_stage_2_14.Po & \adder_32bit_0.operator_B_stage_2_12.Go ;
  assign \adder_32bit_0.operator_B_stage_3_14.Go = \adder_32bit_0.operator_B_stage_2_14.Go | _0199_;
  assign \adder_32bit_0.operator_B_stage_3_15.Po = \adder_32bit_0.operator_B_stage_2_15.Po & \adder_32bit_0.operator_B_stage_2_13.Po ;
  assign _0200_ = \adder_32bit_0.operator_B_stage_2_15.Po & \adder_32bit_0.operator_B_stage_2_13.Go ;
  assign \adder_32bit_0.operator_B_stage_3_15.Go = \adder_32bit_0.operator_B_stage_2_15.Go | _0200_;
  assign \adder_32bit_0.operator_B_stage_3_4.Po = \adder_32bit_0.operator_B_stage_2_4.Po & \adder_32bit_0.operator_B_stage_2_2.Po ;
  assign _0201_ = \adder_32bit_0.operator_B_stage_2_4.Po & \adder_32bit_0.operator_B_stage_2_2.Go ;
  assign \adder_32bit_0.operator_B_stage_3_4.Go = \adder_32bit_0.operator_B_stage_2_4.Go | _0201_;
  assign \adder_32bit_0.operator_B_stage_3_5.Po = \adder_32bit_0.operator_B_stage_2_5.Po & \adder_32bit_0.operator_B_stage_2_3.Po ;
  assign _0202_ = \adder_32bit_0.operator_B_stage_2_5.Po & \adder_32bit_0.operator_B_stage_2_3.Go ;
  assign \adder_32bit_0.operator_B_stage_3_5.Go = \adder_32bit_0.operator_B_stage_2_5.Go | _0202_;
  assign \adder_32bit_0.operator_B_stage_3_6.Po = \adder_32bit_0.operator_B_stage_2_6.Po & \adder_32bit_0.operator_B_stage_2_4.Po ;
  assign _0203_ = \adder_32bit_0.operator_B_stage_2_6.Po & \adder_32bit_0.operator_B_stage_2_4.Go ;
  assign \adder_32bit_0.operator_B_stage_3_6.Go = \adder_32bit_0.operator_B_stage_2_6.Go | _0203_;
  assign \adder_32bit_0.operator_B_stage_3_7.Po = \adder_32bit_0.operator_B_stage_2_7.Po & \adder_32bit_0.operator_B_stage_2_5.Po ;
  assign _0204_ = \adder_32bit_0.operator_B_stage_2_7.Po & \adder_32bit_0.operator_B_stage_2_5.Go ;
  assign \adder_32bit_0.operator_B_stage_3_7.Go = \adder_32bit_0.operator_B_stage_2_7.Go | _0204_;
  assign \adder_32bit_0.operator_B_stage_3_8.Po = \adder_32bit_0.operator_B_stage_2_8.Po & \adder_32bit_0.operator_B_stage_2_6.Po ;
  assign _0205_ = \adder_32bit_0.operator_B_stage_2_8.Po & \adder_32bit_0.operator_B_stage_2_6.Go ;
  assign \adder_32bit_0.operator_B_stage_3_8.Go = \adder_32bit_0.operator_B_stage_2_8.Go | _0205_;
  assign \adder_32bit_0.operator_B_stage_3_9.Po = \adder_32bit_0.operator_B_stage_2_9.Po & \adder_32bit_0.operator_B_stage_2_7.Po ;
  assign _0206_ = \adder_32bit_0.operator_B_stage_2_9.Po & \adder_32bit_0.operator_B_stage_2_7.Go ;
  assign \adder_32bit_0.operator_B_stage_3_9.Go = \adder_32bit_0.operator_B_stage_2_9.Go | _0206_;
  assign \adder_32bit_0.operator_B_stage_4_10.Po = \adder_32bit_0.operator_B_stage_3_10.Po & \adder_32bit_0.operator_B_stage_3_6.Po ;
  assign _0207_ = \adder_32bit_0.operator_B_stage_3_10.Po & \adder_32bit_0.operator_B_stage_3_6.Go ;
  assign \adder_32bit_0.operator_B_stage_4_10.Go = \adder_32bit_0.operator_B_stage_3_10.Go | _0207_;
  assign \adder_32bit_0.operator_B_stage_4_11.Po = \adder_32bit_0.operator_B_stage_3_11.Po & \adder_32bit_0.operator_B_stage_3_7.Po ;
  assign _0208_ = \adder_32bit_0.operator_B_stage_3_11.Po & \adder_32bit_0.operator_B_stage_3_7.Go ;
  assign \adder_32bit_0.operator_B_stage_4_11.Go = \adder_32bit_0.operator_B_stage_3_11.Go | _0208_;
  assign \adder_32bit_0.operator_B_stage_4_12.Po = \adder_32bit_0.operator_B_stage_3_12.Po & \adder_32bit_0.operator_B_stage_3_8.Po ;
  assign _0209_ = \adder_32bit_0.operator_B_stage_3_12.Po & \adder_32bit_0.operator_B_stage_3_8.Go ;
  assign \adder_32bit_0.operator_B_stage_4_12.Go = \adder_32bit_0.operator_B_stage_3_12.Go | _0209_;
  assign \adder_32bit_0.operator_B_stage_4_13.Po = \adder_32bit_0.operator_B_stage_3_13.Po & \adder_32bit_0.operator_B_stage_3_9.Po ;
  assign _0210_ = \adder_32bit_0.operator_B_stage_3_13.Po & \adder_32bit_0.operator_B_stage_3_9.Go ;
  assign \adder_32bit_0.operator_B_stage_4_13.Go = \adder_32bit_0.operator_B_stage_3_13.Go | _0210_;
  assign \adder_32bit_0.operator_B_stage_4_14.Po = \adder_32bit_0.operator_B_stage_3_14.Po & \adder_32bit_0.operator_B_stage_3_10.Po ;
  assign _0211_ = \adder_32bit_0.operator_B_stage_3_14.Po & \adder_32bit_0.operator_B_stage_3_10.Go ;
  assign \adder_32bit_0.operator_B_stage_4_14.Go = \adder_32bit_0.operator_B_stage_3_14.Go | _0211_;
  assign \adder_32bit_0.operator_B_stage_4_15.Po = \adder_32bit_0.operator_B_stage_3_15.Po & \adder_32bit_0.operator_B_stage_3_11.Po ;
  assign _0212_ = \adder_32bit_0.operator_B_stage_3_15.Po & \adder_32bit_0.operator_B_stage_3_11.Go ;
  assign \adder_32bit_0.operator_B_stage_4_15.Go = \adder_32bit_0.operator_B_stage_3_15.Go | _0212_;
  assign \adder_32bit_0.operator_B_stage_4_8.Po = \adder_32bit_0.operator_B_stage_3_8.Po & \adder_32bit_0.operator_B_stage_3_4.Po ;
  assign _0213_ = \adder_32bit_0.operator_B_stage_3_8.Po & \adder_32bit_0.operator_B_stage_3_4.Go ;
  assign \adder_32bit_0.operator_B_stage_4_8.Go = \adder_32bit_0.operator_B_stage_3_8.Go | _0213_;
  assign \adder_32bit_0.operator_B_stage_4_9.Po = \adder_32bit_0.operator_B_stage_3_9.Po & \adder_32bit_0.operator_B_stage_3_5.Po ;
  assign _0214_ = \adder_32bit_0.operator_B_stage_3_9.Po & \adder_32bit_0.operator_B_stage_3_5.Go ;
  assign \adder_32bit_0.operator_B_stage_4_9.Go = \adder_32bit_0.operator_B_stage_3_9.Go | _0214_;
  assign _0215_ = \adder_32bit_0.operator_A_0.P & cout;
  assign \adder_32bit_0.operator_C_stage_1_0.Go = \adder_32bit_0.operator_A_0.G | _0215_;
  assign _0216_ = \adder_32bit_0.operator_B_stage_1_1.Po & \adder_32bit_0.operator_C_stage_1_0.Go ;
  assign \adder_32bit_0.operator_C_stage_2_1.Go = \adder_32bit_0.operator_B_stage_1_1.Go | _0216_;
  assign _0217_ = \adder_32bit_0.operator_B_stage_2_2.Po & \adder_32bit_0.operator_C_stage_1_0.Go ;
  assign \adder_32bit_0.operator_C_stage_3_2.Go = \adder_32bit_0.operator_B_stage_2_2.Go | _0217_;
  assign _0218_ = \adder_32bit_0.operator_B_stage_2_3.Po & \adder_32bit_0.operator_C_stage_2_1.Go ;
  assign \adder_32bit_0.operator_C_stage_3_3.Go = \adder_32bit_0.operator_B_stage_2_3.Go | _0218_;
  assign _0219_ = \adder_32bit_0.operator_B_stage_3_4.Po & \adder_32bit_0.operator_C_stage_1_0.Go ;
  assign \adder_32bit_0.operator_C_stage_4_4.Go = \adder_32bit_0.operator_B_stage_3_4.Go | _0219_;
  assign _0220_ = \adder_32bit_0.operator_B_stage_3_5.Po & \adder_32bit_0.operator_C_stage_2_1.Go ;
  assign \adder_32bit_0.operator_C_stage_4_5.Go = \adder_32bit_0.operator_B_stage_3_5.Go | _0220_;
  assign _0221_ = \adder_32bit_0.operator_B_stage_3_6.Po & \adder_32bit_0.operator_C_stage_3_2.Go ;
  assign \adder_32bit_0.operator_C_stage_4_6.Go = \adder_32bit_0.operator_B_stage_3_6.Go | _0221_;
  assign _0222_ = \adder_32bit_0.operator_B_stage_3_7.Po & \adder_32bit_0.operator_C_stage_3_3.Go ;
  assign \adder_32bit_0.operator_C_stage_4_7.Go = \adder_32bit_0.operator_B_stage_3_7.Go | _0222_;
  assign _0223_ = \adder_32bit_0.operator_B_stage_4_10.Po & \adder_32bit_0.operator_C_stage_3_2.Go ;
  assign \adder_32bit_0.operator_C_stage_5_10.Go = \adder_32bit_0.operator_B_stage_4_10.Go | _0223_;
  assign _0224_ = \adder_32bit_0.operator_B_stage_4_11.Po & \adder_32bit_0.operator_C_stage_3_3.Go ;
  assign \adder_32bit_0.operator_C_stage_5_11.Go = \adder_32bit_0.operator_B_stage_4_11.Go | _0224_;
  assign _0225_ = \adder_32bit_0.operator_B_stage_4_12.Po & \adder_32bit_0.operator_C_stage_4_4.Go ;
  assign \adder_32bit_0.operator_C_stage_5_12.Go = \adder_32bit_0.operator_B_stage_4_12.Go | _0225_;
  assign _0226_ = \adder_32bit_0.operator_B_stage_4_13.Po & \adder_32bit_0.operator_C_stage_4_5.Go ;
  assign \adder_32bit_0.operator_C_stage_5_13.Go = \adder_32bit_0.operator_B_stage_4_13.Go | _0226_;
  assign _0227_ = \adder_32bit_0.operator_B_stage_4_14.Po & \adder_32bit_0.operator_C_stage_4_6.Go ;
  assign \adder_32bit_0.operator_C_stage_5_14.Go = \adder_32bit_0.operator_B_stage_4_14.Go | _0227_;
  assign _0228_ = \adder_32bit_0.operator_B_stage_4_15.Po & \adder_32bit_0.operator_C_stage_4_7.Go ;
  assign \adder_32bit_0.operator_C_stage_5_15.Go = \adder_32bit_0.operator_B_stage_4_15.Go | _0228_;
  assign _0229_ = \adder_32bit_0.operator_B_stage_4_8.Po & \adder_32bit_0.operator_C_stage_1_0.Go ;
  assign \adder_32bit_0.operator_C_stage_5_8.Go = \adder_32bit_0.operator_B_stage_4_8.Go | _0229_;
  assign _0230_ = \adder_32bit_0.operator_B_stage_4_9.Po & \adder_32bit_0.operator_C_stage_2_1.Go ;
  assign \adder_32bit_0.operator_C_stage_5_9.Go = \adder_32bit_0.operator_B_stage_4_9.Go | _0230_;
  assign _0231_ = \adder_32bit_0.operator_A_1.P & \adder_32bit_0.operator_C_stage_1_0.Go ;
  assign \adder_32bit_0.operator_C_stage_6_0.Go = \adder_32bit_0.operator_A_1.G | _0231_;
  assign _0232_ = \adder_32bit_0.operator_A_3.P & \adder_32bit_0.operator_C_stage_2_1.Go ;
  assign \adder_32bit_0.operator_C_stage_6_1.Go = \adder_32bit_0.operator_A_3.G | _0232_;
  assign _0233_ = \adder_32bit_0.operator_A_21.P & \adder_32bit_0.operator_C_stage_5_10.Go ;
  assign \adder_32bit_0.operator_C_stage_6_10.Go = \adder_32bit_0.operator_A_21.G | _0233_;
  assign _0234_ = \adder_32bit_0.operator_A_23.P & \adder_32bit_0.operator_C_stage_5_11.Go ;
  assign \adder_32bit_0.operator_C_stage_6_11.Go = \adder_32bit_0.operator_A_23.G | _0234_;
  assign _0235_ = \adder_32bit_0.operator_A_25.P & \adder_32bit_0.operator_C_stage_5_12.Go ;
  assign \adder_32bit_0.operator_C_stage_6_12.Go = \adder_32bit_0.operator_A_25.G | _0235_;
  assign _0236_ = \adder_32bit_0.operator_A_27.P & \adder_32bit_0.operator_C_stage_5_13.Go ;
  assign \adder_32bit_0.operator_C_stage_6_13.Go = \adder_32bit_0.operator_A_27.G | _0236_;
  assign _0237_ = \adder_32bit_0.operator_A_29.P & \adder_32bit_0.operator_C_stage_5_14.Go ;
  assign \adder_32bit_0.operator_C_stage_6_14.Go = \adder_32bit_0.operator_A_29.G | _0237_;
  assign _0238_ = \adder_32bit_0.operator_A_5.P & \adder_32bit_0.operator_C_stage_3_2.Go ;
  assign \adder_32bit_0.operator_C_stage_6_2.Go = \adder_32bit_0.operator_A_5.G | _0238_;
  assign _0239_ = \adder_32bit_0.operator_A_7.P & \adder_32bit_0.operator_C_stage_3_3.Go ;
  assign \adder_32bit_0.operator_C_stage_6_3.Go = \adder_32bit_0.operator_A_7.G | _0239_;
  assign _0240_ = \adder_32bit_0.operator_A_9.P & \adder_32bit_0.operator_C_stage_4_4.Go ;
  assign \adder_32bit_0.operator_C_stage_6_4.Go = \adder_32bit_0.operator_A_9.G | _0240_;
  assign _0241_ = \adder_32bit_0.operator_A_11.P & \adder_32bit_0.operator_C_stage_4_5.Go ;
  assign \adder_32bit_0.operator_C_stage_6_5.Go = \adder_32bit_0.operator_A_11.G | _0241_;
  assign _0242_ = \adder_32bit_0.operator_A_13.P & \adder_32bit_0.operator_C_stage_4_6.Go ;
  assign \adder_32bit_0.operator_C_stage_6_6.Go = \adder_32bit_0.operator_A_13.G | _0242_;
  assign _0243_ = \adder_32bit_0.operator_A_15.P & \adder_32bit_0.operator_C_stage_4_7.Go ;
  assign \adder_32bit_0.operator_C_stage_6_7.Go = \adder_32bit_0.operator_A_15.G | _0243_;
  assign _0244_ = \adder_32bit_0.operator_A_17.P & \adder_32bit_0.operator_C_stage_5_8.Go ;
  assign \adder_32bit_0.operator_C_stage_6_8.Go = \adder_32bit_0.operator_A_17.G | _0244_;
  assign _0245_ = \adder_32bit_0.operator_A_19.P & \adder_32bit_0.operator_C_stage_5_9.Go ;
  assign \adder_32bit_0.operator_C_stage_6_9.Go = \adder_32bit_0.operator_A_19.G | _0245_;
  always @(posedge i_clk)
    if (!\multiplier_16x16bit_pipelined.i_rst )
      \multiplier_16x16bit_pipelined.reg_layer_2_w0 <= 2'b00;
    else
      \multiplier_16x16bit_pipelined.reg_layer_2_w0 <= _0248_;
  always @(posedge i_clk)
    if (!\multiplier_16x16bit_pipelined.i_rst )
      \multiplier_16x16bit_pipelined.reg_layer_2_w1 <= 1'b0;
    else
      \multiplier_16x16bit_pipelined.reg_layer_2_w1 <= _0259_;
  always @(posedge i_clk)
    if (!\multiplier_16x16bit_pipelined.i_rst )
      \multiplier_16x16bit_pipelined.reg_layer_2_w2 <= 3'b000;
    else
      \multiplier_16x16bit_pipelined.reg_layer_2_w2 <= _0270_;
  always @(posedge i_clk)
    if (!\multiplier_16x16bit_pipelined.i_rst )
      \multiplier_16x16bit_pipelined.reg_layer_2_w3 <= 2'b00;
    else
      \multiplier_16x16bit_pipelined.reg_layer_2_w3 <= _0273_;
  always @(posedge i_clk)
    if (!\multiplier_16x16bit_pipelined.i_rst )
      \multiplier_16x16bit_pipelined.reg_layer_2_w4 <= 2'b00;
    else
      \multiplier_16x16bit_pipelined.reg_layer_2_w4 <= _0274_;
  always @(posedge i_clk)
    if (!\multiplier_16x16bit_pipelined.i_rst )
      \multiplier_16x16bit_pipelined.reg_layer_2_w5 <= 2'b00;
    else
      \multiplier_16x16bit_pipelined.reg_layer_2_w5 <= _0275_;
  always @(posedge i_clk)
    if (!\multiplier_16x16bit_pipelined.i_rst )
      \multiplier_16x16bit_pipelined.reg_layer_2_w6 <= 2'b00;
    else
      \multiplier_16x16bit_pipelined.reg_layer_2_w6 <= _0276_;
  always @(posedge i_clk)
    if (!\multiplier_16x16bit_pipelined.i_rst )
      \multiplier_16x16bit_pipelined.reg_layer_2_w7 <= 2'b00;
    else
      \multiplier_16x16bit_pipelined.reg_layer_2_w7 <= _0277_;
  always @(posedge i_clk)
    if (!\multiplier_16x16bit_pipelined.i_rst )
      \multiplier_16x16bit_pipelined.reg_layer_2_w8 <= 2'b00;
    else
      \multiplier_16x16bit_pipelined.reg_layer_2_w8 <= _0278_;
  always @(posedge i_clk)
    if (!\multiplier_16x16bit_pipelined.i_rst )
      \multiplier_16x16bit_pipelined.reg_layer_2_w9 <= 2'b00;
    else
      \multiplier_16x16bit_pipelined.reg_layer_2_w9 <= _0279_;
  always @(posedge i_clk)
    if (!\multiplier_16x16bit_pipelined.i_rst )
      \multiplier_16x16bit_pipelined.reg_layer_2_w10 <= 2'b00;
    else
      \multiplier_16x16bit_pipelined.reg_layer_2_w10 <= _0249_;
  always @(posedge i_clk)
    if (!\multiplier_16x16bit_pipelined.i_rst )
      \multiplier_16x16bit_pipelined.reg_layer_2_w11 <= 4'b0000;
    else
      \multiplier_16x16bit_pipelined.reg_layer_2_w11 <= _0250_;
  always @(posedge i_clk)
    if (!\multiplier_16x16bit_pipelined.i_rst )
      \multiplier_16x16bit_pipelined.reg_layer_2_w12 <= 3'b000;
    else
      \multiplier_16x16bit_pipelined.reg_layer_2_w12 <= _0251_;
  always @(posedge i_clk)
    if (!\multiplier_16x16bit_pipelined.i_rst )
      \multiplier_16x16bit_pipelined.reg_layer_2_w13 <= 3'b000;
    else
      \multiplier_16x16bit_pipelined.reg_layer_2_w13 <= _0252_;
  always @(posedge i_clk)
    if (!\multiplier_16x16bit_pipelined.i_rst )
      \multiplier_16x16bit_pipelined.reg_layer_2_w14 <= 3'b000;
    else
      \multiplier_16x16bit_pipelined.reg_layer_2_w14 <= _0253_;
  always @(posedge i_clk)
    if (!\multiplier_16x16bit_pipelined.i_rst )
      \multiplier_16x16bit_pipelined.reg_layer_2_w15 <= 3'b000;
    else
      \multiplier_16x16bit_pipelined.reg_layer_2_w15 <= _0254_;
  always @(posedge i_clk)
    if (!\multiplier_16x16bit_pipelined.i_rst )
      \multiplier_16x16bit_pipelined.reg_layer_2_w16 <= 4'b0000;
    else
      \multiplier_16x16bit_pipelined.reg_layer_2_w16 <= _0255_;
  always @(posedge i_clk)
    if (!\multiplier_16x16bit_pipelined.i_rst )
      \multiplier_16x16bit_pipelined.reg_layer_2_w17 <= 3'b000;
    else
      \multiplier_16x16bit_pipelined.reg_layer_2_w17 <= _0256_;
  always @(posedge i_clk)
    if (!\multiplier_16x16bit_pipelined.i_rst )
      \multiplier_16x16bit_pipelined.reg_layer_2_w18 <= 4'b0000;
    else
      \multiplier_16x16bit_pipelined.reg_layer_2_w18 <= _0257_;
  always @(posedge i_clk)
    if (!\multiplier_16x16bit_pipelined.i_rst )
      \multiplier_16x16bit_pipelined.reg_layer_2_w19 <= 3'b000;
    else
      \multiplier_16x16bit_pipelined.reg_layer_2_w19 <= _0258_;
  always @(posedge i_clk)
    if (!\multiplier_16x16bit_pipelined.i_rst )
      \multiplier_16x16bit_pipelined.reg_layer_2_w20 <= 4'b0000;
    else
      \multiplier_16x16bit_pipelined.reg_layer_2_w20 <= _0260_;
  always @(posedge i_clk)
    if (!\multiplier_16x16bit_pipelined.i_rst )
      \multiplier_16x16bit_pipelined.reg_layer_2_w21 <= 3'b000;
    else
      \multiplier_16x16bit_pipelined.reg_layer_2_w21 <= _0261_;
  always @(posedge i_clk)
    if (!\multiplier_16x16bit_pipelined.i_rst )
      \multiplier_16x16bit_pipelined.reg_layer_2_w22 <= 2'b00;
    else
      \multiplier_16x16bit_pipelined.reg_layer_2_w22 <= _0262_;
  always @(posedge i_clk)
    if (!\multiplier_16x16bit_pipelined.i_rst )
      \multiplier_16x16bit_pipelined.reg_layer_2_w23 <= 2'b00;
    else
      \multiplier_16x16bit_pipelined.reg_layer_2_w23 <= _0263_;
  always @(posedge i_clk)
    if (!\multiplier_16x16bit_pipelined.i_rst )
      \multiplier_16x16bit_pipelined.reg_layer_2_w24 <= 3'b000;
    else
      \multiplier_16x16bit_pipelined.reg_layer_2_w24 <= _0264_;
  always @(posedge i_clk)
    if (!\multiplier_16x16bit_pipelined.i_rst )
      \multiplier_16x16bit_pipelined.reg_layer_2_w25 <= 2'b00;
    else
      \multiplier_16x16bit_pipelined.reg_layer_2_w25 <= _0265_;
  always @(posedge i_clk)
    if (!\multiplier_16x16bit_pipelined.i_rst )
      \multiplier_16x16bit_pipelined.reg_layer_2_w26 <= 3'b000;
    else
      \multiplier_16x16bit_pipelined.reg_layer_2_w26 <= _0266_;
  always @(posedge i_clk)
    if (!\multiplier_16x16bit_pipelined.i_rst )
      \multiplier_16x16bit_pipelined.reg_layer_2_w27 <= 2'b00;
    else
      \multiplier_16x16bit_pipelined.reg_layer_2_w27 <= _0267_;
  always @(posedge i_clk)
    if (!\multiplier_16x16bit_pipelined.i_rst )
      \multiplier_16x16bit_pipelined.reg_layer_2_w28 <= 1'b0;
    else
      \multiplier_16x16bit_pipelined.reg_layer_2_w28 <= _0268_;
  always @(posedge i_clk)
    if (!\multiplier_16x16bit_pipelined.i_rst )
      \multiplier_16x16bit_pipelined.reg_layer_2_w29 <= 3'b000;
    else
      \multiplier_16x16bit_pipelined.reg_layer_2_w29 <= _0269_;
  always @(posedge i_clk)
    if (!\multiplier_16x16bit_pipelined.i_rst )
      \multiplier_16x16bit_pipelined.reg_layer_2_w30 <= 1'b0;
    else
      \multiplier_16x16bit_pipelined.reg_layer_2_w30 <= _0271_;
  always @(posedge i_clk)
    if (!\multiplier_16x16bit_pipelined.i_rst )
      \multiplier_16x16bit_pipelined.reg_layer_2_w31 <= 1'b0;
    else
      \multiplier_16x16bit_pipelined.reg_layer_2_w31 <= _0272_;
  always @(posedge i_clk)
    if (!\multiplier_16x16bit_pipelined.i_rst )
      \multiplier_16x16bit_pipelined.md <= 16'b0000000000000000;
    else
      \multiplier_16x16bit_pipelined.md <= _0246_;
  always @(posedge i_clk)
    if (!\multiplier_16x16bit_pipelined.i_rst )
      \multiplier_16x16bit_pipelined.mr <= 16'b0000000000000000;
    else
      \multiplier_16x16bit_pipelined.mr <= _0247_;
  always @(posedge i_clk)
    if (!\multiplier_16x16bit_pipelined.i_rst )
      \multiplier_16x16bit_pipelined.stage_0_ready <= 1'b0;
    else
      \multiplier_16x16bit_pipelined.stage_0_ready <= start;
  assign _0272_ = \multiplier_16x16bit_pipelined.stage_0_ready ? 1'b1 : \multiplier_16x16bit_pipelined.reg_layer_2_w31 ;
  assign _0271_ = \multiplier_16x16bit_pipelined.stage_0_ready ? \multiplier_16x16bit_pipelined.layer_0_w30 : \multiplier_16x16bit_pipelined.reg_layer_2_w30 ;
  wire [2:0] fangyuan46;
  assign fangyuan46 = { 1'b1, \multiplier_16x16bit_pipelined.layer_0_w29[0] , \multiplier_16x16bit_pipelined.layer_2_full_adder_11.cout };

  assign _0269_ = \multiplier_16x16bit_pipelined.stage_0_ready ? fangyuan46 : \multiplier_16x16bit_pipelined.reg_layer_2_w29 ;
  assign _0268_ = \multiplier_16x16bit_pipelined.stage_0_ready ? \multiplier_16x16bit_pipelined.layer_2_full_adder_11.S : \multiplier_16x16bit_pipelined.reg_layer_2_w28 ;
  wire [1:0] fangyuan47;
  assign fangyuan47 = { \multiplier_16x16bit_pipelined.layer_1_full_adder_11.S , \multiplier_16x16bit_pipelined.layer_1_full_adder_10.cout };

  assign _0267_ = \multiplier_16x16bit_pipelined.stage_0_ready ? fangyuan47 : \multiplier_16x16bit_pipelined.reg_layer_2_w27 ;
  wire [2:0] fangyuan48;
  assign fangyuan48 = { \multiplier_16x16bit_pipelined.layer_1_full_adder_10.S , \multiplier_16x16bit_pipelined.layer_1_full_adder_9.cout , \multiplier_16x16bit_pipelined.layer_2_full_adder_10.cout };

  assign _0266_ = \multiplier_16x16bit_pipelined.stage_0_ready ? fangyuan48 : \multiplier_16x16bit_pipelined.reg_layer_2_w26 ;
  wire [1:0] fangyuan49;
  assign fangyuan49 = { \multiplier_16x16bit_pipelined.layer_2_full_adder_10.S , \multiplier_16x16bit_pipelined.layer_2_full_adder_9.cout };

  assign _0265_ = \multiplier_16x16bit_pipelined.stage_0_ready ? fangyuan49 : \multiplier_16x16bit_pipelined.reg_layer_2_w25 ;
  wire [2:0] fangyuan50;
  assign fangyuan50 = { \multiplier_16x16bit_pipelined.layer_0_w24[3] , \multiplier_16x16bit_pipelined.layer_2_full_adder_9.S , \multiplier_16x16bit_pipelined.layer_2_full_adder_8.cout };

  assign _0264_ = \multiplier_16x16bit_pipelined.stage_0_ready ? fangyuan50 : \multiplier_16x16bit_pipelined.reg_layer_2_w24 ;
  wire [1:0] fangyuan51;
  assign fangyuan51 = { \multiplier_16x16bit_pipelined.layer_2_full_adder_8.S , \multiplier_16x16bit_pipelined.layer_2_full_adder_7.cout };

  assign _0263_ = \multiplier_16x16bit_pipelined.stage_0_ready ? fangyuan51 : \multiplier_16x16bit_pipelined.reg_layer_2_w23 ;
  wire [1:0] fangyuan52;
  assign fangyuan52 = { \multiplier_16x16bit_pipelined.layer_2_full_adder_7.S , \multiplier_16x16bit_pipelined.layer_2_full_adder_6.cout };

  assign _0262_ = \multiplier_16x16bit_pipelined.stage_0_ready ? fangyuan52 : \multiplier_16x16bit_pipelined.reg_layer_2_w22 ;
  wire [2:0] fangyuan53;
  assign fangyuan53 = { 1'b1, \multiplier_16x16bit_pipelined.layer_2_full_adder_6.S , \multiplier_16x16bit_pipelined.layer_2_full_adder_5.cout };

  assign _0261_ = \multiplier_16x16bit_pipelined.stage_0_ready ? fangyuan53 : \multiplier_16x16bit_pipelined.reg_layer_2_w21 ;
  wire [3:0] fangyuan54;
  assign fangyuan54 = { \multiplier_16x16bit_pipelined.layer_0_w20[5] , \multiplier_16x16bit_pipelined.layer_2_full_adder_5.S , \multiplier_16x16bit_pipelined.layer_2_compressor42_7.cout , \multiplier_16x16bit_pipelined.layer_2_compressor42_7.carry };

  assign _0260_ = \multiplier_16x16bit_pipelined.stage_0_ready ? fangyuan54 : \multiplier_16x16bit_pipelined.reg_layer_2_w20 ;
  wire [2:0] fangyuan55;
  assign fangyuan55 = { \multiplier_16x16bit_pipelined.layer_2_compressor42_7.S , \multiplier_16x16bit_pipelined.layer_2_compressor42_6.cout , \multiplier_16x16bit_pipelined.layer_2_compressor42_6.carry };

  assign _0258_ = \multiplier_16x16bit_pipelined.stage_0_ready ? fangyuan55 : \multiplier_16x16bit_pipelined.reg_layer_2_w19 ;
  wire [3:0] fangyuan56;
  assign fangyuan56 = { \multiplier_16x16bit_pipelined.layer_0_w18[6] , \multiplier_16x16bit_pipelined.layer_2_compressor42_6.S , \multiplier_16x16bit_pipelined.layer_2_compressor42_5.cout , \multiplier_16x16bit_pipelined.layer_2_compressor42_5.carry };

  assign _0257_ = \multiplier_16x16bit_pipelined.stage_0_ready ? fangyuan56 : \multiplier_16x16bit_pipelined.reg_layer_2_w18 ;
  wire [2:0] fangyuan57;
  assign fangyuan57 = { \multiplier_16x16bit_pipelined.layer_2_compressor42_5.S , \multiplier_16x16bit_pipelined.layer_2_compressor42_4.cout , \multiplier_16x16bit_pipelined.layer_2_compressor42_4.carry };

  assign _0256_ = \multiplier_16x16bit_pipelined.stage_0_ready ? fangyuan57 : \multiplier_16x16bit_pipelined.reg_layer_2_w17 ;
  wire [3:0] fangyuan58;
  assign fangyuan58 = { 1'b1, \multiplier_16x16bit_pipelined.layer_2_compressor42_4.S , \multiplier_16x16bit_pipelined.layer_2_compressor42_3.cout , \multiplier_16x16bit_pipelined.layer_2_compressor42_3.carry };

  assign _0255_ = \multiplier_16x16bit_pipelined.stage_0_ready ? fangyuan58 : \multiplier_16x16bit_pipelined.reg_layer_2_w16 ;
  wire [2:0] fangyuan59;
  assign fangyuan59 = { \multiplier_16x16bit_pipelined.layer_2_compressor42_3.S , \multiplier_16x16bit_pipelined.layer_2_compressor42_2.cout , \multiplier_16x16bit_pipelined.layer_2_compressor42_2.carry };

  assign _0254_ = \multiplier_16x16bit_pipelined.stage_0_ready ? fangyuan59 : \multiplier_16x16bit_pipelined.reg_layer_2_w15 ;
  wire [2:0] fangyuan60;
  assign fangyuan60 = { \multiplier_16x16bit_pipelined.layer_2_compressor42_2.S , \multiplier_16x16bit_pipelined.layer_2_compressor42_1.cout , \multiplier_16x16bit_pipelined.layer_2_compressor42_1.carry };

  assign _0253_ = \multiplier_16x16bit_pipelined.stage_0_ready ? fangyuan60 : \multiplier_16x16bit_pipelined.reg_layer_2_w14 ;
  wire [2:0] fangyuan61;
  assign fangyuan61 = { \multiplier_16x16bit_pipelined.layer_0_w13[6] , \multiplier_16x16bit_pipelined.layer_2_compressor42_1.S , \multiplier_16x16bit_pipelined.layer_2_full_adder_4.cout };

  assign _0252_ = \multiplier_16x16bit_pipelined.stage_0_ready ? fangyuan61 : \multiplier_16x16bit_pipelined.reg_layer_2_w13 ;
  wire [2:0] fangyuan62;
  assign fangyuan62 = { \multiplier_16x16bit_pipelined.layer_1_full_adder_3.S , \multiplier_16x16bit_pipelined.layer_2_full_adder_4.S , \multiplier_16x16bit_pipelined.layer_2_full_adder_3.cout };

  assign _0251_ = \multiplier_16x16bit_pipelined.stage_0_ready ? fangyuan62 : \multiplier_16x16bit_pipelined.reg_layer_2_w12 ;
  wire [3:0] fangyuan63;
  assign fangyuan63 = { \multiplier_16x16bit_pipelined.layer_0_w11[5] , \multiplier_16x16bit_pipelined.layer_2_full_adder_3.S , \multiplier_16x16bit_pipelined.layer_2_compressor42_0.cout , \multiplier_16x16bit_pipelined.layer_2_compressor42_0.carry };

  assign _0250_ = \multiplier_16x16bit_pipelined.stage_0_ready ? fangyuan63 : \multiplier_16x16bit_pipelined.reg_layer_2_w11 ;
  wire [1:0] fangyuan64;
  assign fangyuan64 = { \multiplier_16x16bit_pipelined.layer_2_compressor42_0.S , \multiplier_16x16bit_pipelined.layer_2_full_adder_2.cout };

  assign _0249_ = \multiplier_16x16bit_pipelined.stage_0_ready ? fangyuan64 : \multiplier_16x16bit_pipelined.reg_layer_2_w10 ;
  wire [1:0] fangyuan65;
  assign fangyuan65 = { \multiplier_16x16bit_pipelined.layer_2_full_adder_2.S , \multiplier_16x16bit_pipelined.layer_2_full_adder_1.cout };

  assign _0279_ = \multiplier_16x16bit_pipelined.stage_0_ready ? fangyuan65 : \multiplier_16x16bit_pipelined.reg_layer_2_w9 ;
  wire [1:0] fangyuan66;
  assign fangyuan66 = { \multiplier_16x16bit_pipelined.layer_2_full_adder_1.S , \multiplier_16x16bit_pipelined.layer_2_full_adder_0.cout };

  assign _0278_ = \multiplier_16x16bit_pipelined.stage_0_ready ? fangyuan66 : \multiplier_16x16bit_pipelined.reg_layer_2_w8 ;
  wire [1:0] fangyuan67;
  assign fangyuan67 = { \multiplier_16x16bit_pipelined.layer_0_w7[3] , \multiplier_16x16bit_pipelined.layer_2_full_adder_0.S };

  assign _0277_ = \multiplier_16x16bit_pipelined.stage_0_ready ? fangyuan67 : \multiplier_16x16bit_pipelined.reg_layer_2_w7 ;
  wire [1:0] fangyuan68;
  assign fangyuan68 = { \multiplier_16x16bit_pipelined.layer_1_compressor42_0.S , \multiplier_16x16bit_pipelined.layer_1_full_adder_1.cout };

  assign _0276_ = \multiplier_16x16bit_pipelined.stage_0_ready ? fangyuan68 : \multiplier_16x16bit_pipelined.reg_layer_2_w6 ;
  wire [1:0] fangyuan69;
  assign fangyuan69 = { \multiplier_16x16bit_pipelined.layer_1_full_adder_1.S , \multiplier_16x16bit_pipelined.layer_1_full_adder_0.cout };

  assign _0275_ = \multiplier_16x16bit_pipelined.stage_0_ready ? fangyuan69 : \multiplier_16x16bit_pipelined.reg_layer_2_w5 ;
  wire [1:0] fangyuan70;
  assign fangyuan70 = { \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_2.negation , \multiplier_16x16bit_pipelined.layer_1_full_adder_0.S };

  assign _0274_ = \multiplier_16x16bit_pipelined.stage_0_ready ? fangyuan70 : \multiplier_16x16bit_pipelined.reg_layer_2_w4 ;
  wire [1:0] fangyuan71;
  assign fangyuan71 = { \multiplier_16x16bit_pipelined.layer_0_w3[1] , \multiplier_16x16bit_pipelined.layer_0_w3[0] };

  assign _0273_ = \multiplier_16x16bit_pipelined.stage_0_ready ? fangyuan71 : \multiplier_16x16bit_pipelined.reg_layer_2_w3 ;
  wire [2:0] fangyuan72;
  assign fangyuan72 = { \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_1.negation , \multiplier_16x16bit_pipelined.layer_0_w2[1] , \multiplier_16x16bit_pipelined.layer_0_w2[0] };

  assign _0270_ = \multiplier_16x16bit_pipelined.stage_0_ready ? fangyuan72 : \multiplier_16x16bit_pipelined.reg_layer_2_w2 ;
  assign _0259_ = \multiplier_16x16bit_pipelined.stage_0_ready ? \multiplier_16x16bit_pipelined.layer_0_w1 : \multiplier_16x16bit_pipelined.reg_layer_2_w1 ;
  wire [1:0] fangyuan73;
  assign fangyuan73 = { \multiplier_16x16bit_pipelined.mr [1], \multiplier_16x16bit_pipelined.layer_0_w0[0] };

  assign _0248_ = \multiplier_16x16bit_pipelined.stage_0_ready ? fangyuan73 : \multiplier_16x16bit_pipelined.reg_layer_2_w0 ;
  assign _0247_ = start ? mr : \multiplier_16x16bit_pipelined.mr ;
  assign _0246_ = start ? md : \multiplier_16x16bit_pipelined.md ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.o_s [1] = \multiplier_16x16bit_pipelined.reg_layer_2_w1 ^ \multiplier_16x16bit_pipelined.adder_32bit.operator_A_0.G ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.o_s [2] = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_2.A ^ \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_6_0.Go ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.o_s [3] = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_3.P ^ \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_2_1.Go ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.o_s [4] = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_4.P ^ \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_6_1.Go ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.o_s [5] = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_5.P ^ \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_3_2.Go ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.o_s [6] = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_6.P ^ \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_6_2.Go ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.o_s [7] = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_7.P ^ \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_3_3.Go ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.o_s [8] = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_8.P ^ \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_6_3.Go ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.o_s [9] = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_9.P ^ \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_4_4.Go ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.o_s [10] = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_10.P ^ \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_6_4.Go ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.o_s [11] = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_11.P ^ \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_4_5.Go ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.o_s [12] = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_12.P ^ \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_6_5.Go ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.o_s [13] = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_13.P ^ \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_4_6.Go ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.o_s [14] = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_14.P ^ \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_6_6.Go ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.o_s [15] = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_15.P ^ \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_4_7.Go ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.o_s [16] = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_16.P ^ \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_6_7.Go ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.o_s [17] = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_17.P ^ \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_5_8.Go ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.o_s [18] = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_18.P ^ \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_6_8.Go ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.o_s [19] = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_19.P ^ \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_5_9.Go ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.o_s [20] = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_20.P ^ \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_6_9.Go ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.o_s [21] = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_21.P ^ \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_5_10.Go ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.o_s [22] = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_22.P ^ \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_6_10.Go ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.o_s [23] = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_23.P ^ \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_5_11.Go ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.o_s [24] = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_24.P ^ \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_6_11.Go ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.o_s [25] = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_25.A ^ \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_5_12.Go ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.o_s [26] = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_26.P ^ \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_6_12.Go ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.o_s [27] = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_27.A ^ \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_5_13.Go ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.o_s [28] = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_28.P ^ \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_6_13.Go ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.o_s [29] = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_29.A ^ \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_5_14.Go ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.o_s [30] = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_30.P ^ \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_6_14.Go ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.o_s [31] = \multiplier_16x16bit_pipelined.reg_layer_2_w31 ^ \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_5_15.Go ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_A_0.G = \multiplier_16x16bit_pipelined.reg_layer_2_w0 [0] & \multiplier_16x16bit_pipelined.reg_layer_2_w0 [1];
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_A_0.P = \multiplier_16x16bit_pipelined.reg_layer_2_w0 [0] ^ \multiplier_16x16bit_pipelined.reg_layer_2_w0 [1];
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_A_10.G = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_10.A & \multiplier_16x16bit_pipelined.adder_32bit.operator_A_10.B ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_A_10.P = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_10.A ^ \multiplier_16x16bit_pipelined.adder_32bit.operator_A_10.B ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_A_11.G = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_11.A & \multiplier_16x16bit_pipelined.adder_32bit.operator_A_11.B ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_A_11.P = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_11.A ^ \multiplier_16x16bit_pipelined.adder_32bit.operator_A_11.B ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_A_12.G = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_12.A & \multiplier_16x16bit_pipelined.adder_32bit.operator_A_12.B ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_A_12.P = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_12.A ^ \multiplier_16x16bit_pipelined.adder_32bit.operator_A_12.B ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_A_13.G = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_13.A & \multiplier_16x16bit_pipelined.adder_32bit.operator_A_13.B ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_A_13.P = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_13.A ^ \multiplier_16x16bit_pipelined.adder_32bit.operator_A_13.B ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_A_14.G = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_14.A & \multiplier_16x16bit_pipelined.adder_32bit.operator_A_14.B ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_A_14.P = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_14.A ^ \multiplier_16x16bit_pipelined.adder_32bit.operator_A_14.B ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_A_15.G = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_15.A & \multiplier_16x16bit_pipelined.adder_32bit.operator_A_15.B ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_A_15.P = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_15.A ^ \multiplier_16x16bit_pipelined.adder_32bit.operator_A_15.B ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_A_16.G = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_16.A & \multiplier_16x16bit_pipelined.adder_32bit.operator_A_16.B ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_A_16.P = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_16.A ^ \multiplier_16x16bit_pipelined.adder_32bit.operator_A_16.B ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_A_17.G = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_17.A & \multiplier_16x16bit_pipelined.adder_32bit.operator_A_17.B ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_A_17.P = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_17.A ^ \multiplier_16x16bit_pipelined.adder_32bit.operator_A_17.B ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_A_18.G = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_18.A & \multiplier_16x16bit_pipelined.adder_32bit.operator_A_18.B ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_A_18.P = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_18.A ^ \multiplier_16x16bit_pipelined.adder_32bit.operator_A_18.B ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_A_19.G = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_19.A & \multiplier_16x16bit_pipelined.adder_32bit.operator_A_19.B ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_A_19.P = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_19.A ^ \multiplier_16x16bit_pipelined.adder_32bit.operator_A_19.B ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_A_20.G = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_20.A & \multiplier_16x16bit_pipelined.adder_32bit.operator_A_20.B ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_A_20.P = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_20.A ^ \multiplier_16x16bit_pipelined.adder_32bit.operator_A_20.B ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_A_21.G = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_21.A & \multiplier_16x16bit_pipelined.adder_32bit.operator_A_21.B ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_A_21.P = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_21.A ^ \multiplier_16x16bit_pipelined.adder_32bit.operator_A_21.B ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_A_22.G = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_22.A & \multiplier_16x16bit_pipelined.adder_32bit.operator_A_22.B ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_A_22.P = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_22.A ^ \multiplier_16x16bit_pipelined.adder_32bit.operator_A_22.B ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_A_23.G = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_23.A & \multiplier_16x16bit_pipelined.adder_32bit.operator_A_23.B ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_A_23.P = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_23.A ^ \multiplier_16x16bit_pipelined.adder_32bit.operator_A_23.B ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_A_24.G = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_24.A & \multiplier_16x16bit_pipelined.adder_32bit.operator_A_24.B ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_A_24.P = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_24.A ^ \multiplier_16x16bit_pipelined.adder_32bit.operator_A_24.B ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_A_26.G = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_26.A & \multiplier_16x16bit_pipelined.adder_32bit.operator_A_26.B ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_A_26.P = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_26.A ^ \multiplier_16x16bit_pipelined.adder_32bit.operator_A_26.B ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_A_28.G = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_28.A & \multiplier_16x16bit_pipelined.reg_layer_2_w28 ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_A_28.P = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_28.A ^ \multiplier_16x16bit_pipelined.reg_layer_2_w28 ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_A_3.G = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_3.A & \multiplier_16x16bit_pipelined.adder_32bit.operator_A_3.B ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_A_3.P = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_3.A ^ \multiplier_16x16bit_pipelined.adder_32bit.operator_A_3.B ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_A_30.G = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_30.A & \multiplier_16x16bit_pipelined.reg_layer_2_w30 ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_A_30.P = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_30.A ^ \multiplier_16x16bit_pipelined.reg_layer_2_w30 ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_A_4.G = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_4.A & \multiplier_16x16bit_pipelined.adder_32bit.operator_A_4.B ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_A_4.P = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_4.A ^ \multiplier_16x16bit_pipelined.adder_32bit.operator_A_4.B ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_A_5.G = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_5.A & \multiplier_16x16bit_pipelined.adder_32bit.operator_A_5.B ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_A_5.P = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_5.A ^ \multiplier_16x16bit_pipelined.adder_32bit.operator_A_5.B ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_A_6.G = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_6.A & \multiplier_16x16bit_pipelined.adder_32bit.operator_A_6.B ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_A_6.P = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_6.A ^ \multiplier_16x16bit_pipelined.adder_32bit.operator_A_6.B ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_A_7.G = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_7.A & \multiplier_16x16bit_pipelined.adder_32bit.operator_A_7.B ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_A_7.P = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_7.A ^ \multiplier_16x16bit_pipelined.adder_32bit.operator_A_7.B ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_A_8.G = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_8.A & \multiplier_16x16bit_pipelined.adder_32bit.operator_A_8.B ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_A_8.P = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_8.A ^ \multiplier_16x16bit_pipelined.adder_32bit.operator_A_8.B ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_A_9.G = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_9.A & \multiplier_16x16bit_pipelined.adder_32bit.operator_A_9.B ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_A_9.P = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_9.A ^ \multiplier_16x16bit_pipelined.adder_32bit.operator_A_9.B ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_1.Po = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_2.A & \multiplier_16x16bit_pipelined.reg_layer_2_w1 ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_10.Po = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_20.P & \multiplier_16x16bit_pipelined.adder_32bit.operator_A_19.P ;
  assign _0280_ = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_20.P & \multiplier_16x16bit_pipelined.adder_32bit.operator_A_19.G ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_10.Go = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_20.G | _0280_;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_11.Po = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_22.P & \multiplier_16x16bit_pipelined.adder_32bit.operator_A_21.P ;
  assign _0281_ = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_22.P & \multiplier_16x16bit_pipelined.adder_32bit.operator_A_21.G ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_11.Go = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_22.G | _0281_;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_12.Po = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_24.P & \multiplier_16x16bit_pipelined.adder_32bit.operator_A_23.P ;
  assign _0282_ = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_24.P & \multiplier_16x16bit_pipelined.adder_32bit.operator_A_23.G ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_12.Go = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_24.G | _0282_;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_13.Po = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_26.P & \multiplier_16x16bit_pipelined.adder_32bit.operator_A_25.A ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_14.Po = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_28.P & \multiplier_16x16bit_pipelined.adder_32bit.operator_A_27.A ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_15.Po = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_30.P & \multiplier_16x16bit_pipelined.adder_32bit.operator_A_29.A ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_2.Po = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_4.P & \multiplier_16x16bit_pipelined.adder_32bit.operator_A_3.P ;
  assign _0283_ = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_4.P & \multiplier_16x16bit_pipelined.adder_32bit.operator_A_3.G ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_2.Go = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_4.G | _0283_;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_3.Po = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_6.P & \multiplier_16x16bit_pipelined.adder_32bit.operator_A_5.P ;
  assign _0284_ = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_6.P & \multiplier_16x16bit_pipelined.adder_32bit.operator_A_5.G ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_3.Go = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_6.G | _0284_;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_4.Po = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_8.P & \multiplier_16x16bit_pipelined.adder_32bit.operator_A_7.P ;
  assign _0285_ = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_8.P & \multiplier_16x16bit_pipelined.adder_32bit.operator_A_7.G ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_4.Go = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_8.G | _0285_;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_5.Po = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_10.P & \multiplier_16x16bit_pipelined.adder_32bit.operator_A_9.P ;
  assign _0286_ = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_10.P & \multiplier_16x16bit_pipelined.adder_32bit.operator_A_9.G ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_5.Go = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_10.G | _0286_;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_6.Po = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_12.P & \multiplier_16x16bit_pipelined.adder_32bit.operator_A_11.P ;
  assign _0287_ = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_12.P & \multiplier_16x16bit_pipelined.adder_32bit.operator_A_11.G ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_6.Go = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_12.G | _0287_;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_7.Po = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_14.P & \multiplier_16x16bit_pipelined.adder_32bit.operator_A_13.P ;
  assign _0288_ = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_14.P & \multiplier_16x16bit_pipelined.adder_32bit.operator_A_13.G ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_7.Go = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_14.G | _0288_;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_8.Po = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_16.P & \multiplier_16x16bit_pipelined.adder_32bit.operator_A_15.P ;
  assign _0289_ = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_16.P & \multiplier_16x16bit_pipelined.adder_32bit.operator_A_15.G ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_8.Go = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_16.G | _0289_;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_9.Po = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_18.P & \multiplier_16x16bit_pipelined.adder_32bit.operator_A_17.P ;
  assign _0290_ = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_18.P & \multiplier_16x16bit_pipelined.adder_32bit.operator_A_17.G ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_9.Go = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_18.G | _0290_;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_10.Po = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_10.Po & \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_9.Po ;
  assign _0291_ = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_10.Po & \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_9.Go ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_10.Go = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_10.Go | _0291_;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_11.Po = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_11.Po & \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_10.Po ;
  assign _0292_ = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_11.Po & \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_10.Go ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_11.Go = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_11.Go | _0292_;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_12.Po = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_12.Po & \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_11.Po ;
  assign _0293_ = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_12.Po & \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_11.Go ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_12.Go = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_12.Go | _0293_;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_13.Po = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_13.Po & \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_12.Po ;
  assign _0294_ = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_13.Po & \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_12.Go ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_13.Go = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_26.G | _0294_;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_14.Po = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_14.Po & \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_13.Po ;
  assign _0295_ = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_14.Po & \multiplier_16x16bit_pipelined.adder_32bit.operator_A_26.G ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_14.Go = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_28.G | _0295_;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_15.Po = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_15.Po & \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_14.Po ;
  assign _0296_ = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_15.Po & \multiplier_16x16bit_pipelined.adder_32bit.operator_A_28.G ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_15.Go = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_30.G | _0296_;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_2.Po = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_2.Po & \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_1.Po ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_3.Po = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_3.Po & \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_2.Po ;
  assign _0297_ = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_3.Po & \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_2.Go ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_3.Go = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_3.Go | _0297_;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_4.Po = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_4.Po & \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_3.Po ;
  assign _0298_ = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_4.Po & \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_3.Go ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_4.Go = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_4.Go | _0298_;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_5.Po = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_5.Po & \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_4.Po ;
  assign _0299_ = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_5.Po & \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_4.Go ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_5.Go = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_5.Go | _0299_;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_6.Po = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_6.Po & \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_5.Po ;
  assign _0300_ = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_6.Po & \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_5.Go ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_6.Go = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_6.Go | _0300_;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_7.Po = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_7.Po & \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_6.Po ;
  assign _0301_ = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_7.Po & \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_6.Go ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_7.Go = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_7.Go | _0301_;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_8.Po = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_8.Po & \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_7.Po ;
  assign _0302_ = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_8.Po & \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_7.Go ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_8.Go = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_8.Go | _0302_;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_9.Po = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_9.Po & \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_8.Po ;
  assign _0303_ = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_9.Po & \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_8.Go ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_9.Go = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_9.Go | _0303_;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_10.Po = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_10.Po & \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_8.Po ;
  assign _0304_ = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_10.Po & \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_8.Go ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_10.Go = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_10.Go | _0304_;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_11.Po = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_11.Po & \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_9.Po ;
  assign _0305_ = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_11.Po & \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_9.Go ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_11.Go = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_11.Go | _0305_;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_12.Po = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_12.Po & \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_10.Po ;
  assign _0306_ = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_12.Po & \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_10.Go ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_12.Go = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_12.Go | _0306_;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_13.Po = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_13.Po & \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_11.Po ;
  assign _0307_ = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_13.Po & \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_11.Go ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_13.Go = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_13.Go | _0307_;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_14.Po = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_14.Po & \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_12.Po ;
  assign _0308_ = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_14.Po & \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_12.Go ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_14.Go = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_14.Go | _0308_;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_15.Po = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_15.Po & \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_13.Po ;
  assign _0309_ = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_15.Po & \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_13.Go ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_15.Go = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_15.Go | _0309_;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_4.Po = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_4.Po & \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_2.Po ;
  assign _0310_ = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_4.Po & \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_2.Go ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_4.Go = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_4.Go | _0310_;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_5.Po = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_5.Po & \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_3.Po ;
  assign _0311_ = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_5.Po & \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_3.Go ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_5.Go = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_5.Go | _0311_;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_6.Po = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_6.Po & \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_4.Po ;
  assign _0312_ = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_6.Po & \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_4.Go ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_6.Go = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_6.Go | _0312_;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_7.Po = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_7.Po & \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_5.Po ;
  assign _0313_ = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_7.Po & \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_5.Go ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_7.Go = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_7.Go | _0313_;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_8.Po = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_8.Po & \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_6.Po ;
  assign _0314_ = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_8.Po & \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_6.Go ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_8.Go = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_8.Go | _0314_;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_9.Po = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_9.Po & \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_7.Po ;
  assign _0315_ = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_9.Po & \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_7.Go ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_9.Go = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_9.Go | _0315_;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_4_10.Po = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_10.Po & \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_6.Po ;
  assign _0316_ = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_10.Po & \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_6.Go ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_4_10.Go = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_10.Go | _0316_;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_4_11.Po = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_11.Po & \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_7.Po ;
  assign _0317_ = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_11.Po & \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_7.Go ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_4_11.Go = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_11.Go | _0317_;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_4_12.Po = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_12.Po & \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_8.Po ;
  assign _0318_ = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_12.Po & \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_8.Go ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_4_12.Go = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_12.Go | _0318_;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_4_13.Po = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_13.Po & \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_9.Po ;
  assign _0319_ = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_13.Po & \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_9.Go ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_4_13.Go = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_13.Go | _0319_;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_4_14.Po = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_14.Po & \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_10.Po ;
  assign _0320_ = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_14.Po & \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_10.Go ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_4_14.Go = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_14.Go | _0320_;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_4_15.Po = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_15.Po & \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_11.Po ;
  assign _0321_ = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_15.Po & \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_11.Go ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_4_15.Go = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_15.Go | _0321_;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_4_8.Po = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_8.Po & \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_4.Po ;
  assign _0322_ = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_8.Po & \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_4.Go ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_4_8.Go = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_8.Go | _0322_;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_4_9.Po = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_9.Po & \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_5.Po ;
  assign _0323_ = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_9.Po & \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_5.Go ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_4_9.Go = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_9.Go | _0323_;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_2_1.Go = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_1.Po & \multiplier_16x16bit_pipelined.adder_32bit.operator_A_0.G ;
  assign _0324_ = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_2.Po & \multiplier_16x16bit_pipelined.adder_32bit.operator_A_0.G ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_3_2.Go = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_2.Go | _0324_;
  assign _0325_ = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_3.Po & \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_2_1.Go ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_3_3.Go = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_3.Go | _0325_;
  assign _0326_ = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_4.Po & \multiplier_16x16bit_pipelined.adder_32bit.operator_A_0.G ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_4_4.Go = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_4.Go | _0326_;
  assign _0327_ = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_5.Po & \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_2_1.Go ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_4_5.Go = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_5.Go | _0327_;
  assign _0328_ = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_6.Po & \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_3_2.Go ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_4_6.Go = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_6.Go | _0328_;
  assign _0329_ = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_7.Po & \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_3_3.Go ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_4_7.Go = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_7.Go | _0329_;
  assign _0330_ = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_4_10.Po & \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_3_2.Go ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_5_10.Go = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_4_10.Go | _0330_;
  assign _0331_ = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_4_11.Po & \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_3_3.Go ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_5_11.Go = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_4_11.Go | _0331_;
  assign _0332_ = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_4_12.Po & \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_4_4.Go ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_5_12.Go = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_4_12.Go | _0332_;
  assign _0333_ = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_4_13.Po & \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_4_5.Go ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_5_13.Go = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_4_13.Go | _0333_;
  assign _0334_ = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_4_14.Po & \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_4_6.Go ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_5_14.Go = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_4_14.Go | _0334_;
  assign _0335_ = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_4_15.Po & \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_4_7.Go ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_5_15.Go = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_4_15.Go | _0335_;
  assign _0336_ = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_4_8.Po & \multiplier_16x16bit_pipelined.adder_32bit.operator_A_0.G ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_5_8.Go = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_4_8.Go | _0336_;
  assign _0337_ = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_4_9.Po & \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_2_1.Go ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_5_9.Go = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_4_9.Go | _0337_;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_6_0.Go = \multiplier_16x16bit_pipelined.reg_layer_2_w1 & \multiplier_16x16bit_pipelined.adder_32bit.operator_A_0.G ;
  assign _0338_ = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_3.P & \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_2_1.Go ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_6_1.Go = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_3.G | _0338_;
  assign _0339_ = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_21.P & \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_5_10.Go ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_6_10.Go = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_21.G | _0339_;
  assign _0340_ = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_23.P & \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_5_11.Go ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_6_11.Go = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_23.G | _0340_;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_6_12.Go = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_25.A & \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_5_12.Go ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_6_13.Go = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_27.A & \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_5_13.Go ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_6_14.Go = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_29.A & \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_5_14.Go ;
  assign _0341_ = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_5.P & \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_3_2.Go ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_6_2.Go = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_5.G | _0341_;
  assign _0342_ = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_7.P & \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_3_3.Go ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_6_3.Go = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_7.G | _0342_;
  assign _0343_ = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_9.P & \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_4_4.Go ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_6_4.Go = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_9.G | _0343_;
  assign _0344_ = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_11.P & \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_4_5.Go ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_6_5.Go = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_11.G | _0344_;
  assign _0345_ = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_13.P & \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_4_6.Go ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_6_6.Go = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_13.G | _0345_;
  assign _0346_ = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_15.P & \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_4_7.Go ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_6_7.Go = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_15.G | _0346_;
  assign _0347_ = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_17.P & \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_5_8.Go ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_6_8.Go = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_17.G | _0347_;
  assign _0348_ = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_19.P & \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_5_9.Go ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_6_9.Go = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_19.G | _0348_;
  assign \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_0.double = \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_0.nB & \multiplier_16x16bit_pipelined.mr [1];
  assign \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_0.zero = \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_0.nA & \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_0.nB ;
  assign \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_0.nB = ~ \multiplier_16x16bit_pipelined.mr [0];
  assign \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_0.nA = ~ \multiplier_16x16bit_pipelined.mr [1];
  assign \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_1.BC = \multiplier_16x16bit_pipelined.mr [2] & \multiplier_16x16bit_pipelined.mr [1];
  assign \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_1.nBnC = \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_1.nB & \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_0.nA ;
  assign _0349_ = \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_1.nBnC & \multiplier_16x16bit_pipelined.mr [3];
  assign _0350_ = \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_1.BC & \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_1.nA ;
  assign \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_1.negation = \multiplier_16x16bit_pipelined.mr [3] & \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_1.nBanC ;
  assign _0351_ = \multiplier_16x16bit_pipelined.mr [3] & \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_1.BC ;
  assign _0352_ = \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_1.nA & \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_1.nBnC ;
  assign \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_1.nB = ~ \multiplier_16x16bit_pipelined.mr [2];
  assign \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_1.nA = ~ \multiplier_16x16bit_pipelined.mr [3];
  assign \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_1.nBanC = \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_1.nB | \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_0.nA ;
  assign \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_1.double = _0349_ | _0350_;
  assign \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_1.zero = _0351_ | _0352_;
  assign \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_2.BC = \multiplier_16x16bit_pipelined.mr [4] & \multiplier_16x16bit_pipelined.mr [3];
  assign \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_2.nBnC = \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_2.nB & \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_1.nA ;
  assign _0353_ = \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_2.nBnC & \multiplier_16x16bit_pipelined.mr [5];
  assign _0354_ = \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_2.BC & \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_2.nA ;
  assign \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_2.negation = \multiplier_16x16bit_pipelined.mr [5] & \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_2.nBanC ;
  assign _0355_ = \multiplier_16x16bit_pipelined.mr [5] & \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_2.BC ;
  assign _0356_ = \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_2.nA & \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_2.nBnC ;
  assign \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_2.nB = ~ \multiplier_16x16bit_pipelined.mr [4];
  assign \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_2.nA = ~ \multiplier_16x16bit_pipelined.mr [5];
  assign \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_2.nBanC = \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_2.nB | \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_1.nA ;
  assign \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_2.double = _0353_ | _0354_;
  assign \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_2.zero = _0355_ | _0356_;
  assign \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_3.BC = \multiplier_16x16bit_pipelined.mr [6] & \multiplier_16x16bit_pipelined.mr [5];
  assign \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_3.nBnC = \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_3.nB & \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_2.nA ;
  assign _0357_ = \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_3.nBnC & \multiplier_16x16bit_pipelined.mr [7];
  assign _0358_ = \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_3.BC & \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_3.nA ;
  assign \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_3.negation = \multiplier_16x16bit_pipelined.mr [7] & \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_3.nBanC ;
  assign _0359_ = \multiplier_16x16bit_pipelined.mr [7] & \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_3.BC ;
  assign _0360_ = \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_3.nA & \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_3.nBnC ;
  assign \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_3.nB = ~ \multiplier_16x16bit_pipelined.mr [6];
  assign \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_3.nA = ~ \multiplier_16x16bit_pipelined.mr [7];
  assign \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_3.nBanC = \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_3.nB | \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_2.nA ;
  assign \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_3.double = _0357_ | _0358_;
  assign \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_3.zero = _0359_ | _0360_;
  assign \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_4.BC = \multiplier_16x16bit_pipelined.mr [8] & \multiplier_16x16bit_pipelined.mr [7];
  assign \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_4.nBnC = \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_4.nB & \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_3.nA ;
  assign _0361_ = \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_4.nBnC & \multiplier_16x16bit_pipelined.mr [9];
  assign _0362_ = \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_4.BC & \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_4.nA ;
  assign \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_4.negation = \multiplier_16x16bit_pipelined.mr [9] & \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_4.nBanC ;
  assign _0363_ = \multiplier_16x16bit_pipelined.mr [9] & \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_4.BC ;
  assign _0364_ = \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_4.nA & \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_4.nBnC ;
  assign \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_4.nB = ~ \multiplier_16x16bit_pipelined.mr [8];
  assign \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_4.nA = ~ \multiplier_16x16bit_pipelined.mr [9];
  assign \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_4.nBanC = \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_4.nB | \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_3.nA ;
  assign \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_4.double = _0361_ | _0362_;
  assign \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_4.zero = _0363_ | _0364_;
  assign \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_5.BC = \multiplier_16x16bit_pipelined.mr [10] & \multiplier_16x16bit_pipelined.mr [9];
  assign \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_5.nBnC = \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_5.nB & \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_4.nA ;
  assign _0365_ = \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_5.nBnC & \multiplier_16x16bit_pipelined.mr [11];
  assign _0366_ = \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_5.BC & \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_5.nA ;
  assign \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_5.negation = \multiplier_16x16bit_pipelined.mr [11] & \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_5.nBanC ;
  assign _0367_ = \multiplier_16x16bit_pipelined.mr [11] & \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_5.BC ;
  assign _0368_ = \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_5.nA & \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_5.nBnC ;
  assign \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_5.nB = ~ \multiplier_16x16bit_pipelined.mr [10];
  assign \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_5.nA = ~ \multiplier_16x16bit_pipelined.mr [11];
  assign \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_5.nBanC = \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_5.nB | \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_4.nA ;
  assign \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_5.double = _0365_ | _0366_;
  assign \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_5.zero = _0367_ | _0368_;
  assign \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_6.BC = \multiplier_16x16bit_pipelined.mr [12] & \multiplier_16x16bit_pipelined.mr [11];
  assign \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_6.nBnC = \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_6.nB & \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_5.nA ;
  assign _0369_ = \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_6.nBnC & \multiplier_16x16bit_pipelined.mr [13];
  assign _0370_ = \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_6.BC & \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_6.nA ;
  assign \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_6.negation = \multiplier_16x16bit_pipelined.mr [13] & \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_6.nBanC ;
  assign _0371_ = \multiplier_16x16bit_pipelined.mr [13] & \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_6.BC ;
  assign _0372_ = \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_6.nA & \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_6.nBnC ;
  assign \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_6.nB = ~ \multiplier_16x16bit_pipelined.mr [12];
  assign \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_6.nA = ~ \multiplier_16x16bit_pipelined.mr [13];
  assign \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_6.nBanC = \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_6.nB | \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_5.nA ;
  assign \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_6.double = _0369_ | _0370_;
  assign \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_6.zero = _0371_ | _0372_;
  assign \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_7.BC = \multiplier_16x16bit_pipelined.mr [14] & \multiplier_16x16bit_pipelined.mr [13];
  assign \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_7.nBnC = \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_7.nB & \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_6.nA ;
  assign _0373_ = \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_7.nBnC & \multiplier_16x16bit_pipelined.mr [15];
  assign _0374_ = \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_7.BC & \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_7.nA ;
  assign \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_7.negation = \multiplier_16x16bit_pipelined.mr [15] & \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_7.nBanC ;
  assign _0375_ = \multiplier_16x16bit_pipelined.mr [15] & \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_7.BC ;
  assign _0376_ = \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_7.nA & \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_7.nBnC ;
  assign \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_7.nB = ~ \multiplier_16x16bit_pipelined.mr [14];
  assign \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_7.nA = ~ \multiplier_16x16bit_pipelined.mr [15];
  assign \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_7.nBanC = \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_7.nB | \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_6.nA ;
  assign \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_7.double = _0373_ | _0374_;
  assign \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_7.zero = _0375_ | _0376_;
  assign \multiplier_16x16bit_pipelined.layer_1_compressor42_0.AB = \multiplier_16x16bit_pipelined.layer_1_compressor42_0.A & \multiplier_16x16bit_pipelined.layer_1_compressor42_0.B ;
  assign \multiplier_16x16bit_pipelined.layer_1_compressor42_0.CD = \multiplier_16x16bit_pipelined.layer_1_compressor42_0.C & \multiplier_16x16bit_pipelined.layer_1_compressor42_0.D ;
  assign _0377_ = \multiplier_16x16bit_pipelined.layer_1_compressor42_0.AB & \multiplier_16x16bit_pipelined.layer_1_compressor42_0.CD ;
  assign _0378_ = \multiplier_16x16bit_pipelined.layer_1_compressor42_0.AxorB & \multiplier_16x16bit_pipelined.layer_1_compressor42_0.CxorD ;
  assign _0379_ = \multiplier_16x16bit_pipelined.layer_1_compressor42_0.AxBxCxD & \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_3.negation ;
  assign \multiplier_16x16bit_pipelined.layer_1_compressor42_0.cout = \multiplier_16x16bit_pipelined.layer_1_compressor42_0.AB | \multiplier_16x16bit_pipelined.layer_1_compressor42_0.CD ;
  assign _0380_ = _0377_ | _0378_;
  assign \multiplier_16x16bit_pipelined.layer_1_compressor42_0.carry = _0380_ | _0379_;
  assign \multiplier_16x16bit_pipelined.layer_1_compressor42_0.AxorB = \multiplier_16x16bit_pipelined.layer_1_compressor42_0.A ^ \multiplier_16x16bit_pipelined.layer_1_compressor42_0.B ;
  assign \multiplier_16x16bit_pipelined.layer_1_compressor42_0.CxorD = \multiplier_16x16bit_pipelined.layer_1_compressor42_0.C ^ \multiplier_16x16bit_pipelined.layer_1_compressor42_0.D ;
  assign \multiplier_16x16bit_pipelined.layer_1_compressor42_0.AxBxCxD = \multiplier_16x16bit_pipelined.layer_1_compressor42_0.AxorB ^ \multiplier_16x16bit_pipelined.layer_1_compressor42_0.CxorD ;
  assign \multiplier_16x16bit_pipelined.layer_1_compressor42_0.S = \multiplier_16x16bit_pipelined.layer_1_compressor42_0.AxBxCxD ^ \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_3.negation ;
  assign \multiplier_16x16bit_pipelined.layer_1_compressor42_1.AB = \multiplier_16x16bit_pipelined.layer_1_compressor42_1.A & \multiplier_16x16bit_pipelined.layer_1_compressor42_1.B ;
  assign \multiplier_16x16bit_pipelined.layer_1_compressor42_1.CD = \multiplier_16x16bit_pipelined.layer_1_compressor42_1.C & \multiplier_16x16bit_pipelined.layer_1_compressor42_1.D ;
  assign _0381_ = \multiplier_16x16bit_pipelined.layer_1_compressor42_1.AB & \multiplier_16x16bit_pipelined.layer_1_compressor42_1.CD ;
  assign _0382_ = \multiplier_16x16bit_pipelined.layer_1_compressor42_1.AxorB & \multiplier_16x16bit_pipelined.layer_1_compressor42_1.CxorD ;
  assign _0383_ = \multiplier_16x16bit_pipelined.layer_1_compressor42_1.AxBxCxD & \multiplier_16x16bit_pipelined.layer_1_compressor42_1.cin ;
  assign \multiplier_16x16bit_pipelined.layer_1_compressor42_1.cout = \multiplier_16x16bit_pipelined.layer_1_compressor42_1.AB | \multiplier_16x16bit_pipelined.layer_1_compressor42_1.CD ;
  assign _0384_ = _0381_ | _0382_;
  assign \multiplier_16x16bit_pipelined.layer_1_compressor42_1.carry = _0384_ | _0383_;
  assign \multiplier_16x16bit_pipelined.layer_1_compressor42_1.AxorB = \multiplier_16x16bit_pipelined.layer_1_compressor42_1.A ^ \multiplier_16x16bit_pipelined.layer_1_compressor42_1.B ;
  assign \multiplier_16x16bit_pipelined.layer_1_compressor42_1.CxorD = \multiplier_16x16bit_pipelined.layer_1_compressor42_1.C ^ \multiplier_16x16bit_pipelined.layer_1_compressor42_1.D ;
  assign \multiplier_16x16bit_pipelined.layer_1_compressor42_1.AxBxCxD = \multiplier_16x16bit_pipelined.layer_1_compressor42_1.AxorB ^ \multiplier_16x16bit_pipelined.layer_1_compressor42_1.CxorD ;
  assign \multiplier_16x16bit_pipelined.layer_1_compressor42_1.S = \multiplier_16x16bit_pipelined.layer_1_compressor42_1.AxBxCxD ^ \multiplier_16x16bit_pipelined.layer_1_compressor42_1.cin ;
  assign \multiplier_16x16bit_pipelined.layer_1_compressor42_10.AB = \multiplier_16x16bit_pipelined.layer_1_compressor42_10.A & \multiplier_16x16bit_pipelined.layer_1_compressor42_10.B ;
  assign \multiplier_16x16bit_pipelined.layer_1_compressor42_10.CD = \multiplier_16x16bit_pipelined.layer_1_compressor42_10.C & \multiplier_16x16bit_pipelined.layer_1_compressor42_10.D ;
  assign _0385_ = \multiplier_16x16bit_pipelined.layer_1_compressor42_10.AB & \multiplier_16x16bit_pipelined.layer_1_compressor42_10.CD ;
  assign _0386_ = \multiplier_16x16bit_pipelined.layer_1_compressor42_10.AxorB & \multiplier_16x16bit_pipelined.layer_1_compressor42_10.CxorD ;
  assign _0387_ = \multiplier_16x16bit_pipelined.layer_1_compressor42_10.AxBxCxD & \multiplier_16x16bit_pipelined.layer_1_compressor42_10.cin ;
  assign \multiplier_16x16bit_pipelined.layer_1_compressor42_10.cout = \multiplier_16x16bit_pipelined.layer_1_compressor42_10.AB | \multiplier_16x16bit_pipelined.layer_1_compressor42_10.CD ;
  assign _0388_ = _0385_ | _0386_;
  assign \multiplier_16x16bit_pipelined.layer_1_compressor42_10.carry = _0388_ | _0387_;
  assign \multiplier_16x16bit_pipelined.layer_1_compressor42_10.AxorB = \multiplier_16x16bit_pipelined.layer_1_compressor42_10.A ^ \multiplier_16x16bit_pipelined.layer_1_compressor42_10.B ;
  assign \multiplier_16x16bit_pipelined.layer_1_compressor42_10.CxorD = \multiplier_16x16bit_pipelined.layer_1_compressor42_10.C ^ \multiplier_16x16bit_pipelined.layer_1_compressor42_10.D ;
  assign \multiplier_16x16bit_pipelined.layer_1_compressor42_10.AxBxCxD = \multiplier_16x16bit_pipelined.layer_1_compressor42_10.AxorB ^ \multiplier_16x16bit_pipelined.layer_1_compressor42_10.CxorD ;
  assign \multiplier_16x16bit_pipelined.layer_1_compressor42_10.S = \multiplier_16x16bit_pipelined.layer_1_compressor42_10.AxBxCxD ^ \multiplier_16x16bit_pipelined.layer_1_compressor42_10.cin ;
  assign \multiplier_16x16bit_pipelined.layer_1_compressor42_11.AB = \multiplier_16x16bit_pipelined.layer_1_compressor42_11.A & \multiplier_16x16bit_pipelined.layer_1_compressor42_11.B ;
  assign \multiplier_16x16bit_pipelined.layer_1_compressor42_11.CD = \multiplier_16x16bit_pipelined.layer_1_compressor42_11.C & \multiplier_16x16bit_pipelined.layer_1_compressor42_11.D ;
  assign _0389_ = \multiplier_16x16bit_pipelined.layer_1_compressor42_11.AB & \multiplier_16x16bit_pipelined.layer_1_compressor42_11.CD ;
  assign _0390_ = \multiplier_16x16bit_pipelined.layer_1_compressor42_11.AxorB & \multiplier_16x16bit_pipelined.layer_1_compressor42_11.CxorD ;
  assign _0391_ = \multiplier_16x16bit_pipelined.layer_1_compressor42_11.AxBxCxD & \multiplier_16x16bit_pipelined.layer_1_compressor42_11.cin ;
  assign \multiplier_16x16bit_pipelined.layer_1_compressor42_11.cout = \multiplier_16x16bit_pipelined.layer_1_compressor42_11.AB | \multiplier_16x16bit_pipelined.layer_1_compressor42_11.CD ;
  assign _0392_ = _0389_ | _0390_;
  assign \multiplier_16x16bit_pipelined.layer_1_compressor42_11.carry = _0392_ | _0391_;
  assign \multiplier_16x16bit_pipelined.layer_1_compressor42_11.AxorB = \multiplier_16x16bit_pipelined.layer_1_compressor42_11.A ^ \multiplier_16x16bit_pipelined.layer_1_compressor42_11.B ;
  assign \multiplier_16x16bit_pipelined.layer_1_compressor42_11.CxorD = \multiplier_16x16bit_pipelined.layer_1_compressor42_11.C ^ \multiplier_16x16bit_pipelined.layer_1_compressor42_11.D ;
  assign \multiplier_16x16bit_pipelined.layer_1_compressor42_11.AxBxCxD = \multiplier_16x16bit_pipelined.layer_1_compressor42_11.AxorB ^ \multiplier_16x16bit_pipelined.layer_1_compressor42_11.CxorD ;
  assign \multiplier_16x16bit_pipelined.layer_1_compressor42_11.S = \multiplier_16x16bit_pipelined.layer_1_compressor42_11.AxBxCxD ^ \multiplier_16x16bit_pipelined.layer_1_compressor42_11.cin ;
  assign \multiplier_16x16bit_pipelined.layer_1_compressor42_12.AB = \multiplier_16x16bit_pipelined.layer_1_compressor42_12.A & \multiplier_16x16bit_pipelined.layer_1_compressor42_12.B ;
  assign \multiplier_16x16bit_pipelined.layer_1_compressor42_12.CD = \multiplier_16x16bit_pipelined.layer_1_compressor42_12.C & \multiplier_16x16bit_pipelined.layer_1_compressor42_12.D ;
  assign _0393_ = \multiplier_16x16bit_pipelined.layer_1_compressor42_12.AB & \multiplier_16x16bit_pipelined.layer_1_compressor42_12.CD ;
  assign _0394_ = \multiplier_16x16bit_pipelined.layer_1_compressor42_12.AxorB & \multiplier_16x16bit_pipelined.layer_1_compressor42_12.CxorD ;
  assign _0395_ = \multiplier_16x16bit_pipelined.layer_1_compressor42_12.AxBxCxD & \multiplier_16x16bit_pipelined.layer_1_compressor42_12.cin ;
  assign \multiplier_16x16bit_pipelined.layer_1_compressor42_12.cout = \multiplier_16x16bit_pipelined.layer_1_compressor42_12.AB | \multiplier_16x16bit_pipelined.layer_1_compressor42_12.CD ;
  assign _0396_ = _0393_ | _0394_;
  assign \multiplier_16x16bit_pipelined.layer_1_compressor42_12.carry = _0396_ | _0395_;
  assign \multiplier_16x16bit_pipelined.layer_1_compressor42_12.AxorB = \multiplier_16x16bit_pipelined.layer_1_compressor42_12.A ^ \multiplier_16x16bit_pipelined.layer_1_compressor42_12.B ;
  assign \multiplier_16x16bit_pipelined.layer_1_compressor42_12.CxorD = \multiplier_16x16bit_pipelined.layer_1_compressor42_12.C ^ \multiplier_16x16bit_pipelined.layer_1_compressor42_12.D ;
  assign \multiplier_16x16bit_pipelined.layer_1_compressor42_12.AxBxCxD = \multiplier_16x16bit_pipelined.layer_1_compressor42_12.AxorB ^ \multiplier_16x16bit_pipelined.layer_1_compressor42_12.CxorD ;
  assign \multiplier_16x16bit_pipelined.layer_1_compressor42_12.S = \multiplier_16x16bit_pipelined.layer_1_compressor42_12.AxBxCxD ^ \multiplier_16x16bit_pipelined.layer_1_compressor42_12.cin ;
  assign \multiplier_16x16bit_pipelined.layer_1_compressor42_13.AB = \multiplier_16x16bit_pipelined.layer_1_compressor42_13.A & \multiplier_16x16bit_pipelined.layer_1_compressor42_13.B ;
  assign \multiplier_16x16bit_pipelined.layer_1_compressor42_13.CD = \multiplier_16x16bit_pipelined.layer_1_compressor42_13.C & \multiplier_16x16bit_pipelined.layer_1_compressor42_13.D ;
  assign _0397_ = \multiplier_16x16bit_pipelined.layer_1_compressor42_13.AB & \multiplier_16x16bit_pipelined.layer_1_compressor42_13.CD ;
  assign _0398_ = \multiplier_16x16bit_pipelined.layer_1_compressor42_13.AxorB & \multiplier_16x16bit_pipelined.layer_1_compressor42_13.CxorD ;
  assign _0399_ = \multiplier_16x16bit_pipelined.layer_1_compressor42_13.AxBxCxD & \multiplier_16x16bit_pipelined.layer_1_compressor42_13.cin ;
  assign \multiplier_16x16bit_pipelined.layer_1_compressor42_13.cout = \multiplier_16x16bit_pipelined.layer_1_compressor42_13.AB | \multiplier_16x16bit_pipelined.layer_1_compressor42_13.CD ;
  assign _0400_ = _0397_ | _0398_;
  assign \multiplier_16x16bit_pipelined.layer_1_compressor42_13.carry = _0400_ | _0399_;
  assign \multiplier_16x16bit_pipelined.layer_1_compressor42_13.AxorB = \multiplier_16x16bit_pipelined.layer_1_compressor42_13.A ^ \multiplier_16x16bit_pipelined.layer_1_compressor42_13.B ;
  assign \multiplier_16x16bit_pipelined.layer_1_compressor42_13.CxorD = \multiplier_16x16bit_pipelined.layer_1_compressor42_13.C ^ \multiplier_16x16bit_pipelined.layer_1_compressor42_13.D ;
  assign \multiplier_16x16bit_pipelined.layer_1_compressor42_13.AxBxCxD = \multiplier_16x16bit_pipelined.layer_1_compressor42_13.AxorB ^ \multiplier_16x16bit_pipelined.layer_1_compressor42_13.CxorD ;
  assign \multiplier_16x16bit_pipelined.layer_1_compressor42_13.S = \multiplier_16x16bit_pipelined.layer_1_compressor42_13.AxBxCxD ^ \multiplier_16x16bit_pipelined.layer_1_compressor42_13.cin ;
  assign \multiplier_16x16bit_pipelined.layer_1_compressor42_14.AB = \multiplier_16x16bit_pipelined.layer_1_compressor42_14.A & \multiplier_16x16bit_pipelined.layer_1_compressor42_14.B ;
  assign \multiplier_16x16bit_pipelined.layer_1_compressor42_14.CD = \multiplier_16x16bit_pipelined.layer_1_compressor42_14.C & \multiplier_16x16bit_pipelined.layer_1_compressor42_14.D ;
  assign _0401_ = \multiplier_16x16bit_pipelined.layer_1_compressor42_14.AB & \multiplier_16x16bit_pipelined.layer_1_compressor42_14.CD ;
  assign _0402_ = \multiplier_16x16bit_pipelined.layer_1_compressor42_14.AxorB & \multiplier_16x16bit_pipelined.layer_1_compressor42_14.CxorD ;
  assign _0403_ = \multiplier_16x16bit_pipelined.layer_1_compressor42_14.AxBxCxD & \multiplier_16x16bit_pipelined.layer_1_compressor42_14.cin ;
  assign \multiplier_16x16bit_pipelined.layer_1_compressor42_14.cout = \multiplier_16x16bit_pipelined.layer_1_compressor42_14.AB | \multiplier_16x16bit_pipelined.layer_1_compressor42_14.CD ;
  assign _0404_ = _0401_ | _0402_;
  assign \multiplier_16x16bit_pipelined.layer_1_compressor42_14.carry = _0404_ | _0403_;
  assign \multiplier_16x16bit_pipelined.layer_1_compressor42_14.AxorB = \multiplier_16x16bit_pipelined.layer_1_compressor42_14.A ^ \multiplier_16x16bit_pipelined.layer_1_compressor42_14.B ;
  assign \multiplier_16x16bit_pipelined.layer_1_compressor42_14.CxorD = \multiplier_16x16bit_pipelined.layer_1_compressor42_14.C ^ \multiplier_16x16bit_pipelined.layer_1_compressor42_14.D ;
  assign \multiplier_16x16bit_pipelined.layer_1_compressor42_14.AxBxCxD = \multiplier_16x16bit_pipelined.layer_1_compressor42_14.AxorB ^ \multiplier_16x16bit_pipelined.layer_1_compressor42_14.CxorD ;
  assign \multiplier_16x16bit_pipelined.layer_1_compressor42_14.S = \multiplier_16x16bit_pipelined.layer_1_compressor42_14.AxBxCxD ^ \multiplier_16x16bit_pipelined.layer_1_compressor42_14.cin ;
  assign \multiplier_16x16bit_pipelined.layer_1_compressor42_15.AB = \multiplier_16x16bit_pipelined.layer_1_compressor42_15.A & \multiplier_16x16bit_pipelined.layer_1_compressor42_15.B ;
  assign \multiplier_16x16bit_pipelined.layer_1_compressor42_15.CD = \multiplier_16x16bit_pipelined.layer_1_compressor42_15.C & \multiplier_16x16bit_pipelined.layer_1_compressor42_15.D ;
  assign _0405_ = \multiplier_16x16bit_pipelined.layer_1_compressor42_15.AB & \multiplier_16x16bit_pipelined.layer_1_compressor42_15.CD ;
  assign _0406_ = \multiplier_16x16bit_pipelined.layer_1_compressor42_15.AxorB & \multiplier_16x16bit_pipelined.layer_1_compressor42_15.CxorD ;
  assign _0407_ = \multiplier_16x16bit_pipelined.layer_1_compressor42_15.AxBxCxD & \multiplier_16x16bit_pipelined.layer_1_compressor42_15.cin ;
  assign \multiplier_16x16bit_pipelined.layer_1_compressor42_15.cout = \multiplier_16x16bit_pipelined.layer_1_compressor42_15.AB | \multiplier_16x16bit_pipelined.layer_1_compressor42_15.CD ;
  assign _0408_ = _0405_ | _0406_;
  assign \multiplier_16x16bit_pipelined.layer_1_compressor42_15.carry = _0408_ | _0407_;
  assign \multiplier_16x16bit_pipelined.layer_1_compressor42_15.AxorB = \multiplier_16x16bit_pipelined.layer_1_compressor42_15.A ^ \multiplier_16x16bit_pipelined.layer_1_compressor42_15.B ;
  assign \multiplier_16x16bit_pipelined.layer_1_compressor42_15.CxorD = \multiplier_16x16bit_pipelined.layer_1_compressor42_15.C ^ \multiplier_16x16bit_pipelined.layer_1_compressor42_15.D ;
  assign \multiplier_16x16bit_pipelined.layer_1_compressor42_15.AxBxCxD = \multiplier_16x16bit_pipelined.layer_1_compressor42_15.AxorB ^ \multiplier_16x16bit_pipelined.layer_1_compressor42_15.CxorD ;
  assign \multiplier_16x16bit_pipelined.layer_1_compressor42_15.S = \multiplier_16x16bit_pipelined.layer_1_compressor42_15.AxBxCxD ^ \multiplier_16x16bit_pipelined.layer_1_compressor42_15.cin ;
  assign \multiplier_16x16bit_pipelined.layer_1_compressor42_16.AB = \multiplier_16x16bit_pipelined.layer_1_compressor42_16.A & \multiplier_16x16bit_pipelined.layer_1_compressor42_16.B ;
  assign \multiplier_16x16bit_pipelined.layer_1_compressor42_16.CD = \multiplier_16x16bit_pipelined.layer_1_compressor42_16.C & \multiplier_16x16bit_pipelined.layer_1_compressor42_16.D ;
  assign _0409_ = \multiplier_16x16bit_pipelined.layer_1_compressor42_16.AB & \multiplier_16x16bit_pipelined.layer_1_compressor42_16.CD ;
  assign _0410_ = \multiplier_16x16bit_pipelined.layer_1_compressor42_16.AxorB & \multiplier_16x16bit_pipelined.layer_1_compressor42_16.CxorD ;
  assign \multiplier_16x16bit_pipelined.layer_1_compressor42_16.cout = \multiplier_16x16bit_pipelined.layer_1_compressor42_16.AB | \multiplier_16x16bit_pipelined.layer_1_compressor42_16.CD ;
  assign _0411_ = _0409_ | _0410_;
  assign \multiplier_16x16bit_pipelined.layer_1_compressor42_16.carry = _0411_ | \multiplier_16x16bit_pipelined.layer_1_compressor42_16.AxBxCxD ;
  assign \multiplier_16x16bit_pipelined.layer_1_compressor42_16.AxorB = \multiplier_16x16bit_pipelined.layer_1_compressor42_16.A ^ \multiplier_16x16bit_pipelined.layer_1_compressor42_16.B ;
  assign \multiplier_16x16bit_pipelined.layer_1_compressor42_16.CxorD = \multiplier_16x16bit_pipelined.layer_1_compressor42_16.C ^ \multiplier_16x16bit_pipelined.layer_1_compressor42_16.D ;
  assign \multiplier_16x16bit_pipelined.layer_1_compressor42_16.AxBxCxD = \multiplier_16x16bit_pipelined.layer_1_compressor42_16.AxorB ^ \multiplier_16x16bit_pipelined.layer_1_compressor42_16.CxorD ;
  assign \multiplier_16x16bit_pipelined.layer_1_compressor42_16.S = \multiplier_16x16bit_pipelined.layer_1_compressor42_16.AxBxCxD ^ 1'b1;
  assign \multiplier_16x16bit_pipelined.layer_1_compressor42_2.AB = \multiplier_16x16bit_pipelined.layer_1_compressor42_2.A & \multiplier_16x16bit_pipelined.layer_1_compressor42_2.B ;
  assign \multiplier_16x16bit_pipelined.layer_1_compressor42_2.CD = \multiplier_16x16bit_pipelined.layer_1_compressor42_2.C & \multiplier_16x16bit_pipelined.layer_1_compressor42_2.D ;
  assign _0412_ = \multiplier_16x16bit_pipelined.layer_1_compressor42_2.AB & \multiplier_16x16bit_pipelined.layer_1_compressor42_2.CD ;
  assign _0413_ = \multiplier_16x16bit_pipelined.layer_1_compressor42_2.AxorB & \multiplier_16x16bit_pipelined.layer_1_compressor42_2.CxorD ;
  assign _0414_ = \multiplier_16x16bit_pipelined.layer_1_compressor42_2.AxBxCxD & \multiplier_16x16bit_pipelined.layer_1_compressor42_2.cin ;
  assign \multiplier_16x16bit_pipelined.layer_1_compressor42_2.cout = \multiplier_16x16bit_pipelined.layer_1_compressor42_2.AB | \multiplier_16x16bit_pipelined.layer_1_compressor42_2.CD ;
  assign _0415_ = _0412_ | _0413_;
  assign \multiplier_16x16bit_pipelined.layer_1_compressor42_2.carry = _0415_ | _0414_;
  assign \multiplier_16x16bit_pipelined.layer_1_compressor42_2.AxorB = \multiplier_16x16bit_pipelined.layer_1_compressor42_2.A ^ \multiplier_16x16bit_pipelined.layer_1_compressor42_2.B ;
  assign \multiplier_16x16bit_pipelined.layer_1_compressor42_2.CxorD = \multiplier_16x16bit_pipelined.layer_1_compressor42_2.C ^ \multiplier_16x16bit_pipelined.layer_1_compressor42_2.D ;
  assign \multiplier_16x16bit_pipelined.layer_1_compressor42_2.AxBxCxD = \multiplier_16x16bit_pipelined.layer_1_compressor42_2.AxorB ^ \multiplier_16x16bit_pipelined.layer_1_compressor42_2.CxorD ;
  assign \multiplier_16x16bit_pipelined.layer_1_compressor42_2.S = \multiplier_16x16bit_pipelined.layer_1_compressor42_2.AxBxCxD ^ \multiplier_16x16bit_pipelined.layer_1_compressor42_2.cin ;
  assign \multiplier_16x16bit_pipelined.layer_1_compressor42_3.AB = \multiplier_16x16bit_pipelined.layer_1_compressor42_3.A & \multiplier_16x16bit_pipelined.layer_1_compressor42_3.B ;
  assign \multiplier_16x16bit_pipelined.layer_1_compressor42_3.CD = \multiplier_16x16bit_pipelined.layer_1_compressor42_3.C & \multiplier_16x16bit_pipelined.layer_1_compressor42_3.D ;
  assign _0416_ = \multiplier_16x16bit_pipelined.layer_1_compressor42_3.AB & \multiplier_16x16bit_pipelined.layer_1_compressor42_3.CD ;
  assign _0417_ = \multiplier_16x16bit_pipelined.layer_1_compressor42_3.AxorB & \multiplier_16x16bit_pipelined.layer_1_compressor42_3.CxorD ;
  assign _0418_ = \multiplier_16x16bit_pipelined.layer_1_compressor42_3.AxBxCxD & \multiplier_16x16bit_pipelined.layer_1_compressor42_3.cin ;
  assign \multiplier_16x16bit_pipelined.layer_1_compressor42_3.cout = \multiplier_16x16bit_pipelined.layer_1_compressor42_3.AB | \multiplier_16x16bit_pipelined.layer_1_compressor42_3.CD ;
  assign _0419_ = _0416_ | _0417_;
  assign \multiplier_16x16bit_pipelined.layer_1_compressor42_3.carry = _0419_ | _0418_;
  assign \multiplier_16x16bit_pipelined.layer_1_compressor42_3.AxorB = \multiplier_16x16bit_pipelined.layer_1_compressor42_3.A ^ \multiplier_16x16bit_pipelined.layer_1_compressor42_3.B ;
  assign \multiplier_16x16bit_pipelined.layer_1_compressor42_3.CxorD = \multiplier_16x16bit_pipelined.layer_1_compressor42_3.C ^ \multiplier_16x16bit_pipelined.layer_1_compressor42_3.D ;
  assign \multiplier_16x16bit_pipelined.layer_1_compressor42_3.AxBxCxD = \multiplier_16x16bit_pipelined.layer_1_compressor42_3.AxorB ^ \multiplier_16x16bit_pipelined.layer_1_compressor42_3.CxorD ;
  assign \multiplier_16x16bit_pipelined.layer_1_compressor42_3.S = \multiplier_16x16bit_pipelined.layer_1_compressor42_3.AxBxCxD ^ \multiplier_16x16bit_pipelined.layer_1_compressor42_3.cin ;
  assign \multiplier_16x16bit_pipelined.layer_1_compressor42_4.AB = \multiplier_16x16bit_pipelined.layer_1_compressor42_4.A & \multiplier_16x16bit_pipelined.layer_1_compressor42_4.B ;
  assign \multiplier_16x16bit_pipelined.layer_1_compressor42_4.CD = \multiplier_16x16bit_pipelined.layer_1_compressor42_4.C & \multiplier_16x16bit_pipelined.layer_1_compressor42_4.D ;
  assign _0420_ = \multiplier_16x16bit_pipelined.layer_1_compressor42_4.AB & \multiplier_16x16bit_pipelined.layer_1_compressor42_4.CD ;
  assign _0421_ = \multiplier_16x16bit_pipelined.layer_1_compressor42_4.AxorB & \multiplier_16x16bit_pipelined.layer_1_compressor42_4.CxorD ;
  assign _0422_ = \multiplier_16x16bit_pipelined.layer_1_compressor42_4.AxBxCxD & \multiplier_16x16bit_pipelined.layer_1_compressor42_4.cin ;
  assign \multiplier_16x16bit_pipelined.layer_1_compressor42_4.cout = \multiplier_16x16bit_pipelined.layer_1_compressor42_4.AB | \multiplier_16x16bit_pipelined.layer_1_compressor42_4.CD ;
  assign _0423_ = _0420_ | _0421_;
  assign \multiplier_16x16bit_pipelined.layer_1_compressor42_4.carry = _0423_ | _0422_;
  assign \multiplier_16x16bit_pipelined.layer_1_compressor42_4.AxorB = \multiplier_16x16bit_pipelined.layer_1_compressor42_4.A ^ \multiplier_16x16bit_pipelined.layer_1_compressor42_4.B ;
  assign \multiplier_16x16bit_pipelined.layer_1_compressor42_4.CxorD = \multiplier_16x16bit_pipelined.layer_1_compressor42_4.C ^ \multiplier_16x16bit_pipelined.layer_1_compressor42_4.D ;
  assign \multiplier_16x16bit_pipelined.layer_1_compressor42_4.AxBxCxD = \multiplier_16x16bit_pipelined.layer_1_compressor42_4.AxorB ^ \multiplier_16x16bit_pipelined.layer_1_compressor42_4.CxorD ;
  assign \multiplier_16x16bit_pipelined.layer_1_compressor42_4.S = \multiplier_16x16bit_pipelined.layer_1_compressor42_4.AxBxCxD ^ \multiplier_16x16bit_pipelined.layer_1_compressor42_4.cin ;
  assign \multiplier_16x16bit_pipelined.layer_1_compressor42_5.AB = \multiplier_16x16bit_pipelined.layer_1_compressor42_5.A & \multiplier_16x16bit_pipelined.layer_1_compressor42_5.B ;
  assign \multiplier_16x16bit_pipelined.layer_1_compressor42_5.CD = \multiplier_16x16bit_pipelined.layer_1_compressor42_5.C & \multiplier_16x16bit_pipelined.layer_1_compressor42_5.D ;
  assign _0424_ = \multiplier_16x16bit_pipelined.layer_1_compressor42_5.AB & \multiplier_16x16bit_pipelined.layer_1_compressor42_5.CD ;
  assign _0425_ = \multiplier_16x16bit_pipelined.layer_1_compressor42_5.AxorB & \multiplier_16x16bit_pipelined.layer_1_compressor42_5.CxorD ;
  assign _0426_ = \multiplier_16x16bit_pipelined.layer_1_compressor42_5.AxBxCxD & \multiplier_16x16bit_pipelined.layer_1_compressor42_5.cin ;
  assign \multiplier_16x16bit_pipelined.layer_1_compressor42_5.cout = \multiplier_16x16bit_pipelined.layer_1_compressor42_5.AB | \multiplier_16x16bit_pipelined.layer_1_compressor42_5.CD ;
  assign _0427_ = _0424_ | _0425_;
  assign \multiplier_16x16bit_pipelined.layer_1_compressor42_5.carry = _0427_ | _0426_;
  assign \multiplier_16x16bit_pipelined.layer_1_compressor42_5.AxorB = \multiplier_16x16bit_pipelined.layer_1_compressor42_5.A ^ \multiplier_16x16bit_pipelined.layer_1_compressor42_5.B ;
  assign \multiplier_16x16bit_pipelined.layer_1_compressor42_5.CxorD = \multiplier_16x16bit_pipelined.layer_1_compressor42_5.C ^ \multiplier_16x16bit_pipelined.layer_1_compressor42_5.D ;
  assign \multiplier_16x16bit_pipelined.layer_1_compressor42_5.AxBxCxD = \multiplier_16x16bit_pipelined.layer_1_compressor42_5.AxorB ^ \multiplier_16x16bit_pipelined.layer_1_compressor42_5.CxorD ;
  assign \multiplier_16x16bit_pipelined.layer_1_compressor42_5.S = \multiplier_16x16bit_pipelined.layer_1_compressor42_5.AxBxCxD ^ \multiplier_16x16bit_pipelined.layer_1_compressor42_5.cin ;
  assign \multiplier_16x16bit_pipelined.layer_1_compressor42_6.AB = \multiplier_16x16bit_pipelined.layer_1_compressor42_6.A & \multiplier_16x16bit_pipelined.layer_1_compressor42_6.B ;
  assign \multiplier_16x16bit_pipelined.layer_1_compressor42_6.CD = \multiplier_16x16bit_pipelined.layer_1_compressor42_6.C & \multiplier_16x16bit_pipelined.layer_1_compressor42_6.D ;
  assign _0428_ = \multiplier_16x16bit_pipelined.layer_1_compressor42_6.AB & \multiplier_16x16bit_pipelined.layer_1_compressor42_6.CD ;
  assign _0429_ = \multiplier_16x16bit_pipelined.layer_1_compressor42_6.AxorB & \multiplier_16x16bit_pipelined.layer_1_compressor42_6.CxorD ;
  assign _0430_ = \multiplier_16x16bit_pipelined.layer_1_compressor42_6.AxBxCxD & \multiplier_16x16bit_pipelined.layer_1_compressor42_6.cin ;
  assign \multiplier_16x16bit_pipelined.layer_1_compressor42_6.cout = \multiplier_16x16bit_pipelined.layer_1_compressor42_6.AB | \multiplier_16x16bit_pipelined.layer_1_compressor42_6.CD ;
  assign _0431_ = _0428_ | _0429_;
  assign \multiplier_16x16bit_pipelined.layer_1_compressor42_6.carry = _0431_ | _0430_;
  assign \multiplier_16x16bit_pipelined.layer_1_compressor42_6.AxorB = \multiplier_16x16bit_pipelined.layer_1_compressor42_6.A ^ \multiplier_16x16bit_pipelined.layer_1_compressor42_6.B ;
  assign \multiplier_16x16bit_pipelined.layer_1_compressor42_6.CxorD = \multiplier_16x16bit_pipelined.layer_1_compressor42_6.C ^ \multiplier_16x16bit_pipelined.layer_1_compressor42_6.D ;
  assign \multiplier_16x16bit_pipelined.layer_1_compressor42_6.AxBxCxD = \multiplier_16x16bit_pipelined.layer_1_compressor42_6.AxorB ^ \multiplier_16x16bit_pipelined.layer_1_compressor42_6.CxorD ;
  assign \multiplier_16x16bit_pipelined.layer_1_compressor42_6.S = \multiplier_16x16bit_pipelined.layer_1_compressor42_6.AxBxCxD ^ \multiplier_16x16bit_pipelined.layer_1_compressor42_6.cin ;
  assign \multiplier_16x16bit_pipelined.layer_1_compressor42_7.AB = \multiplier_16x16bit_pipelined.layer_1_compressor42_7.A & \multiplier_16x16bit_pipelined.layer_1_compressor42_7.B ;
  assign \multiplier_16x16bit_pipelined.layer_1_compressor42_7.CD = \multiplier_16x16bit_pipelined.layer_1_compressor42_7.C & \multiplier_16x16bit_pipelined.layer_1_compressor42_7.D ;
  assign _0432_ = \multiplier_16x16bit_pipelined.layer_1_compressor42_7.AB & \multiplier_16x16bit_pipelined.layer_1_compressor42_7.CD ;
  assign _0433_ = \multiplier_16x16bit_pipelined.layer_1_compressor42_7.AxorB & \multiplier_16x16bit_pipelined.layer_1_compressor42_7.CxorD ;
  assign _0434_ = \multiplier_16x16bit_pipelined.layer_1_compressor42_7.AxBxCxD & \multiplier_16x16bit_pipelined.layer_1_compressor42_7.cin ;
  assign \multiplier_16x16bit_pipelined.layer_1_compressor42_7.cout = \multiplier_16x16bit_pipelined.layer_1_compressor42_7.AB | \multiplier_16x16bit_pipelined.layer_1_compressor42_7.CD ;
  assign _0435_ = _0432_ | _0433_;
  assign \multiplier_16x16bit_pipelined.layer_1_compressor42_7.carry = _0435_ | _0434_;
  assign \multiplier_16x16bit_pipelined.layer_1_compressor42_7.AxorB = \multiplier_16x16bit_pipelined.layer_1_compressor42_7.A ^ \multiplier_16x16bit_pipelined.layer_1_compressor42_7.B ;
  assign \multiplier_16x16bit_pipelined.layer_1_compressor42_7.CxorD = \multiplier_16x16bit_pipelined.layer_1_compressor42_7.C ^ \multiplier_16x16bit_pipelined.layer_1_compressor42_7.D ;
  assign \multiplier_16x16bit_pipelined.layer_1_compressor42_7.AxBxCxD = \multiplier_16x16bit_pipelined.layer_1_compressor42_7.AxorB ^ \multiplier_16x16bit_pipelined.layer_1_compressor42_7.CxorD ;
  assign \multiplier_16x16bit_pipelined.layer_1_compressor42_7.S = \multiplier_16x16bit_pipelined.layer_1_compressor42_7.AxBxCxD ^ \multiplier_16x16bit_pipelined.layer_1_compressor42_7.cin ;
  assign \multiplier_16x16bit_pipelined.layer_1_compressor42_8.AB = \multiplier_16x16bit_pipelined.layer_1_compressor42_8.A & \multiplier_16x16bit_pipelined.layer_1_compressor42_8.B ;
  assign \multiplier_16x16bit_pipelined.layer_1_compressor42_8.CD = \multiplier_16x16bit_pipelined.layer_1_compressor42_8.C & \multiplier_16x16bit_pipelined.layer_1_compressor42_8.D ;
  assign _0436_ = \multiplier_16x16bit_pipelined.layer_1_compressor42_8.AB & \multiplier_16x16bit_pipelined.layer_1_compressor42_8.CD ;
  assign _0437_ = \multiplier_16x16bit_pipelined.layer_1_compressor42_8.AxorB & \multiplier_16x16bit_pipelined.layer_1_compressor42_8.CxorD ;
  assign _0438_ = \multiplier_16x16bit_pipelined.layer_1_compressor42_8.AxBxCxD & \multiplier_16x16bit_pipelined.layer_1_compressor42_8.cin ;
  assign \multiplier_16x16bit_pipelined.layer_1_compressor42_8.cout = \multiplier_16x16bit_pipelined.layer_1_compressor42_8.AB | \multiplier_16x16bit_pipelined.layer_1_compressor42_8.CD ;
  assign _0439_ = _0436_ | _0437_;
  assign \multiplier_16x16bit_pipelined.layer_1_compressor42_8.carry = _0439_ | _0438_;
  assign \multiplier_16x16bit_pipelined.layer_1_compressor42_8.AxorB = \multiplier_16x16bit_pipelined.layer_1_compressor42_8.A ^ \multiplier_16x16bit_pipelined.layer_1_compressor42_8.B ;
  assign \multiplier_16x16bit_pipelined.layer_1_compressor42_8.CxorD = \multiplier_16x16bit_pipelined.layer_1_compressor42_8.C ^ \multiplier_16x16bit_pipelined.layer_1_compressor42_8.D ;
  assign \multiplier_16x16bit_pipelined.layer_1_compressor42_8.AxBxCxD = \multiplier_16x16bit_pipelined.layer_1_compressor42_8.AxorB ^ \multiplier_16x16bit_pipelined.layer_1_compressor42_8.CxorD ;
  assign \multiplier_16x16bit_pipelined.layer_1_compressor42_8.S = \multiplier_16x16bit_pipelined.layer_1_compressor42_8.AxBxCxD ^ \multiplier_16x16bit_pipelined.layer_1_compressor42_8.cin ;
  assign \multiplier_16x16bit_pipelined.layer_1_compressor42_9.AB = \multiplier_16x16bit_pipelined.layer_1_compressor42_9.A & \multiplier_16x16bit_pipelined.layer_1_compressor42_9.B ;
  assign \multiplier_16x16bit_pipelined.layer_1_compressor42_9.CD = \multiplier_16x16bit_pipelined.layer_1_compressor42_9.C & \multiplier_16x16bit_pipelined.layer_1_compressor42_9.D ;
  assign _0440_ = \multiplier_16x16bit_pipelined.layer_1_compressor42_9.AB & \multiplier_16x16bit_pipelined.layer_1_compressor42_9.CD ;
  assign _0441_ = \multiplier_16x16bit_pipelined.layer_1_compressor42_9.AxorB & \multiplier_16x16bit_pipelined.layer_1_compressor42_9.CxorD ;
  assign _0442_ = \multiplier_16x16bit_pipelined.layer_1_compressor42_9.AxBxCxD & \multiplier_16x16bit_pipelined.layer_1_compressor42_9.cin ;
  assign \multiplier_16x16bit_pipelined.layer_1_compressor42_9.cout = \multiplier_16x16bit_pipelined.layer_1_compressor42_9.AB | \multiplier_16x16bit_pipelined.layer_1_compressor42_9.CD ;
  assign _0443_ = _0440_ | _0441_;
  assign \multiplier_16x16bit_pipelined.layer_1_compressor42_9.carry = _0443_ | _0442_;
  assign \multiplier_16x16bit_pipelined.layer_1_compressor42_9.AxorB = \multiplier_16x16bit_pipelined.layer_1_compressor42_9.A ^ \multiplier_16x16bit_pipelined.layer_1_compressor42_9.B ;
  assign \multiplier_16x16bit_pipelined.layer_1_compressor42_9.CxorD = \multiplier_16x16bit_pipelined.layer_1_compressor42_9.C ^ \multiplier_16x16bit_pipelined.layer_1_compressor42_9.D ;
  assign \multiplier_16x16bit_pipelined.layer_1_compressor42_9.AxBxCxD = \multiplier_16x16bit_pipelined.layer_1_compressor42_9.AxorB ^ \multiplier_16x16bit_pipelined.layer_1_compressor42_9.CxorD ;
  assign \multiplier_16x16bit_pipelined.layer_1_compressor42_9.S = \multiplier_16x16bit_pipelined.layer_1_compressor42_9.AxBxCxD ^ \multiplier_16x16bit_pipelined.layer_1_compressor42_9.cin ;
  assign \multiplier_16x16bit_pipelined.layer_1_full_adder_0.AB = \multiplier_16x16bit_pipelined.layer_1_full_adder_0.A & \multiplier_16x16bit_pipelined.layer_1_full_adder_0.B ;
  assign _0444_ = \multiplier_16x16bit_pipelined.layer_1_full_adder_0.AxorB & \multiplier_16x16bit_pipelined.layer_1_full_adder_0.cin ;
  assign \multiplier_16x16bit_pipelined.layer_1_full_adder_0.cout = \multiplier_16x16bit_pipelined.layer_1_full_adder_0.AB | _0444_;
  assign \multiplier_16x16bit_pipelined.layer_1_full_adder_0.AxorB = \multiplier_16x16bit_pipelined.layer_1_full_adder_0.A ^ \multiplier_16x16bit_pipelined.layer_1_full_adder_0.B ;
  assign \multiplier_16x16bit_pipelined.layer_1_full_adder_0.S = \multiplier_16x16bit_pipelined.layer_1_full_adder_0.AxorB ^ \multiplier_16x16bit_pipelined.layer_1_full_adder_0.cin ;
  assign \multiplier_16x16bit_pipelined.layer_1_full_adder_1.AB = \multiplier_16x16bit_pipelined.layer_1_full_adder_1.A & \multiplier_16x16bit_pipelined.layer_1_full_adder_1.B ;
  assign _0445_ = \multiplier_16x16bit_pipelined.layer_1_full_adder_1.AxorB & \multiplier_16x16bit_pipelined.layer_1_full_adder_1.cin ;
  assign \multiplier_16x16bit_pipelined.layer_1_full_adder_1.cout = \multiplier_16x16bit_pipelined.layer_1_full_adder_1.AB | _0445_;
  assign \multiplier_16x16bit_pipelined.layer_1_full_adder_1.AxorB = \multiplier_16x16bit_pipelined.layer_1_full_adder_1.A ^ \multiplier_16x16bit_pipelined.layer_1_full_adder_1.B ;
  assign \multiplier_16x16bit_pipelined.layer_1_full_adder_1.S = \multiplier_16x16bit_pipelined.layer_1_full_adder_1.AxorB ^ \multiplier_16x16bit_pipelined.layer_1_full_adder_1.cin ;
  assign \multiplier_16x16bit_pipelined.layer_1_full_adder_10.AB = \multiplier_16x16bit_pipelined.layer_1_full_adder_10.A & \multiplier_16x16bit_pipelined.layer_1_full_adder_10.B ;
  assign _0446_ = \multiplier_16x16bit_pipelined.layer_1_full_adder_10.AxorB & \multiplier_16x16bit_pipelined.layer_1_full_adder_10.cin ;
  assign \multiplier_16x16bit_pipelined.layer_1_full_adder_10.cout = \multiplier_16x16bit_pipelined.layer_1_full_adder_10.AB | _0446_;
  assign \multiplier_16x16bit_pipelined.layer_1_full_adder_10.AxorB = \multiplier_16x16bit_pipelined.layer_1_full_adder_10.A ^ \multiplier_16x16bit_pipelined.layer_1_full_adder_10.B ;
  assign \multiplier_16x16bit_pipelined.layer_1_full_adder_10.S = \multiplier_16x16bit_pipelined.layer_1_full_adder_10.AxorB ^ \multiplier_16x16bit_pipelined.layer_1_full_adder_10.cin ;
  assign \multiplier_16x16bit_pipelined.layer_1_full_adder_11.AB = \multiplier_16x16bit_pipelined.layer_1_full_adder_11.A & \multiplier_16x16bit_pipelined.layer_1_full_adder_11.B ;
  assign \multiplier_16x16bit_pipelined.layer_1_full_adder_11.cout = \multiplier_16x16bit_pipelined.layer_1_full_adder_11.AB | \multiplier_16x16bit_pipelined.layer_1_full_adder_11.AxorB ;
  assign \multiplier_16x16bit_pipelined.layer_1_full_adder_11.AxorB = \multiplier_16x16bit_pipelined.layer_1_full_adder_11.A ^ \multiplier_16x16bit_pipelined.layer_1_full_adder_11.B ;
  assign \multiplier_16x16bit_pipelined.layer_1_full_adder_11.S = \multiplier_16x16bit_pipelined.layer_1_full_adder_11.AxorB ^ 1'b1;
  assign \multiplier_16x16bit_pipelined.layer_1_full_adder_2.AB = \multiplier_16x16bit_pipelined.layer_1_full_adder_2.A & \multiplier_16x16bit_pipelined.layer_1_full_adder_2.B ;
  assign _0447_ = \multiplier_16x16bit_pipelined.layer_1_full_adder_2.AxorB & \multiplier_16x16bit_pipelined.layer_1_full_adder_2.cin ;
  assign \multiplier_16x16bit_pipelined.layer_1_full_adder_2.cout = \multiplier_16x16bit_pipelined.layer_1_full_adder_2.AB | _0447_;
  assign \multiplier_16x16bit_pipelined.layer_1_full_adder_2.AxorB = \multiplier_16x16bit_pipelined.layer_1_full_adder_2.A ^ \multiplier_16x16bit_pipelined.layer_1_full_adder_2.B ;
  assign \multiplier_16x16bit_pipelined.layer_1_full_adder_2.S = \multiplier_16x16bit_pipelined.layer_1_full_adder_2.AxorB ^ \multiplier_16x16bit_pipelined.layer_1_full_adder_2.cin ;
  assign \multiplier_16x16bit_pipelined.layer_1_full_adder_3.AB = \multiplier_16x16bit_pipelined.layer_1_full_adder_3.A & \multiplier_16x16bit_pipelined.layer_1_full_adder_3.B ;
  assign _0448_ = \multiplier_16x16bit_pipelined.layer_1_full_adder_3.AxorB & \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_6.negation ;
  assign \multiplier_16x16bit_pipelined.layer_1_full_adder_3.cout = \multiplier_16x16bit_pipelined.layer_1_full_adder_3.AB | _0448_;
  assign \multiplier_16x16bit_pipelined.layer_1_full_adder_3.AxorB = \multiplier_16x16bit_pipelined.layer_1_full_adder_3.A ^ \multiplier_16x16bit_pipelined.layer_1_full_adder_3.B ;
  assign \multiplier_16x16bit_pipelined.layer_1_full_adder_3.S = \multiplier_16x16bit_pipelined.layer_1_full_adder_3.AxorB ^ \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_6.negation ;
  assign \multiplier_16x16bit_pipelined.layer_1_full_adder_4.AB = \multiplier_16x16bit_pipelined.layer_1_full_adder_4.A & \multiplier_16x16bit_pipelined.layer_1_full_adder_4.B ;
  assign _0449_ = \multiplier_16x16bit_pipelined.layer_1_full_adder_4.AxorB & \multiplier_16x16bit_pipelined.layer_1_full_adder_4.cin ;
  assign \multiplier_16x16bit_pipelined.layer_1_full_adder_4.cout = \multiplier_16x16bit_pipelined.layer_1_full_adder_4.AB | _0449_;
  assign \multiplier_16x16bit_pipelined.layer_1_full_adder_4.AxorB = \multiplier_16x16bit_pipelined.layer_1_full_adder_4.A ^ \multiplier_16x16bit_pipelined.layer_1_full_adder_4.B ;
  assign \multiplier_16x16bit_pipelined.layer_1_full_adder_4.S = \multiplier_16x16bit_pipelined.layer_1_full_adder_4.AxorB ^ \multiplier_16x16bit_pipelined.layer_1_full_adder_4.cin ;
  assign \multiplier_16x16bit_pipelined.layer_1_full_adder_5.AB = \multiplier_16x16bit_pipelined.layer_1_full_adder_5.A & \multiplier_16x16bit_pipelined.layer_1_full_adder_5.B ;
  assign _0450_ = \multiplier_16x16bit_pipelined.layer_1_full_adder_5.AxorB & \multiplier_16x16bit_pipelined.layer_1_full_adder_5.cin ;
  assign \multiplier_16x16bit_pipelined.layer_1_full_adder_5.cout = \multiplier_16x16bit_pipelined.layer_1_full_adder_5.AB | _0450_;
  assign \multiplier_16x16bit_pipelined.layer_1_full_adder_5.AxorB = \multiplier_16x16bit_pipelined.layer_1_full_adder_5.A ^ \multiplier_16x16bit_pipelined.layer_1_full_adder_5.B ;
  assign \multiplier_16x16bit_pipelined.layer_1_full_adder_5.S = \multiplier_16x16bit_pipelined.layer_1_full_adder_5.AxorB ^ \multiplier_16x16bit_pipelined.layer_1_full_adder_5.cin ;
  assign \multiplier_16x16bit_pipelined.layer_1_full_adder_6.AB = \multiplier_16x16bit_pipelined.layer_1_full_adder_6.A & \multiplier_16x16bit_pipelined.layer_1_full_adder_6.B ;
  assign _0451_ = \multiplier_16x16bit_pipelined.layer_1_full_adder_6.AxorB & \multiplier_16x16bit_pipelined.layer_1_full_adder_6.cin ;
  assign \multiplier_16x16bit_pipelined.layer_1_full_adder_6.cout = \multiplier_16x16bit_pipelined.layer_1_full_adder_6.AB | _0451_;
  assign \multiplier_16x16bit_pipelined.layer_1_full_adder_6.AxorB = \multiplier_16x16bit_pipelined.layer_1_full_adder_6.A ^ \multiplier_16x16bit_pipelined.layer_1_full_adder_6.B ;
  assign \multiplier_16x16bit_pipelined.layer_1_full_adder_6.S = \multiplier_16x16bit_pipelined.layer_1_full_adder_6.AxorB ^ \multiplier_16x16bit_pipelined.layer_1_full_adder_6.cin ;
  assign \multiplier_16x16bit_pipelined.layer_1_full_adder_7.AB = \multiplier_16x16bit_pipelined.layer_1_full_adder_7.A & \multiplier_16x16bit_pipelined.layer_1_full_adder_7.B ;
  assign \multiplier_16x16bit_pipelined.layer_1_full_adder_7.cout = \multiplier_16x16bit_pipelined.layer_1_full_adder_7.AB | \multiplier_16x16bit_pipelined.layer_1_full_adder_7.AxorB ;
  assign \multiplier_16x16bit_pipelined.layer_1_full_adder_7.AxorB = \multiplier_16x16bit_pipelined.layer_1_full_adder_7.A ^ \multiplier_16x16bit_pipelined.layer_1_full_adder_7.B ;
  assign \multiplier_16x16bit_pipelined.layer_1_full_adder_7.S = \multiplier_16x16bit_pipelined.layer_1_full_adder_7.AxorB ^ 1'b1;
  assign \multiplier_16x16bit_pipelined.layer_1_full_adder_8.AB = \multiplier_16x16bit_pipelined.layer_1_full_adder_8.A & \multiplier_16x16bit_pipelined.layer_1_full_adder_8.B ;
  assign _0452_ = \multiplier_16x16bit_pipelined.layer_1_full_adder_8.AxorB & \multiplier_16x16bit_pipelined.layer_1_full_adder_8.cin ;
  assign \multiplier_16x16bit_pipelined.layer_1_full_adder_8.cout = \multiplier_16x16bit_pipelined.layer_1_full_adder_8.AB | _0452_;
  assign \multiplier_16x16bit_pipelined.layer_1_full_adder_8.AxorB = \multiplier_16x16bit_pipelined.layer_1_full_adder_8.A ^ \multiplier_16x16bit_pipelined.layer_1_full_adder_8.B ;
  assign \multiplier_16x16bit_pipelined.layer_1_full_adder_8.S = \multiplier_16x16bit_pipelined.layer_1_full_adder_8.AxorB ^ \multiplier_16x16bit_pipelined.layer_1_full_adder_8.cin ;
  assign \multiplier_16x16bit_pipelined.layer_1_full_adder_9.AB = \multiplier_16x16bit_pipelined.layer_1_full_adder_9.A & \multiplier_16x16bit_pipelined.layer_1_full_adder_9.B ;
  assign _0453_ = \multiplier_16x16bit_pipelined.layer_1_full_adder_9.AxorB & \multiplier_16x16bit_pipelined.layer_1_full_adder_9.cin ;
  assign \multiplier_16x16bit_pipelined.layer_1_full_adder_9.cout = \multiplier_16x16bit_pipelined.layer_1_full_adder_9.AB | _0453_;
  assign \multiplier_16x16bit_pipelined.layer_1_full_adder_9.AxorB = \multiplier_16x16bit_pipelined.layer_1_full_adder_9.A ^ \multiplier_16x16bit_pipelined.layer_1_full_adder_9.B ;
  assign \multiplier_16x16bit_pipelined.layer_1_full_adder_9.S = \multiplier_16x16bit_pipelined.layer_1_full_adder_9.AxorB ^ \multiplier_16x16bit_pipelined.layer_1_full_adder_9.cin ;
  assign \multiplier_16x16bit_pipelined.layer_2_compressor42_0.AB = \multiplier_16x16bit_pipelined.layer_1_compressor42_2.carry & \multiplier_16x16bit_pipelined.layer_1_compressor42_2.cout ;
  assign \multiplier_16x16bit_pipelined.layer_2_compressor42_0.CD = \multiplier_16x16bit_pipelined.layer_1_compressor42_3.S & \multiplier_16x16bit_pipelined.layer_2_compressor42_0.D ;
  assign _0454_ = \multiplier_16x16bit_pipelined.layer_2_compressor42_0.AB & \multiplier_16x16bit_pipelined.layer_2_compressor42_0.CD ;
  assign _0455_ = \multiplier_16x16bit_pipelined.layer_2_compressor42_0.AxorB & \multiplier_16x16bit_pipelined.layer_2_compressor42_0.CxorD ;
  assign _0456_ = \multiplier_16x16bit_pipelined.layer_2_compressor42_0.AxBxCxD & \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_5.negation ;
  assign \multiplier_16x16bit_pipelined.layer_2_compressor42_0.cout = \multiplier_16x16bit_pipelined.layer_2_compressor42_0.AB | \multiplier_16x16bit_pipelined.layer_2_compressor42_0.CD ;
  assign _0457_ = _0454_ | _0455_;
  assign \multiplier_16x16bit_pipelined.layer_2_compressor42_0.carry = _0457_ | _0456_;
  assign \multiplier_16x16bit_pipelined.layer_2_compressor42_0.AxorB = \multiplier_16x16bit_pipelined.layer_1_compressor42_2.carry ^ \multiplier_16x16bit_pipelined.layer_1_compressor42_2.cout ;
  assign \multiplier_16x16bit_pipelined.layer_2_compressor42_0.CxorD = \multiplier_16x16bit_pipelined.layer_1_compressor42_3.S ^ \multiplier_16x16bit_pipelined.layer_2_compressor42_0.D ;
  assign \multiplier_16x16bit_pipelined.layer_2_compressor42_0.AxBxCxD = \multiplier_16x16bit_pipelined.layer_2_compressor42_0.AxorB ^ \multiplier_16x16bit_pipelined.layer_2_compressor42_0.CxorD ;
  assign \multiplier_16x16bit_pipelined.layer_2_compressor42_0.S = \multiplier_16x16bit_pipelined.layer_2_compressor42_0.AxBxCxD ^ \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_5.negation ;
  assign \multiplier_16x16bit_pipelined.layer_2_compressor42_1.AB = \multiplier_16x16bit_pipelined.layer_1_compressor42_5.carry & \multiplier_16x16bit_pipelined.layer_1_compressor42_5.cout ;
  assign \multiplier_16x16bit_pipelined.layer_2_compressor42_1.CD = \multiplier_16x16bit_pipelined.layer_1_full_adder_3.cout & \multiplier_16x16bit_pipelined.layer_1_compressor42_6.S ;
  assign _0458_ = \multiplier_16x16bit_pipelined.layer_2_compressor42_1.AB & \multiplier_16x16bit_pipelined.layer_2_compressor42_1.CD ;
  assign _0459_ = \multiplier_16x16bit_pipelined.layer_2_compressor42_1.AxorB & \multiplier_16x16bit_pipelined.layer_2_compressor42_1.CxorD ;
  assign _0460_ = \multiplier_16x16bit_pipelined.layer_2_compressor42_1.AxBxCxD & \multiplier_16x16bit_pipelined.layer_2_compressor42_1.cin ;
  assign \multiplier_16x16bit_pipelined.layer_2_compressor42_1.cout = \multiplier_16x16bit_pipelined.layer_2_compressor42_1.AB | \multiplier_16x16bit_pipelined.layer_2_compressor42_1.CD ;
  assign _0461_ = _0458_ | _0459_;
  assign \multiplier_16x16bit_pipelined.layer_2_compressor42_1.carry = _0461_ | _0460_;
  assign \multiplier_16x16bit_pipelined.layer_2_compressor42_1.AxorB = \multiplier_16x16bit_pipelined.layer_1_compressor42_5.carry ^ \multiplier_16x16bit_pipelined.layer_1_compressor42_5.cout ;
  assign \multiplier_16x16bit_pipelined.layer_2_compressor42_1.CxorD = \multiplier_16x16bit_pipelined.layer_1_full_adder_3.cout ^ \multiplier_16x16bit_pipelined.layer_1_compressor42_6.S ;
  assign \multiplier_16x16bit_pipelined.layer_2_compressor42_1.AxBxCxD = \multiplier_16x16bit_pipelined.layer_2_compressor42_1.AxorB ^ \multiplier_16x16bit_pipelined.layer_2_compressor42_1.CxorD ;
  assign \multiplier_16x16bit_pipelined.layer_2_compressor42_1.S = \multiplier_16x16bit_pipelined.layer_2_compressor42_1.AxBxCxD ^ \multiplier_16x16bit_pipelined.layer_2_compressor42_1.cin ;
  assign \multiplier_16x16bit_pipelined.layer_2_compressor42_2.AB = \multiplier_16x16bit_pipelined.layer_1_compressor42_6.carry & \multiplier_16x16bit_pipelined.layer_1_compressor42_6.cout ;
  assign \multiplier_16x16bit_pipelined.layer_2_compressor42_2.CD = \multiplier_16x16bit_pipelined.layer_1_compressor42_7.S & \multiplier_16x16bit_pipelined.layer_1_full_adder_4.S ;
  assign _0462_ = \multiplier_16x16bit_pipelined.layer_2_compressor42_2.AB & \multiplier_16x16bit_pipelined.layer_2_compressor42_2.CD ;
  assign _0463_ = \multiplier_16x16bit_pipelined.layer_2_compressor42_2.AxorB & \multiplier_16x16bit_pipelined.layer_2_compressor42_2.CxorD ;
  assign _0464_ = \multiplier_16x16bit_pipelined.layer_2_compressor42_2.AxBxCxD & \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_7.negation ;
  assign \multiplier_16x16bit_pipelined.layer_2_compressor42_2.cout = \multiplier_16x16bit_pipelined.layer_2_compressor42_2.AB | \multiplier_16x16bit_pipelined.layer_2_compressor42_2.CD ;
  assign _0465_ = _0462_ | _0463_;
  assign \multiplier_16x16bit_pipelined.layer_2_compressor42_2.carry = _0465_ | _0464_;
  assign \multiplier_16x16bit_pipelined.layer_2_compressor42_2.AxorB = \multiplier_16x16bit_pipelined.layer_1_compressor42_6.carry ^ \multiplier_16x16bit_pipelined.layer_1_compressor42_6.cout ;
  assign \multiplier_16x16bit_pipelined.layer_2_compressor42_2.CxorD = \multiplier_16x16bit_pipelined.layer_1_compressor42_7.S ^ \multiplier_16x16bit_pipelined.layer_1_full_adder_4.S ;
  assign \multiplier_16x16bit_pipelined.layer_2_compressor42_2.AxBxCxD = \multiplier_16x16bit_pipelined.layer_2_compressor42_2.AxorB ^ \multiplier_16x16bit_pipelined.layer_2_compressor42_2.CxorD ;
  assign \multiplier_16x16bit_pipelined.layer_2_compressor42_2.S = \multiplier_16x16bit_pipelined.layer_2_compressor42_2.AxBxCxD ^ \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_7.negation ;
  assign \multiplier_16x16bit_pipelined.layer_2_compressor42_3.AB = \multiplier_16x16bit_pipelined.layer_1_compressor42_7.carry & \multiplier_16x16bit_pipelined.layer_1_compressor42_7.cout ;
  assign \multiplier_16x16bit_pipelined.layer_2_compressor42_3.CD = \multiplier_16x16bit_pipelined.layer_1_full_adder_4.cout & \multiplier_16x16bit_pipelined.layer_1_compressor42_8.S ;
  assign _0466_ = \multiplier_16x16bit_pipelined.layer_2_compressor42_3.AB & \multiplier_16x16bit_pipelined.layer_2_compressor42_3.CD ;
  assign _0467_ = \multiplier_16x16bit_pipelined.layer_2_compressor42_3.AxorB & \multiplier_16x16bit_pipelined.layer_2_compressor42_3.CxorD ;
  assign _0468_ = \multiplier_16x16bit_pipelined.layer_2_compressor42_3.AxBxCxD & \multiplier_16x16bit_pipelined.layer_1_full_adder_5.S ;
  assign \multiplier_16x16bit_pipelined.layer_2_compressor42_3.cout = \multiplier_16x16bit_pipelined.layer_2_compressor42_3.AB | \multiplier_16x16bit_pipelined.layer_2_compressor42_3.CD ;
  assign _0469_ = _0466_ | _0467_;
  assign \multiplier_16x16bit_pipelined.layer_2_compressor42_3.carry = _0469_ | _0468_;
  assign \multiplier_16x16bit_pipelined.layer_2_compressor42_3.AxorB = \multiplier_16x16bit_pipelined.layer_1_compressor42_7.carry ^ \multiplier_16x16bit_pipelined.layer_1_compressor42_7.cout ;
  assign \multiplier_16x16bit_pipelined.layer_2_compressor42_3.CxorD = \multiplier_16x16bit_pipelined.layer_1_full_adder_4.cout ^ \multiplier_16x16bit_pipelined.layer_1_compressor42_8.S ;
  assign \multiplier_16x16bit_pipelined.layer_2_compressor42_3.AxBxCxD = \multiplier_16x16bit_pipelined.layer_2_compressor42_3.AxorB ^ \multiplier_16x16bit_pipelined.layer_2_compressor42_3.CxorD ;
  assign \multiplier_16x16bit_pipelined.layer_2_compressor42_3.S = \multiplier_16x16bit_pipelined.layer_2_compressor42_3.AxBxCxD ^ \multiplier_16x16bit_pipelined.layer_1_full_adder_5.S ;
  assign \multiplier_16x16bit_pipelined.layer_2_compressor42_4.AB = \multiplier_16x16bit_pipelined.layer_1_compressor42_8.carry & \multiplier_16x16bit_pipelined.layer_1_compressor42_8.cout ;
  assign \multiplier_16x16bit_pipelined.layer_2_compressor42_4.CD = \multiplier_16x16bit_pipelined.layer_1_full_adder_5.cout & \multiplier_16x16bit_pipelined.layer_1_compressor42_9.S ;
  assign _0470_ = \multiplier_16x16bit_pipelined.layer_2_compressor42_4.AB & \multiplier_16x16bit_pipelined.layer_2_compressor42_4.CD ;
  assign _0471_ = \multiplier_16x16bit_pipelined.layer_2_compressor42_4.AxorB & \multiplier_16x16bit_pipelined.layer_2_compressor42_4.CxorD ;
  assign _0472_ = \multiplier_16x16bit_pipelined.layer_2_compressor42_4.AxBxCxD & \multiplier_16x16bit_pipelined.layer_1_full_adder_6.S ;
  assign \multiplier_16x16bit_pipelined.layer_2_compressor42_4.cout = \multiplier_16x16bit_pipelined.layer_2_compressor42_4.AB | \multiplier_16x16bit_pipelined.layer_2_compressor42_4.CD ;
  assign _0473_ = _0470_ | _0471_;
  assign \multiplier_16x16bit_pipelined.layer_2_compressor42_4.carry = _0473_ | _0472_;
  assign \multiplier_16x16bit_pipelined.layer_2_compressor42_4.AxorB = \multiplier_16x16bit_pipelined.layer_1_compressor42_8.carry ^ \multiplier_16x16bit_pipelined.layer_1_compressor42_8.cout ;
  assign \multiplier_16x16bit_pipelined.layer_2_compressor42_4.CxorD = \multiplier_16x16bit_pipelined.layer_1_full_adder_5.cout ^ \multiplier_16x16bit_pipelined.layer_1_compressor42_9.S ;
  assign \multiplier_16x16bit_pipelined.layer_2_compressor42_4.AxBxCxD = \multiplier_16x16bit_pipelined.layer_2_compressor42_4.AxorB ^ \multiplier_16x16bit_pipelined.layer_2_compressor42_4.CxorD ;
  assign \multiplier_16x16bit_pipelined.layer_2_compressor42_4.S = \multiplier_16x16bit_pipelined.layer_2_compressor42_4.AxBxCxD ^ \multiplier_16x16bit_pipelined.layer_1_full_adder_6.S ;
  assign \multiplier_16x16bit_pipelined.layer_2_compressor42_5.AB = \multiplier_16x16bit_pipelined.layer_1_compressor42_9.carry & \multiplier_16x16bit_pipelined.layer_1_compressor42_9.cout ;
  assign \multiplier_16x16bit_pipelined.layer_2_compressor42_5.CD = \multiplier_16x16bit_pipelined.layer_1_full_adder_6.cout & \multiplier_16x16bit_pipelined.layer_1_compressor42_10.S ;
  assign _0474_ = \multiplier_16x16bit_pipelined.layer_2_compressor42_5.AB & \multiplier_16x16bit_pipelined.layer_2_compressor42_5.CD ;
  assign _0475_ = \multiplier_16x16bit_pipelined.layer_2_compressor42_5.AxorB & \multiplier_16x16bit_pipelined.layer_2_compressor42_5.CxorD ;
  assign _0476_ = \multiplier_16x16bit_pipelined.layer_2_compressor42_5.AxBxCxD & \multiplier_16x16bit_pipelined.layer_1_full_adder_7.S ;
  assign \multiplier_16x16bit_pipelined.layer_2_compressor42_5.cout = \multiplier_16x16bit_pipelined.layer_2_compressor42_5.AB | \multiplier_16x16bit_pipelined.layer_2_compressor42_5.CD ;
  assign _0477_ = _0474_ | _0475_;
  assign \multiplier_16x16bit_pipelined.layer_2_compressor42_5.carry = _0477_ | _0476_;
  assign \multiplier_16x16bit_pipelined.layer_2_compressor42_5.AxorB = \multiplier_16x16bit_pipelined.layer_1_compressor42_9.carry ^ \multiplier_16x16bit_pipelined.layer_1_compressor42_9.cout ;
  assign \multiplier_16x16bit_pipelined.layer_2_compressor42_5.CxorD = \multiplier_16x16bit_pipelined.layer_1_full_adder_6.cout ^ \multiplier_16x16bit_pipelined.layer_1_compressor42_10.S ;
  assign \multiplier_16x16bit_pipelined.layer_2_compressor42_5.AxBxCxD = \multiplier_16x16bit_pipelined.layer_2_compressor42_5.AxorB ^ \multiplier_16x16bit_pipelined.layer_2_compressor42_5.CxorD ;
  assign \multiplier_16x16bit_pipelined.layer_2_compressor42_5.S = \multiplier_16x16bit_pipelined.layer_2_compressor42_5.AxBxCxD ^ \multiplier_16x16bit_pipelined.layer_1_full_adder_7.S ;
  assign \multiplier_16x16bit_pipelined.layer_2_compressor42_6.AB = \multiplier_16x16bit_pipelined.layer_1_compressor42_10.carry & \multiplier_16x16bit_pipelined.layer_1_compressor42_10.cout ;
  assign \multiplier_16x16bit_pipelined.layer_2_compressor42_6.CD = \multiplier_16x16bit_pipelined.layer_1_full_adder_7.cout & \multiplier_16x16bit_pipelined.layer_1_compressor42_11.S ;
  assign _0478_ = \multiplier_16x16bit_pipelined.layer_2_compressor42_6.AB & \multiplier_16x16bit_pipelined.layer_2_compressor42_6.CD ;
  assign _0479_ = \multiplier_16x16bit_pipelined.layer_2_compressor42_6.AxorB & \multiplier_16x16bit_pipelined.layer_2_compressor42_6.CxorD ;
  assign _0480_ = \multiplier_16x16bit_pipelined.layer_2_compressor42_6.AxBxCxD & \multiplier_16x16bit_pipelined.layer_2_compressor42_6.cin ;
  assign \multiplier_16x16bit_pipelined.layer_2_compressor42_6.cout = \multiplier_16x16bit_pipelined.layer_2_compressor42_6.AB | \multiplier_16x16bit_pipelined.layer_2_compressor42_6.CD ;
  assign _0481_ = _0478_ | _0479_;
  assign \multiplier_16x16bit_pipelined.layer_2_compressor42_6.carry = _0481_ | _0480_;
  assign \multiplier_16x16bit_pipelined.layer_2_compressor42_6.AxorB = \multiplier_16x16bit_pipelined.layer_1_compressor42_10.carry ^ \multiplier_16x16bit_pipelined.layer_1_compressor42_10.cout ;
  assign \multiplier_16x16bit_pipelined.layer_2_compressor42_6.CxorD = \multiplier_16x16bit_pipelined.layer_1_full_adder_7.cout ^ \multiplier_16x16bit_pipelined.layer_1_compressor42_11.S ;
  assign \multiplier_16x16bit_pipelined.layer_2_compressor42_6.AxBxCxD = \multiplier_16x16bit_pipelined.layer_2_compressor42_6.AxorB ^ \multiplier_16x16bit_pipelined.layer_2_compressor42_6.CxorD ;
  assign \multiplier_16x16bit_pipelined.layer_2_compressor42_6.S = \multiplier_16x16bit_pipelined.layer_2_compressor42_6.AxBxCxD ^ \multiplier_16x16bit_pipelined.layer_2_compressor42_6.cin ;
  assign \multiplier_16x16bit_pipelined.layer_2_compressor42_7.AB = \multiplier_16x16bit_pipelined.layer_1_compressor42_11.carry & \multiplier_16x16bit_pipelined.layer_1_compressor42_11.cout ;
  assign \multiplier_16x16bit_pipelined.layer_2_compressor42_7.CD = \multiplier_16x16bit_pipelined.layer_1_compressor42_12.S & \multiplier_16x16bit_pipelined.layer_2_compressor42_7.D ;
  assign _0482_ = \multiplier_16x16bit_pipelined.layer_2_compressor42_7.AB & \multiplier_16x16bit_pipelined.layer_2_compressor42_7.CD ;
  assign _0483_ = \multiplier_16x16bit_pipelined.layer_2_compressor42_7.AxorB & \multiplier_16x16bit_pipelined.layer_2_compressor42_7.CxorD ;
  assign \multiplier_16x16bit_pipelined.layer_2_compressor42_7.cout = \multiplier_16x16bit_pipelined.layer_2_compressor42_7.AB | \multiplier_16x16bit_pipelined.layer_2_compressor42_7.CD ;
  assign _0484_ = _0482_ | _0483_;
  assign \multiplier_16x16bit_pipelined.layer_2_compressor42_7.carry = _0484_ | \multiplier_16x16bit_pipelined.layer_2_compressor42_7.AxBxCxD ;
  assign \multiplier_16x16bit_pipelined.layer_2_compressor42_7.AxorB = \multiplier_16x16bit_pipelined.layer_1_compressor42_11.carry ^ \multiplier_16x16bit_pipelined.layer_1_compressor42_11.cout ;
  assign \multiplier_16x16bit_pipelined.layer_2_compressor42_7.CxorD = \multiplier_16x16bit_pipelined.layer_1_compressor42_12.S ^ \multiplier_16x16bit_pipelined.layer_2_compressor42_7.D ;
  assign \multiplier_16x16bit_pipelined.layer_2_compressor42_7.AxBxCxD = \multiplier_16x16bit_pipelined.layer_2_compressor42_7.AxorB ^ \multiplier_16x16bit_pipelined.layer_2_compressor42_7.CxorD ;
  assign \multiplier_16x16bit_pipelined.layer_2_compressor42_7.S = \multiplier_16x16bit_pipelined.layer_2_compressor42_7.AxBxCxD ^ 1'b1;
  assign \multiplier_16x16bit_pipelined.layer_2_full_adder_0.AB = \multiplier_16x16bit_pipelined.layer_1_compressor42_0.carry & \multiplier_16x16bit_pipelined.layer_1_compressor42_0.cout ;
  assign _0485_ = \multiplier_16x16bit_pipelined.layer_2_full_adder_0.AxorB & \multiplier_16x16bit_pipelined.layer_1_full_adder_2.S ;
  assign \multiplier_16x16bit_pipelined.layer_2_full_adder_0.cout = \multiplier_16x16bit_pipelined.layer_2_full_adder_0.AB | _0485_;
  assign \multiplier_16x16bit_pipelined.layer_2_full_adder_0.AxorB = \multiplier_16x16bit_pipelined.layer_1_compressor42_0.carry ^ \multiplier_16x16bit_pipelined.layer_1_compressor42_0.cout ;
  assign \multiplier_16x16bit_pipelined.layer_2_full_adder_0.S = \multiplier_16x16bit_pipelined.layer_2_full_adder_0.AxorB ^ \multiplier_16x16bit_pipelined.layer_1_full_adder_2.S ;
  assign \multiplier_16x16bit_pipelined.layer_2_full_adder_1.AB = \multiplier_16x16bit_pipelined.layer_1_full_adder_2.cout & \multiplier_16x16bit_pipelined.layer_1_compressor42_1.S ;
  assign _0486_ = \multiplier_16x16bit_pipelined.layer_2_full_adder_1.AxorB & \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_4.negation ;
  assign \multiplier_16x16bit_pipelined.layer_2_full_adder_1.cout = \multiplier_16x16bit_pipelined.layer_2_full_adder_1.AB | _0486_;
  assign \multiplier_16x16bit_pipelined.layer_2_full_adder_1.AxorB = \multiplier_16x16bit_pipelined.layer_1_full_adder_2.cout ^ \multiplier_16x16bit_pipelined.layer_1_compressor42_1.S ;
  assign \multiplier_16x16bit_pipelined.layer_2_full_adder_1.S = \multiplier_16x16bit_pipelined.layer_2_full_adder_1.AxorB ^ \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_4.negation ;
  assign \multiplier_16x16bit_pipelined.layer_2_full_adder_10.AB = \multiplier_16x16bit_pipelined.layer_1_full_adder_8.cout & \multiplier_16x16bit_pipelined.layer_1_full_adder_9.S ;
  assign \multiplier_16x16bit_pipelined.layer_2_full_adder_10.cout = \multiplier_16x16bit_pipelined.layer_2_full_adder_10.AB | \multiplier_16x16bit_pipelined.layer_2_full_adder_10.AxorB ;
  assign \multiplier_16x16bit_pipelined.layer_2_full_adder_10.AxorB = \multiplier_16x16bit_pipelined.layer_1_full_adder_8.cout ^ \multiplier_16x16bit_pipelined.layer_1_full_adder_9.S ;
  assign \multiplier_16x16bit_pipelined.layer_2_full_adder_10.S = \multiplier_16x16bit_pipelined.layer_2_full_adder_10.AxorB ^ 1'b1;
  assign \multiplier_16x16bit_pipelined.layer_2_full_adder_11.AB = \multiplier_16x16bit_pipelined.layer_1_full_adder_11.cout & \multiplier_16x16bit_pipelined.layer_2_full_adder_11.B ;
  assign _0487_ = \multiplier_16x16bit_pipelined.layer_2_full_adder_11.AxorB & \multiplier_16x16bit_pipelined.layer_2_full_adder_11.cin ;
  assign \multiplier_16x16bit_pipelined.layer_2_full_adder_11.cout = \multiplier_16x16bit_pipelined.layer_2_full_adder_11.AB | _0487_;
  assign \multiplier_16x16bit_pipelined.layer_2_full_adder_11.AxorB = \multiplier_16x16bit_pipelined.layer_1_full_adder_11.cout ^ \multiplier_16x16bit_pipelined.layer_2_full_adder_11.B ;
  assign \multiplier_16x16bit_pipelined.layer_2_full_adder_11.S = \multiplier_16x16bit_pipelined.layer_2_full_adder_11.AxorB ^ \multiplier_16x16bit_pipelined.layer_2_full_adder_11.cin ;
  assign \multiplier_16x16bit_pipelined.layer_2_full_adder_2.AB = \multiplier_16x16bit_pipelined.layer_1_compressor42_1.carry & \multiplier_16x16bit_pipelined.layer_1_compressor42_1.cout ;
  assign _0488_ = \multiplier_16x16bit_pipelined.layer_2_full_adder_2.AxorB & \multiplier_16x16bit_pipelined.layer_1_compressor42_2.S ;
  assign \multiplier_16x16bit_pipelined.layer_2_full_adder_2.cout = \multiplier_16x16bit_pipelined.layer_2_full_adder_2.AB | _0488_;
  assign \multiplier_16x16bit_pipelined.layer_2_full_adder_2.AxorB = \multiplier_16x16bit_pipelined.layer_1_compressor42_1.carry ^ \multiplier_16x16bit_pipelined.layer_1_compressor42_1.cout ;
  assign \multiplier_16x16bit_pipelined.layer_2_full_adder_2.S = \multiplier_16x16bit_pipelined.layer_2_full_adder_2.AxorB ^ \multiplier_16x16bit_pipelined.layer_1_compressor42_2.S ;
  assign \multiplier_16x16bit_pipelined.layer_2_full_adder_3.AB = \multiplier_16x16bit_pipelined.layer_1_compressor42_3.carry & \multiplier_16x16bit_pipelined.layer_1_compressor42_3.cout ;
  assign _0489_ = \multiplier_16x16bit_pipelined.layer_2_full_adder_3.AxorB & \multiplier_16x16bit_pipelined.layer_1_compressor42_4.S ;
  assign \multiplier_16x16bit_pipelined.layer_2_full_adder_3.cout = \multiplier_16x16bit_pipelined.layer_2_full_adder_3.AB | _0489_;
  assign \multiplier_16x16bit_pipelined.layer_2_full_adder_3.AxorB = \multiplier_16x16bit_pipelined.layer_1_compressor42_3.carry ^ \multiplier_16x16bit_pipelined.layer_1_compressor42_3.cout ;
  assign \multiplier_16x16bit_pipelined.layer_2_full_adder_3.S = \multiplier_16x16bit_pipelined.layer_2_full_adder_3.AxorB ^ \multiplier_16x16bit_pipelined.layer_1_compressor42_4.S ;
  assign \multiplier_16x16bit_pipelined.layer_2_full_adder_4.AB = \multiplier_16x16bit_pipelined.layer_1_compressor42_4.carry & \multiplier_16x16bit_pipelined.layer_1_compressor42_4.cout ;
  assign _0490_ = \multiplier_16x16bit_pipelined.layer_2_full_adder_4.AxorB & \multiplier_16x16bit_pipelined.layer_1_compressor42_5.S ;
  assign \multiplier_16x16bit_pipelined.layer_2_full_adder_4.cout = \multiplier_16x16bit_pipelined.layer_2_full_adder_4.AB | _0490_;
  assign \multiplier_16x16bit_pipelined.layer_2_full_adder_4.AxorB = \multiplier_16x16bit_pipelined.layer_1_compressor42_4.carry ^ \multiplier_16x16bit_pipelined.layer_1_compressor42_4.cout ;
  assign \multiplier_16x16bit_pipelined.layer_2_full_adder_4.S = \multiplier_16x16bit_pipelined.layer_2_full_adder_4.AxorB ^ \multiplier_16x16bit_pipelined.layer_1_compressor42_5.S ;
  assign \multiplier_16x16bit_pipelined.layer_2_full_adder_5.AB = \multiplier_16x16bit_pipelined.layer_1_compressor42_12.carry & \multiplier_16x16bit_pipelined.layer_1_compressor42_12.cout ;
  assign _0491_ = \multiplier_16x16bit_pipelined.layer_2_full_adder_5.AxorB & \multiplier_16x16bit_pipelined.layer_1_compressor42_13.S ;
  assign \multiplier_16x16bit_pipelined.layer_2_full_adder_5.cout = \multiplier_16x16bit_pipelined.layer_2_full_adder_5.AB | _0491_;
  assign \multiplier_16x16bit_pipelined.layer_2_full_adder_5.AxorB = \multiplier_16x16bit_pipelined.layer_1_compressor42_12.carry ^ \multiplier_16x16bit_pipelined.layer_1_compressor42_12.cout ;
  assign \multiplier_16x16bit_pipelined.layer_2_full_adder_5.S = \multiplier_16x16bit_pipelined.layer_2_full_adder_5.AxorB ^ \multiplier_16x16bit_pipelined.layer_1_compressor42_13.S ;
  assign \multiplier_16x16bit_pipelined.layer_2_full_adder_6.AB = \multiplier_16x16bit_pipelined.layer_1_compressor42_13.carry & \multiplier_16x16bit_pipelined.layer_1_compressor42_13.cout ;
  assign _0492_ = \multiplier_16x16bit_pipelined.layer_2_full_adder_6.AxorB & \multiplier_16x16bit_pipelined.layer_1_compressor42_14.S ;
  assign \multiplier_16x16bit_pipelined.layer_2_full_adder_6.cout = \multiplier_16x16bit_pipelined.layer_2_full_adder_6.AB | _0492_;
  assign \multiplier_16x16bit_pipelined.layer_2_full_adder_6.AxorB = \multiplier_16x16bit_pipelined.layer_1_compressor42_13.carry ^ \multiplier_16x16bit_pipelined.layer_1_compressor42_13.cout ;
  assign \multiplier_16x16bit_pipelined.layer_2_full_adder_6.S = \multiplier_16x16bit_pipelined.layer_2_full_adder_6.AxorB ^ \multiplier_16x16bit_pipelined.layer_1_compressor42_14.S ;
  assign \multiplier_16x16bit_pipelined.layer_2_full_adder_7.AB = \multiplier_16x16bit_pipelined.layer_1_compressor42_14.carry & \multiplier_16x16bit_pipelined.layer_1_compressor42_14.cout ;
  assign _0493_ = \multiplier_16x16bit_pipelined.layer_2_full_adder_7.AxorB & \multiplier_16x16bit_pipelined.layer_1_compressor42_15.S ;
  assign \multiplier_16x16bit_pipelined.layer_2_full_adder_7.cout = \multiplier_16x16bit_pipelined.layer_2_full_adder_7.AB | _0493_;
  assign \multiplier_16x16bit_pipelined.layer_2_full_adder_7.AxorB = \multiplier_16x16bit_pipelined.layer_1_compressor42_14.carry ^ \multiplier_16x16bit_pipelined.layer_1_compressor42_14.cout ;
  assign \multiplier_16x16bit_pipelined.layer_2_full_adder_7.S = \multiplier_16x16bit_pipelined.layer_2_full_adder_7.AxorB ^ \multiplier_16x16bit_pipelined.layer_1_compressor42_15.S ;
  assign \multiplier_16x16bit_pipelined.layer_2_full_adder_8.AB = \multiplier_16x16bit_pipelined.layer_1_compressor42_15.carry & \multiplier_16x16bit_pipelined.layer_1_compressor42_15.cout ;
  assign _0494_ = \multiplier_16x16bit_pipelined.layer_2_full_adder_8.AxorB & \multiplier_16x16bit_pipelined.layer_1_compressor42_16.S ;
  assign \multiplier_16x16bit_pipelined.layer_2_full_adder_8.cout = \multiplier_16x16bit_pipelined.layer_2_full_adder_8.AB | _0494_;
  assign \multiplier_16x16bit_pipelined.layer_2_full_adder_8.AxorB = \multiplier_16x16bit_pipelined.layer_1_compressor42_15.carry ^ \multiplier_16x16bit_pipelined.layer_1_compressor42_15.cout ;
  assign \multiplier_16x16bit_pipelined.layer_2_full_adder_8.S = \multiplier_16x16bit_pipelined.layer_2_full_adder_8.AxorB ^ \multiplier_16x16bit_pipelined.layer_1_compressor42_16.S ;
  assign \multiplier_16x16bit_pipelined.layer_2_full_adder_9.AB = \multiplier_16x16bit_pipelined.layer_1_compressor42_16.carry & \multiplier_16x16bit_pipelined.layer_1_compressor42_16.cout ;
  assign _0495_ = \multiplier_16x16bit_pipelined.layer_2_full_adder_9.AxorB & \multiplier_16x16bit_pipelined.layer_1_full_adder_8.S ;
  assign \multiplier_16x16bit_pipelined.layer_2_full_adder_9.cout = \multiplier_16x16bit_pipelined.layer_2_full_adder_9.AB | _0495_;
  assign \multiplier_16x16bit_pipelined.layer_2_full_adder_9.AxorB = \multiplier_16x16bit_pipelined.layer_1_compressor42_16.carry ^ \multiplier_16x16bit_pipelined.layer_1_compressor42_16.cout ;
  assign \multiplier_16x16bit_pipelined.layer_2_full_adder_9.S = \multiplier_16x16bit_pipelined.layer_2_full_adder_9.AxorB ^ \multiplier_16x16bit_pipelined.layer_1_full_adder_8.S ;
  assign \multiplier_16x16bit_pipelined.layer_3_full_adder_0.AB = \multiplier_16x16bit_pipelined.reg_layer_2_w11 [0] & \multiplier_16x16bit_pipelined.reg_layer_2_w11 [1];
  assign _0496_ = \multiplier_16x16bit_pipelined.layer_3_full_adder_0.AxorB & \multiplier_16x16bit_pipelined.reg_layer_2_w11 [2];
  assign \multiplier_16x16bit_pipelined.layer_3_full_adder_0.cout = \multiplier_16x16bit_pipelined.layer_3_full_adder_0.AB | _0496_;
  assign \multiplier_16x16bit_pipelined.layer_3_full_adder_0.AxorB = \multiplier_16x16bit_pipelined.reg_layer_2_w11 [0] ^ \multiplier_16x16bit_pipelined.reg_layer_2_w11 [1];
  assign \multiplier_16x16bit_pipelined.layer_3_full_adder_0.S = \multiplier_16x16bit_pipelined.layer_3_full_adder_0.AxorB ^ \multiplier_16x16bit_pipelined.reg_layer_2_w11 [2];
  assign \multiplier_16x16bit_pipelined.layer_3_full_adder_1.AB = \multiplier_16x16bit_pipelined.reg_layer_2_w12 [0] & \multiplier_16x16bit_pipelined.reg_layer_2_w12 [1];
  assign _0497_ = \multiplier_16x16bit_pipelined.layer_3_full_adder_1.AxorB & \multiplier_16x16bit_pipelined.reg_layer_2_w12 [2];
  assign \multiplier_16x16bit_pipelined.layer_3_full_adder_1.cout = \multiplier_16x16bit_pipelined.layer_3_full_adder_1.AB | _0497_;
  assign \multiplier_16x16bit_pipelined.layer_3_full_adder_1.AxorB = \multiplier_16x16bit_pipelined.reg_layer_2_w12 [0] ^ \multiplier_16x16bit_pipelined.reg_layer_2_w12 [1];
  assign \multiplier_16x16bit_pipelined.layer_3_full_adder_1.S = \multiplier_16x16bit_pipelined.layer_3_full_adder_1.AxorB ^ \multiplier_16x16bit_pipelined.reg_layer_2_w12 [2];
  assign \multiplier_16x16bit_pipelined.layer_3_full_adder_10.AB = \multiplier_16x16bit_pipelined.reg_layer_2_w21 [0] & \multiplier_16x16bit_pipelined.reg_layer_2_w21 [1];
  assign _0498_ = \multiplier_16x16bit_pipelined.layer_3_full_adder_10.AxorB & \multiplier_16x16bit_pipelined.reg_layer_2_w21 [2];
  assign \multiplier_16x16bit_pipelined.layer_3_full_adder_10.cout = \multiplier_16x16bit_pipelined.layer_3_full_adder_10.AB | _0498_;
  assign \multiplier_16x16bit_pipelined.layer_3_full_adder_10.AxorB = \multiplier_16x16bit_pipelined.reg_layer_2_w21 [0] ^ \multiplier_16x16bit_pipelined.reg_layer_2_w21 [1];
  assign \multiplier_16x16bit_pipelined.layer_3_full_adder_10.S = \multiplier_16x16bit_pipelined.layer_3_full_adder_10.AxorB ^ \multiplier_16x16bit_pipelined.reg_layer_2_w21 [2];
  assign \multiplier_16x16bit_pipelined.layer_3_full_adder_11.AB = \multiplier_16x16bit_pipelined.reg_layer_2_w24 [0] & \multiplier_16x16bit_pipelined.reg_layer_2_w24 [1];
  assign _0499_ = \multiplier_16x16bit_pipelined.layer_3_full_adder_11.AxorB & \multiplier_16x16bit_pipelined.reg_layer_2_w24 [2];
  assign \multiplier_16x16bit_pipelined.layer_3_full_adder_11.cout = \multiplier_16x16bit_pipelined.layer_3_full_adder_11.AB | _0499_;
  assign \multiplier_16x16bit_pipelined.layer_3_full_adder_11.AxorB = \multiplier_16x16bit_pipelined.reg_layer_2_w24 [0] ^ \multiplier_16x16bit_pipelined.reg_layer_2_w24 [1];
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_A_24.B = \multiplier_16x16bit_pipelined.layer_3_full_adder_11.AxorB ^ \multiplier_16x16bit_pipelined.reg_layer_2_w24 [2];
  assign \multiplier_16x16bit_pipelined.layer_3_full_adder_12.AB = \multiplier_16x16bit_pipelined.reg_layer_2_w26 [0] & \multiplier_16x16bit_pipelined.reg_layer_2_w26 [1];
  assign _0500_ = \multiplier_16x16bit_pipelined.layer_3_full_adder_12.AxorB & \multiplier_16x16bit_pipelined.reg_layer_2_w26 [2];
  assign \multiplier_16x16bit_pipelined.layer_3_full_adder_12.cout = \multiplier_16x16bit_pipelined.layer_3_full_adder_12.AB | _0500_;
  assign \multiplier_16x16bit_pipelined.layer_3_full_adder_12.AxorB = \multiplier_16x16bit_pipelined.reg_layer_2_w26 [0] ^ \multiplier_16x16bit_pipelined.reg_layer_2_w26 [1];
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_A_26.B = \multiplier_16x16bit_pipelined.layer_3_full_adder_12.AxorB ^ \multiplier_16x16bit_pipelined.reg_layer_2_w26 [2];
  assign \multiplier_16x16bit_pipelined.layer_3_full_adder_13.AB = \multiplier_16x16bit_pipelined.reg_layer_2_w29 [0] & \multiplier_16x16bit_pipelined.reg_layer_2_w29 [1];
  assign _0501_ = \multiplier_16x16bit_pipelined.layer_3_full_adder_13.AxorB & \multiplier_16x16bit_pipelined.reg_layer_2_w29 [2];
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_A_30.A = \multiplier_16x16bit_pipelined.layer_3_full_adder_13.AB | _0501_;
  assign \multiplier_16x16bit_pipelined.layer_3_full_adder_13.AxorB = \multiplier_16x16bit_pipelined.reg_layer_2_w29 [0] ^ \multiplier_16x16bit_pipelined.reg_layer_2_w29 [1];
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_A_29.A = \multiplier_16x16bit_pipelined.layer_3_full_adder_13.AxorB ^ \multiplier_16x16bit_pipelined.reg_layer_2_w29 [2];
  assign \multiplier_16x16bit_pipelined.layer_3_full_adder_2.AB = \multiplier_16x16bit_pipelined.reg_layer_2_w13 [0] & \multiplier_16x16bit_pipelined.reg_layer_2_w13 [1];
  assign _0502_ = \multiplier_16x16bit_pipelined.layer_3_full_adder_2.AxorB & \multiplier_16x16bit_pipelined.reg_layer_2_w13 [2];
  assign \multiplier_16x16bit_pipelined.layer_3_full_adder_2.cout = \multiplier_16x16bit_pipelined.layer_3_full_adder_2.AB | _0502_;
  assign \multiplier_16x16bit_pipelined.layer_3_full_adder_2.AxorB = \multiplier_16x16bit_pipelined.reg_layer_2_w13 [0] ^ \multiplier_16x16bit_pipelined.reg_layer_2_w13 [1];
  assign \multiplier_16x16bit_pipelined.layer_3_full_adder_2.S = \multiplier_16x16bit_pipelined.layer_3_full_adder_2.AxorB ^ \multiplier_16x16bit_pipelined.reg_layer_2_w13 [2];
  assign \multiplier_16x16bit_pipelined.layer_3_full_adder_3.AB = \multiplier_16x16bit_pipelined.reg_layer_2_w14 [0] & \multiplier_16x16bit_pipelined.reg_layer_2_w14 [1];
  assign _0503_ = \multiplier_16x16bit_pipelined.layer_3_full_adder_3.AxorB & \multiplier_16x16bit_pipelined.reg_layer_2_w14 [2];
  assign \multiplier_16x16bit_pipelined.layer_3_full_adder_3.cout = \multiplier_16x16bit_pipelined.layer_3_full_adder_3.AB | _0503_;
  assign \multiplier_16x16bit_pipelined.layer_3_full_adder_3.AxorB = \multiplier_16x16bit_pipelined.reg_layer_2_w14 [0] ^ \multiplier_16x16bit_pipelined.reg_layer_2_w14 [1];
  assign \multiplier_16x16bit_pipelined.layer_3_full_adder_3.S = \multiplier_16x16bit_pipelined.layer_3_full_adder_3.AxorB ^ \multiplier_16x16bit_pipelined.reg_layer_2_w14 [2];
  assign \multiplier_16x16bit_pipelined.layer_3_full_adder_4.AB = \multiplier_16x16bit_pipelined.reg_layer_2_w15 [0] & \multiplier_16x16bit_pipelined.reg_layer_2_w15 [1];
  assign _0504_ = \multiplier_16x16bit_pipelined.layer_3_full_adder_4.AxorB & \multiplier_16x16bit_pipelined.reg_layer_2_w15 [2];
  assign \multiplier_16x16bit_pipelined.layer_3_full_adder_4.cout = \multiplier_16x16bit_pipelined.layer_3_full_adder_4.AB | _0504_;
  assign \multiplier_16x16bit_pipelined.layer_3_full_adder_4.AxorB = \multiplier_16x16bit_pipelined.reg_layer_2_w15 [0] ^ \multiplier_16x16bit_pipelined.reg_layer_2_w15 [1];
  assign \multiplier_16x16bit_pipelined.layer_3_full_adder_4.S = \multiplier_16x16bit_pipelined.layer_3_full_adder_4.AxorB ^ \multiplier_16x16bit_pipelined.reg_layer_2_w15 [2];
  assign \multiplier_16x16bit_pipelined.layer_3_full_adder_5.AB = \multiplier_16x16bit_pipelined.reg_layer_2_w16 [0] & \multiplier_16x16bit_pipelined.reg_layer_2_w16 [1];
  assign _0505_ = \multiplier_16x16bit_pipelined.layer_3_full_adder_5.AxorB & \multiplier_16x16bit_pipelined.reg_layer_2_w16 [2];
  assign \multiplier_16x16bit_pipelined.layer_3_full_adder_5.cout = \multiplier_16x16bit_pipelined.layer_3_full_adder_5.AB | _0505_;
  assign \multiplier_16x16bit_pipelined.layer_3_full_adder_5.AxorB = \multiplier_16x16bit_pipelined.reg_layer_2_w16 [0] ^ \multiplier_16x16bit_pipelined.reg_layer_2_w16 [1];
  assign \multiplier_16x16bit_pipelined.layer_3_full_adder_5.S = \multiplier_16x16bit_pipelined.layer_3_full_adder_5.AxorB ^ \multiplier_16x16bit_pipelined.reg_layer_2_w16 [2];
  assign \multiplier_16x16bit_pipelined.layer_3_full_adder_6.AB = \multiplier_16x16bit_pipelined.reg_layer_2_w17 [0] & \multiplier_16x16bit_pipelined.reg_layer_2_w17 [1];
  assign _0506_ = \multiplier_16x16bit_pipelined.layer_3_full_adder_6.AxorB & \multiplier_16x16bit_pipelined.reg_layer_2_w17 [2];
  assign \multiplier_16x16bit_pipelined.layer_3_full_adder_6.cout = \multiplier_16x16bit_pipelined.layer_3_full_adder_6.AB | _0506_;
  assign \multiplier_16x16bit_pipelined.layer_3_full_adder_6.AxorB = \multiplier_16x16bit_pipelined.reg_layer_2_w17 [0] ^ \multiplier_16x16bit_pipelined.reg_layer_2_w17 [1];
  assign \multiplier_16x16bit_pipelined.layer_3_full_adder_6.S = \multiplier_16x16bit_pipelined.layer_3_full_adder_6.AxorB ^ \multiplier_16x16bit_pipelined.reg_layer_2_w17 [2];
  assign \multiplier_16x16bit_pipelined.layer_3_full_adder_7.AB = \multiplier_16x16bit_pipelined.reg_layer_2_w18 [0] & \multiplier_16x16bit_pipelined.reg_layer_2_w18 [1];
  assign _0507_ = \multiplier_16x16bit_pipelined.layer_3_full_adder_7.AxorB & \multiplier_16x16bit_pipelined.reg_layer_2_w18 [2];
  assign \multiplier_16x16bit_pipelined.layer_3_full_adder_7.cout = \multiplier_16x16bit_pipelined.layer_3_full_adder_7.AB | _0507_;
  assign \multiplier_16x16bit_pipelined.layer_3_full_adder_7.AxorB = \multiplier_16x16bit_pipelined.reg_layer_2_w18 [0] ^ \multiplier_16x16bit_pipelined.reg_layer_2_w18 [1];
  assign \multiplier_16x16bit_pipelined.layer_3_full_adder_7.S = \multiplier_16x16bit_pipelined.layer_3_full_adder_7.AxorB ^ \multiplier_16x16bit_pipelined.reg_layer_2_w18 [2];
  assign \multiplier_16x16bit_pipelined.layer_3_full_adder_8.AB = \multiplier_16x16bit_pipelined.reg_layer_2_w19 [0] & \multiplier_16x16bit_pipelined.reg_layer_2_w19 [1];
  assign _0508_ = \multiplier_16x16bit_pipelined.layer_3_full_adder_8.AxorB & \multiplier_16x16bit_pipelined.reg_layer_2_w19 [2];
  assign \multiplier_16x16bit_pipelined.layer_3_full_adder_8.cout = \multiplier_16x16bit_pipelined.layer_3_full_adder_8.AB | _0508_;
  assign \multiplier_16x16bit_pipelined.layer_3_full_adder_8.AxorB = \multiplier_16x16bit_pipelined.reg_layer_2_w19 [0] ^ \multiplier_16x16bit_pipelined.reg_layer_2_w19 [1];
  assign \multiplier_16x16bit_pipelined.layer_3_full_adder_8.S = \multiplier_16x16bit_pipelined.layer_3_full_adder_8.AxorB ^ \multiplier_16x16bit_pipelined.reg_layer_2_w19 [2];
  assign \multiplier_16x16bit_pipelined.layer_3_full_adder_9.AB = \multiplier_16x16bit_pipelined.reg_layer_2_w20 [0] & \multiplier_16x16bit_pipelined.reg_layer_2_w20 [1];
  assign _0509_ = \multiplier_16x16bit_pipelined.layer_3_full_adder_9.AxorB & \multiplier_16x16bit_pipelined.reg_layer_2_w20 [2];
  assign \multiplier_16x16bit_pipelined.layer_3_full_adder_9.cout = \multiplier_16x16bit_pipelined.layer_3_full_adder_9.AB | _0509_;
  assign \multiplier_16x16bit_pipelined.layer_3_full_adder_9.AxorB = \multiplier_16x16bit_pipelined.reg_layer_2_w20 [0] ^ \multiplier_16x16bit_pipelined.reg_layer_2_w20 [1];
  assign \multiplier_16x16bit_pipelined.layer_3_full_adder_9.S = \multiplier_16x16bit_pipelined.layer_3_full_adder_9.AxorB ^ \multiplier_16x16bit_pipelined.reg_layer_2_w20 [2];
  assign \multiplier_16x16bit_pipelined.layer_4_full_adder_0.AB = \multiplier_16x16bit_pipelined.reg_layer_2_w2 [0] & \multiplier_16x16bit_pipelined.reg_layer_2_w2 [1];
  assign _0510_ = \multiplier_16x16bit_pipelined.layer_4_full_adder_0.AxorB & \multiplier_16x16bit_pipelined.reg_layer_2_w2 [2];
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_A_3.A = \multiplier_16x16bit_pipelined.layer_4_full_adder_0.AB | _0510_;
  assign \multiplier_16x16bit_pipelined.layer_4_full_adder_0.AxorB = \multiplier_16x16bit_pipelined.reg_layer_2_w2 [0] ^ \multiplier_16x16bit_pipelined.reg_layer_2_w2 [1];
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_A_2.A = \multiplier_16x16bit_pipelined.layer_4_full_adder_0.AxorB ^ \multiplier_16x16bit_pipelined.reg_layer_2_w2 [2];
  assign \multiplier_16x16bit_pipelined.layer_4_full_adder_1.AB = \multiplier_16x16bit_pipelined.layer_3_full_adder_4.cout & \multiplier_16x16bit_pipelined.layer_3_full_adder_5.S ;
  assign _0511_ = \multiplier_16x16bit_pipelined.layer_4_full_adder_1.AxorB & \multiplier_16x16bit_pipelined.reg_layer_2_w16 [3];
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_A_17.A = \multiplier_16x16bit_pipelined.layer_4_full_adder_1.AB | _0511_;
  assign \multiplier_16x16bit_pipelined.layer_4_full_adder_1.AxorB = \multiplier_16x16bit_pipelined.layer_3_full_adder_4.cout ^ \multiplier_16x16bit_pipelined.layer_3_full_adder_5.S ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_A_16.B = \multiplier_16x16bit_pipelined.layer_4_full_adder_1.AxorB ^ \multiplier_16x16bit_pipelined.reg_layer_2_w16 [3];
  assign \multiplier_16x16bit_pipelined.layer_4_full_adder_2.AB = \multiplier_16x16bit_pipelined.layer_3_full_adder_6.cout & \multiplier_16x16bit_pipelined.layer_3_full_adder_7.S ;
  assign _0512_ = \multiplier_16x16bit_pipelined.layer_4_full_adder_2.AxorB & \multiplier_16x16bit_pipelined.reg_layer_2_w18 [3];
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_A_19.A = \multiplier_16x16bit_pipelined.layer_4_full_adder_2.AB | _0512_;
  assign \multiplier_16x16bit_pipelined.layer_4_full_adder_2.AxorB = \multiplier_16x16bit_pipelined.layer_3_full_adder_6.cout ^ \multiplier_16x16bit_pipelined.layer_3_full_adder_7.S ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_A_18.B = \multiplier_16x16bit_pipelined.layer_4_full_adder_2.AxorB ^ \multiplier_16x16bit_pipelined.reg_layer_2_w18 [3];
  assign \multiplier_16x16bit_pipelined.layer_4_full_adder_3.AB = \multiplier_16x16bit_pipelined.layer_3_full_adder_8.cout & \multiplier_16x16bit_pipelined.layer_3_full_adder_9.S ;
  assign _0513_ = \multiplier_16x16bit_pipelined.layer_4_full_adder_3.AxorB & \multiplier_16x16bit_pipelined.reg_layer_2_w20 [3];
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_A_21.A = \multiplier_16x16bit_pipelined.layer_4_full_adder_3.AB | _0513_;
  assign \multiplier_16x16bit_pipelined.layer_4_full_adder_3.AxorB = \multiplier_16x16bit_pipelined.layer_3_full_adder_8.cout ^ \multiplier_16x16bit_pipelined.layer_3_full_adder_9.S ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_A_20.B = \multiplier_16x16bit_pipelined.layer_4_full_adder_3.AxorB ^ \multiplier_16x16bit_pipelined.reg_layer_2_w20 [3];
  assign \multiplier_16x16bit_pipelined.layer_4_full_adder_4.AB = \multiplier_16x16bit_pipelined.layer_3_full_adder_10.cout & \multiplier_16x16bit_pipelined.reg_layer_2_w22 [0];
  assign _0514_ = \multiplier_16x16bit_pipelined.layer_4_full_adder_4.AxorB & \multiplier_16x16bit_pipelined.reg_layer_2_w22 [1];
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_A_23.A = \multiplier_16x16bit_pipelined.layer_4_full_adder_4.AB | _0514_;
  assign \multiplier_16x16bit_pipelined.layer_4_full_adder_4.AxorB = \multiplier_16x16bit_pipelined.layer_3_full_adder_10.cout ^ \multiplier_16x16bit_pipelined.reg_layer_2_w22 [0];
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_A_22.B = \multiplier_16x16bit_pipelined.layer_4_full_adder_4.AxorB ^ \multiplier_16x16bit_pipelined.reg_layer_2_w22 [1];
  assign \multiplier_16x16bit_pipelined.layer_4_full_adder_5.AB = \multiplier_16x16bit_pipelined.layer_3_full_adder_11.cout & \multiplier_16x16bit_pipelined.reg_layer_2_w25 [0];
  assign _0515_ = \multiplier_16x16bit_pipelined.layer_4_full_adder_5.AxorB & \multiplier_16x16bit_pipelined.reg_layer_2_w25 [1];
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_A_26.A = \multiplier_16x16bit_pipelined.layer_4_full_adder_5.AB | _0515_;
  assign \multiplier_16x16bit_pipelined.layer_4_full_adder_5.AxorB = \multiplier_16x16bit_pipelined.layer_3_full_adder_11.cout ^ \multiplier_16x16bit_pipelined.reg_layer_2_w25 [0];
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_A_25.A = \multiplier_16x16bit_pipelined.layer_4_full_adder_5.AxorB ^ \multiplier_16x16bit_pipelined.reg_layer_2_w25 [1];
  assign \multiplier_16x16bit_pipelined.layer_4_full_adder_6.AB = \multiplier_16x16bit_pipelined.layer_3_full_adder_12.cout & \multiplier_16x16bit_pipelined.reg_layer_2_w27 [0];
  assign _0516_ = \multiplier_16x16bit_pipelined.layer_4_full_adder_6.AxorB & \multiplier_16x16bit_pipelined.reg_layer_2_w27 [1];
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_A_28.A = \multiplier_16x16bit_pipelined.layer_4_full_adder_6.AB | _0516_;
  assign \multiplier_16x16bit_pipelined.layer_4_full_adder_6.AxorB = \multiplier_16x16bit_pipelined.layer_3_full_adder_12.cout ^ \multiplier_16x16bit_pipelined.reg_layer_2_w27 [0];
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_A_27.A = \multiplier_16x16bit_pipelined.layer_4_full_adder_6.AxorB ^ \multiplier_16x16bit_pipelined.reg_layer_2_w27 [1];
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_A_4.A = \multiplier_16x16bit_pipelined.reg_layer_2_w3 [0] & \multiplier_16x16bit_pipelined.reg_layer_2_w3 [1];
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_A_3.B = \multiplier_16x16bit_pipelined.reg_layer_2_w3 [0] ^ \multiplier_16x16bit_pipelined.reg_layer_2_w3 [1];
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_A_5.A = \multiplier_16x16bit_pipelined.reg_layer_2_w4 [0] & \multiplier_16x16bit_pipelined.reg_layer_2_w4 [1];
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_A_4.B = \multiplier_16x16bit_pipelined.reg_layer_2_w4 [0] ^ \multiplier_16x16bit_pipelined.reg_layer_2_w4 [1];
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_A_14.A = \multiplier_16x16bit_pipelined.layer_3_full_adder_1.cout & \multiplier_16x16bit_pipelined.layer_3_full_adder_2.S ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_A_13.B = \multiplier_16x16bit_pipelined.layer_3_full_adder_1.cout ^ \multiplier_16x16bit_pipelined.layer_3_full_adder_2.S ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_A_15.A = \multiplier_16x16bit_pipelined.layer_3_full_adder_2.cout & \multiplier_16x16bit_pipelined.layer_3_full_adder_3.S ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_A_14.B = \multiplier_16x16bit_pipelined.layer_3_full_adder_2.cout ^ \multiplier_16x16bit_pipelined.layer_3_full_adder_3.S ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_A_16.A = \multiplier_16x16bit_pipelined.layer_3_full_adder_3.cout & \multiplier_16x16bit_pipelined.layer_3_full_adder_4.S ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_A_15.B = \multiplier_16x16bit_pipelined.layer_3_full_adder_3.cout ^ \multiplier_16x16bit_pipelined.layer_3_full_adder_4.S ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_A_18.A = \multiplier_16x16bit_pipelined.layer_3_full_adder_5.cout & \multiplier_16x16bit_pipelined.layer_3_full_adder_6.S ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_A_17.B = \multiplier_16x16bit_pipelined.layer_3_full_adder_5.cout ^ \multiplier_16x16bit_pipelined.layer_3_full_adder_6.S ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_A_20.A = \multiplier_16x16bit_pipelined.layer_3_full_adder_7.cout & \multiplier_16x16bit_pipelined.layer_3_full_adder_8.S ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_A_19.B = \multiplier_16x16bit_pipelined.layer_3_full_adder_7.cout ^ \multiplier_16x16bit_pipelined.layer_3_full_adder_8.S ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_A_22.A = \multiplier_16x16bit_pipelined.layer_3_full_adder_9.cout & \multiplier_16x16bit_pipelined.layer_3_full_adder_10.S ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_A_21.B = \multiplier_16x16bit_pipelined.layer_3_full_adder_9.cout ^ \multiplier_16x16bit_pipelined.layer_3_full_adder_10.S ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_A_24.A = \multiplier_16x16bit_pipelined.reg_layer_2_w23 [0] & \multiplier_16x16bit_pipelined.reg_layer_2_w23 [1];
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_A_23.B = \multiplier_16x16bit_pipelined.reg_layer_2_w23 [0] ^ \multiplier_16x16bit_pipelined.reg_layer_2_w23 [1];
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_A_6.A = \multiplier_16x16bit_pipelined.reg_layer_2_w5 [0] & \multiplier_16x16bit_pipelined.reg_layer_2_w5 [1];
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_A_5.B = \multiplier_16x16bit_pipelined.reg_layer_2_w5 [0] ^ \multiplier_16x16bit_pipelined.reg_layer_2_w5 [1];
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_A_7.A = \multiplier_16x16bit_pipelined.reg_layer_2_w6 [0] & \multiplier_16x16bit_pipelined.reg_layer_2_w6 [1];
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_A_6.B = \multiplier_16x16bit_pipelined.reg_layer_2_w6 [0] ^ \multiplier_16x16bit_pipelined.reg_layer_2_w6 [1];
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_A_8.A = \multiplier_16x16bit_pipelined.reg_layer_2_w7 [0] & \multiplier_16x16bit_pipelined.reg_layer_2_w7 [1];
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_A_7.B = \multiplier_16x16bit_pipelined.reg_layer_2_w7 [0] ^ \multiplier_16x16bit_pipelined.reg_layer_2_w7 [1];
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_A_9.A = \multiplier_16x16bit_pipelined.reg_layer_2_w8 [0] & \multiplier_16x16bit_pipelined.reg_layer_2_w8 [1];
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_A_8.B = \multiplier_16x16bit_pipelined.reg_layer_2_w8 [0] ^ \multiplier_16x16bit_pipelined.reg_layer_2_w8 [1];
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_A_10.A = \multiplier_16x16bit_pipelined.reg_layer_2_w9 [0] & \multiplier_16x16bit_pipelined.reg_layer_2_w9 [1];
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_A_9.B = \multiplier_16x16bit_pipelined.reg_layer_2_w9 [0] ^ \multiplier_16x16bit_pipelined.reg_layer_2_w9 [1];
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_A_11.A = \multiplier_16x16bit_pipelined.reg_layer_2_w10 [0] & \multiplier_16x16bit_pipelined.reg_layer_2_w10 [1];
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_A_10.B = \multiplier_16x16bit_pipelined.reg_layer_2_w10 [0] ^ \multiplier_16x16bit_pipelined.reg_layer_2_w10 [1];
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_A_12.A = \multiplier_16x16bit_pipelined.layer_3_full_adder_0.S & \multiplier_16x16bit_pipelined.reg_layer_2_w11 [3];
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_A_11.B = \multiplier_16x16bit_pipelined.layer_3_full_adder_0.S ^ \multiplier_16x16bit_pipelined.reg_layer_2_w11 [3];
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_A_13.A = \multiplier_16x16bit_pipelined.layer_3_full_adder_0.cout & \multiplier_16x16bit_pipelined.layer_3_full_adder_1.S ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_A_12.B = \multiplier_16x16bit_pipelined.layer_3_full_adder_0.cout ^ \multiplier_16x16bit_pipelined.layer_3_full_adder_1.S ;
  assign _0517_ = ~ \multiplier_16x16bit_pipelined.md ;
  assign \multiplier_16x16bit_pipelined.layer_1_compressor42_9.A = ~ \multiplier_16x16bit_pipelined.partial_product_gen_0.zmd [15];
  assign \multiplier_16x16bit_pipelined.partial_product_gen_0.nmd = \multiplier_16x16bit_pipelined.mr [1] ? _0517_ : \multiplier_16x16bit_pipelined.md ;
  assign \multiplier_16x16bit_pipelined.partial_product_gen_0.zmd = \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_0.zero ? 16'b0000000000000000 : \multiplier_16x16bit_pipelined.partial_product_gen_0.nmd ;
  wire [15:0] fangyuan74;
  assign { \multiplier_16x16bit_pipelined.layer_1_compressor42_8.A , \multiplier_16x16bit_pipelined.layer_1_compressor42_7.A , \multiplier_16x16bit_pipelined.layer_1_compressor42_6.A , \multiplier_16x16bit_pipelined.layer_1_compressor42_5.A , \multiplier_16x16bit_pipelined.layer_1_compressor42_4.A , \multiplier_16x16bit_pipelined.layer_1_compressor42_3.A , \multiplier_16x16bit_pipelined.layer_1_compressor42_2.A , \multiplier_16x16bit_pipelined.layer_1_compressor42_1.A , \multiplier_16x16bit_pipelined.layer_1_full_adder_2.A , \multiplier_16x16bit_pipelined.layer_1_compressor42_0.A , \multiplier_16x16bit_pipelined.layer_1_full_adder_1.A , \multiplier_16x16bit_pipelined.layer_1_full_adder_0.A , \multiplier_16x16bit_pipelined.layer_0_w3[0] , \multiplier_16x16bit_pipelined.layer_0_w2[0] , \multiplier_16x16bit_pipelined.layer_0_w1 , \multiplier_16x16bit_pipelined.layer_0_w0[0] } = fangyuan74;
  wire [15:0] fangyuan75;
  assign fangyuan75 = { \multiplier_16x16bit_pipelined.partial_product_gen_0.zmd [14:0], \multiplier_16x16bit_pipelined.mr [1] };

  assign fangyuan74 = \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_0.double ? fangyuan75 : \multiplier_16x16bit_pipelined.partial_product_gen_0.zmd ;
  assign \multiplier_16x16bit_pipelined.layer_1_compressor42_11.A = ~ \multiplier_16x16bit_pipelined.partial_product_gen_1.zmd [15];
  assign \multiplier_16x16bit_pipelined.partial_product_gen_1.nmd = \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_1.negation ? _0517_ : \multiplier_16x16bit_pipelined.md ;
  assign \multiplier_16x16bit_pipelined.partial_product_gen_1.zmd = \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_1.zero ? 16'b0000000000000000 : \multiplier_16x16bit_pipelined.partial_product_gen_1.nmd ;
  wire [15:0] fangyuan76;
  assign { \multiplier_16x16bit_pipelined.layer_1_compressor42_10.A , \multiplier_16x16bit_pipelined.layer_1_compressor42_9.B , \multiplier_16x16bit_pipelined.layer_1_compressor42_8.B , \multiplier_16x16bit_pipelined.layer_1_compressor42_7.B , \multiplier_16x16bit_pipelined.layer_1_compressor42_6.B , \multiplier_16x16bit_pipelined.layer_1_compressor42_5.B , \multiplier_16x16bit_pipelined.layer_1_compressor42_4.B , \multiplier_16x16bit_pipelined.layer_1_compressor42_3.B , \multiplier_16x16bit_pipelined.layer_1_compressor42_2.B , \multiplier_16x16bit_pipelined.layer_1_compressor42_1.B , \multiplier_16x16bit_pipelined.layer_1_full_adder_2.B , \multiplier_16x16bit_pipelined.layer_1_compressor42_0.B , \multiplier_16x16bit_pipelined.layer_1_full_adder_1.B , \multiplier_16x16bit_pipelined.layer_1_full_adder_0.B , \multiplier_16x16bit_pipelined.layer_0_w3[1] , \multiplier_16x16bit_pipelined.layer_0_w2[1] } = fangyuan76;
  wire [15:0] fangyuan77;
  assign fangyuan77 = { \multiplier_16x16bit_pipelined.partial_product_gen_1.zmd [14:0], \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_1.negation };

  assign fangyuan76 = \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_1.double ? fangyuan77 : \multiplier_16x16bit_pipelined.partial_product_gen_1.zmd ;
  assign \multiplier_16x16bit_pipelined.layer_1_compressor42_13.A = ~ \multiplier_16x16bit_pipelined.partial_product_gen_2.zmd [15];
  assign \multiplier_16x16bit_pipelined.partial_product_gen_2.nmd = \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_2.negation ? _0517_ : \multiplier_16x16bit_pipelined.md ;
  assign \multiplier_16x16bit_pipelined.partial_product_gen_2.zmd = \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_2.zero ? 16'b0000000000000000 : \multiplier_16x16bit_pipelined.partial_product_gen_2.nmd ;
  wire [15:0] fangyuan78;
  assign { \multiplier_16x16bit_pipelined.layer_1_compressor42_12.A , \multiplier_16x16bit_pipelined.layer_1_compressor42_11.B , \multiplier_16x16bit_pipelined.layer_1_compressor42_10.B , \multiplier_16x16bit_pipelined.layer_1_compressor42_9.C , \multiplier_16x16bit_pipelined.layer_1_compressor42_8.C , \multiplier_16x16bit_pipelined.layer_1_compressor42_7.C , \multiplier_16x16bit_pipelined.layer_1_compressor42_6.C , \multiplier_16x16bit_pipelined.layer_1_compressor42_5.C , \multiplier_16x16bit_pipelined.layer_1_compressor42_4.C , \multiplier_16x16bit_pipelined.layer_1_compressor42_3.C , \multiplier_16x16bit_pipelined.layer_1_compressor42_2.C , \multiplier_16x16bit_pipelined.layer_1_compressor42_1.C , \multiplier_16x16bit_pipelined.layer_1_full_adder_2.cin , \multiplier_16x16bit_pipelined.layer_1_compressor42_0.C , \multiplier_16x16bit_pipelined.layer_1_full_adder_1.cin , \multiplier_16x16bit_pipelined.layer_1_full_adder_0.cin } = fangyuan78;
  wire [15:0] fangyuan79;
  assign fangyuan79 = { \multiplier_16x16bit_pipelined.partial_product_gen_2.zmd [14:0], \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_2.negation };

  assign fangyuan78 = \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_2.double ? fangyuan79 : \multiplier_16x16bit_pipelined.partial_product_gen_2.zmd ;
  assign \multiplier_16x16bit_pipelined.layer_1_compressor42_15.A = ~ \multiplier_16x16bit_pipelined.partial_product_gen_3.zmd [15];
  assign \multiplier_16x16bit_pipelined.partial_product_gen_3.nmd = \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_3.negation ? _0517_ : \multiplier_16x16bit_pipelined.md ;
  assign \multiplier_16x16bit_pipelined.partial_product_gen_3.zmd = \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_3.zero ? 16'b0000000000000000 : \multiplier_16x16bit_pipelined.partial_product_gen_3.nmd ;
  wire [15:0] fangyuan80;
  assign { \multiplier_16x16bit_pipelined.layer_1_compressor42_14.A , \multiplier_16x16bit_pipelined.layer_1_compressor42_13.B , \multiplier_16x16bit_pipelined.layer_1_compressor42_12.B , \multiplier_16x16bit_pipelined.layer_1_compressor42_11.C , \multiplier_16x16bit_pipelined.layer_1_compressor42_10.C , \multiplier_16x16bit_pipelined.layer_1_compressor42_9.D , \multiplier_16x16bit_pipelined.layer_1_compressor42_8.D , \multiplier_16x16bit_pipelined.layer_1_compressor42_7.D , \multiplier_16x16bit_pipelined.layer_1_compressor42_6.D , \multiplier_16x16bit_pipelined.layer_1_compressor42_5.D , \multiplier_16x16bit_pipelined.layer_1_compressor42_4.D , \multiplier_16x16bit_pipelined.layer_1_compressor42_3.D , \multiplier_16x16bit_pipelined.layer_1_compressor42_2.D , \multiplier_16x16bit_pipelined.layer_1_compressor42_1.D , \multiplier_16x16bit_pipelined.layer_0_w7[3] , \multiplier_16x16bit_pipelined.layer_1_compressor42_0.D } = fangyuan80;
  wire [15:0] fangyuan81;
  assign fangyuan81 = { \multiplier_16x16bit_pipelined.partial_product_gen_3.zmd [14:0], \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_3.negation };

  assign fangyuan80 = \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_3.double ? fangyuan81 : \multiplier_16x16bit_pipelined.partial_product_gen_3.zmd ;
  assign \multiplier_16x16bit_pipelined.layer_1_full_adder_8.A = ~ \multiplier_16x16bit_pipelined.partial_product_gen_4.zmd [15];
  assign \multiplier_16x16bit_pipelined.partial_product_gen_4.nmd = \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_4.negation ? _0517_ : \multiplier_16x16bit_pipelined.md ;
  assign \multiplier_16x16bit_pipelined.partial_product_gen_4.zmd = \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_4.zero ? 16'b0000000000000000 : \multiplier_16x16bit_pipelined.partial_product_gen_4.nmd ;
  wire [15:0] fangyuan82;
  assign { \multiplier_16x16bit_pipelined.layer_1_compressor42_16.A , \multiplier_16x16bit_pipelined.layer_1_compressor42_15.B , \multiplier_16x16bit_pipelined.layer_1_compressor42_14.B , \multiplier_16x16bit_pipelined.layer_1_compressor42_13.C , \multiplier_16x16bit_pipelined.layer_1_compressor42_12.C , \multiplier_16x16bit_pipelined.layer_1_compressor42_11.D , \multiplier_16x16bit_pipelined.layer_1_compressor42_10.D , \multiplier_16x16bit_pipelined.layer_1_compressor42_9.cin , \multiplier_16x16bit_pipelined.layer_1_compressor42_8.cin , \multiplier_16x16bit_pipelined.layer_1_compressor42_7.cin , \multiplier_16x16bit_pipelined.layer_1_compressor42_6.cin , \multiplier_16x16bit_pipelined.layer_1_compressor42_5.cin , \multiplier_16x16bit_pipelined.layer_1_compressor42_4.cin , \multiplier_16x16bit_pipelined.layer_1_compressor42_3.cin , \multiplier_16x16bit_pipelined.layer_1_compressor42_2.cin , \multiplier_16x16bit_pipelined.layer_1_compressor42_1.cin } = fangyuan82;
  wire [15:0] fangyuan83;
  assign fangyuan83 = { \multiplier_16x16bit_pipelined.partial_product_gen_4.zmd [14:0], \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_4.negation };

  assign fangyuan82 = \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_4.double ? fangyuan83 : \multiplier_16x16bit_pipelined.partial_product_gen_4.zmd ;
  assign \multiplier_16x16bit_pipelined.layer_1_full_adder_10.A = ~ \multiplier_16x16bit_pipelined.partial_product_gen_5.zmd [15];
  assign \multiplier_16x16bit_pipelined.partial_product_gen_5.nmd = \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_5.negation ? _0517_ : \multiplier_16x16bit_pipelined.md ;
  assign \multiplier_16x16bit_pipelined.partial_product_gen_5.zmd = \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_5.zero ? 16'b0000000000000000 : \multiplier_16x16bit_pipelined.partial_product_gen_5.nmd ;
  wire [15:0] fangyuan84;
  assign { \multiplier_16x16bit_pipelined.layer_1_full_adder_9.A , \multiplier_16x16bit_pipelined.layer_1_full_adder_8.B , \multiplier_16x16bit_pipelined.layer_1_compressor42_16.B , \multiplier_16x16bit_pipelined.layer_1_compressor42_15.C , \multiplier_16x16bit_pipelined.layer_1_compressor42_14.C , \multiplier_16x16bit_pipelined.layer_1_compressor42_13.D , \multiplier_16x16bit_pipelined.layer_1_compressor42_12.D , \multiplier_16x16bit_pipelined.layer_1_compressor42_11.cin , \multiplier_16x16bit_pipelined.layer_1_compressor42_10.cin , \multiplier_16x16bit_pipelined.layer_1_full_adder_6.A , \multiplier_16x16bit_pipelined.layer_1_full_adder_5.A , \multiplier_16x16bit_pipelined.layer_1_full_adder_4.A , \multiplier_16x16bit_pipelined.layer_2_compressor42_1.cin , \multiplier_16x16bit_pipelined.layer_1_full_adder_3.A , \multiplier_16x16bit_pipelined.layer_0_w11[5] , \multiplier_16x16bit_pipelined.layer_2_compressor42_0.D } = fangyuan84;
  wire [15:0] fangyuan85;
  assign fangyuan85 = { \multiplier_16x16bit_pipelined.partial_product_gen_5.zmd [14:0], \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_5.negation };

  assign fangyuan84 = \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_5.double ? fangyuan85 : \multiplier_16x16bit_pipelined.partial_product_gen_5.zmd ;
  assign \multiplier_16x16bit_pipelined.layer_2_full_adder_11.B = ~ \multiplier_16x16bit_pipelined.partial_product_gen_6.zmd [15];
  assign \multiplier_16x16bit_pipelined.partial_product_gen_6.nmd = \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_6.negation ? _0517_ : \multiplier_16x16bit_pipelined.md ;
  assign \multiplier_16x16bit_pipelined.partial_product_gen_6.zmd = \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_6.zero ? 16'b0000000000000000 : \multiplier_16x16bit_pipelined.partial_product_gen_6.nmd ;
  wire [15:0] fangyuan86;
  assign { \multiplier_16x16bit_pipelined.layer_1_full_adder_11.A , \multiplier_16x16bit_pipelined.layer_1_full_adder_10.B , \multiplier_16x16bit_pipelined.layer_1_full_adder_9.B , \multiplier_16x16bit_pipelined.layer_1_full_adder_8.cin , \multiplier_16x16bit_pipelined.layer_1_compressor42_16.C , \multiplier_16x16bit_pipelined.layer_1_compressor42_15.D , \multiplier_16x16bit_pipelined.layer_1_compressor42_14.D , \multiplier_16x16bit_pipelined.layer_1_compressor42_13.cin , \multiplier_16x16bit_pipelined.layer_1_compressor42_12.cin , \multiplier_16x16bit_pipelined.layer_2_compressor42_6.cin , \multiplier_16x16bit_pipelined.layer_1_full_adder_7.A , \multiplier_16x16bit_pipelined.layer_1_full_adder_6.B , \multiplier_16x16bit_pipelined.layer_1_full_adder_5.B , \multiplier_16x16bit_pipelined.layer_1_full_adder_4.B , \multiplier_16x16bit_pipelined.layer_0_w13[6] , \multiplier_16x16bit_pipelined.layer_1_full_adder_3.B } = fangyuan86;
  wire [15:0] fangyuan87;
  assign fangyuan87 = { \multiplier_16x16bit_pipelined.partial_product_gen_6.zmd [14:0], \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_6.negation };

  assign fangyuan86 = \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_6.double ? fangyuan87 : \multiplier_16x16bit_pipelined.partial_product_gen_6.zmd ;
  assign \multiplier_16x16bit_pipelined.layer_0_w30 = ~ \multiplier_16x16bit_pipelined.partial_product_gen_7.zmd [15];
  assign \multiplier_16x16bit_pipelined.partial_product_gen_7.nmd = \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_7.negation ? _0517_ : \multiplier_16x16bit_pipelined.md ;
  assign \multiplier_16x16bit_pipelined.partial_product_gen_7.zmd = \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_7.zero ? 16'b0000000000000000 : \multiplier_16x16bit_pipelined.partial_product_gen_7.nmd ;
  wire [15:0] fangyuan88;
  assign { \multiplier_16x16bit_pipelined.layer_0_w29[0] , \multiplier_16x16bit_pipelined.layer_2_full_adder_11.cin , \multiplier_16x16bit_pipelined.layer_1_full_adder_11.B , \multiplier_16x16bit_pipelined.layer_1_full_adder_10.cin , \multiplier_16x16bit_pipelined.layer_1_full_adder_9.cin , \multiplier_16x16bit_pipelined.layer_0_w24[3] , \multiplier_16x16bit_pipelined.layer_1_compressor42_16.D , \multiplier_16x16bit_pipelined.layer_1_compressor42_15.cin , \multiplier_16x16bit_pipelined.layer_1_compressor42_14.cin , \multiplier_16x16bit_pipelined.layer_0_w20[5] , \multiplier_16x16bit_pipelined.layer_2_compressor42_7.D , \multiplier_16x16bit_pipelined.layer_0_w18[6] , \multiplier_16x16bit_pipelined.layer_1_full_adder_7.B , \multiplier_16x16bit_pipelined.layer_1_full_adder_6.cin , \multiplier_16x16bit_pipelined.layer_1_full_adder_5.cin , \multiplier_16x16bit_pipelined.layer_1_full_adder_4.cin } = fangyuan88;
  wire [15:0] fangyuan89;
  assign fangyuan89 = { \multiplier_16x16bit_pipelined.partial_product_gen_7.zmd [14:0], \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_7.negation };

  assign fangyuan88 = \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_7.double ? fangyuan89 : \multiplier_16x16bit_pipelined.partial_product_gen_7.zmd ;
  assign _0518_ = _0043_ ? kd : ki;
  assign mr = _0042_ ? kpd : _0518_;
  assign _0519_ = _0045_ ? \err[0] : \adder_32bit_0.o_s [15:0];
  assign md = _0044_ ? \err[1] : _0519_;
  assign o_wb_data = adr_check_1 ? _0000_ : 32'd0;
  assign \adder_32bit_0.G0 [30:0] = { \adder_32bit_0.operator_A_30.G , \adder_32bit_0.operator_A_29.G , \adder_32bit_0.operator_A_28.G , \adder_32bit_0.operator_A_27.G , \adder_32bit_0.operator_A_26.G , \adder_32bit_0.operator_A_25.G , \adder_32bit_0.operator_A_24.G , \adder_32bit_0.operator_A_23.G , \adder_32bit_0.operator_A_22.G , \adder_32bit_0.operator_A_21.G , \adder_32bit_0.operator_A_20.G , \adder_32bit_0.operator_A_19.G , \adder_32bit_0.operator_A_18.G , \adder_32bit_0.operator_A_17.G , \adder_32bit_0.operator_A_16.G , \adder_32bit_0.operator_A_15.G , \adder_32bit_0.operator_A_14.G , \adder_32bit_0.operator_A_13.G , \adder_32bit_0.operator_A_12.G , \adder_32bit_0.operator_A_11.G , \adder_32bit_0.operator_A_10.G , \adder_32bit_0.operator_A_9.G , \adder_32bit_0.operator_A_8.G , \adder_32bit_0.operator_A_7.G , \adder_32bit_0.operator_A_6.G , \adder_32bit_0.operator_A_5.G , \adder_32bit_0.operator_A_4.G , \adder_32bit_0.operator_A_3.G , \adder_32bit_0.operator_A_2.G , \adder_32bit_0.operator_A_1.G , \adder_32bit_0.operator_A_0.G };
  assign \adder_32bit_0.G1 = { \adder_32bit_0.operator_B_stage_1_15.Go , \adder_32bit_0.operator_B_stage_1_14.Go , \adder_32bit_0.operator_B_stage_1_13.Go , \adder_32bit_0.operator_B_stage_1_12.Go , \adder_32bit_0.operator_B_stage_1_11.Go , \adder_32bit_0.operator_B_stage_1_10.Go , \adder_32bit_0.operator_B_stage_1_9.Go , \adder_32bit_0.operator_B_stage_1_8.Go , \adder_32bit_0.operator_B_stage_1_7.Go , \adder_32bit_0.operator_B_stage_1_6.Go , \adder_32bit_0.operator_B_stage_1_5.Go , \adder_32bit_0.operator_B_stage_1_4.Go , \adder_32bit_0.operator_B_stage_1_3.Go , \adder_32bit_0.operator_B_stage_1_2.Go , \adder_32bit_0.operator_B_stage_1_1.Go , \adder_32bit_0.operator_C_stage_1_0.Go };
  assign \adder_32bit_0.G2 = { \adder_32bit_0.operator_B_stage_2_15.Go , \adder_32bit_0.operator_B_stage_2_14.Go , \adder_32bit_0.operator_B_stage_2_13.Go , \adder_32bit_0.operator_B_stage_2_12.Go , \adder_32bit_0.operator_B_stage_2_11.Go , \adder_32bit_0.operator_B_stage_2_10.Go , \adder_32bit_0.operator_B_stage_2_9.Go , \adder_32bit_0.operator_B_stage_2_8.Go , \adder_32bit_0.operator_B_stage_2_7.Go , \adder_32bit_0.operator_B_stage_2_6.Go , \adder_32bit_0.operator_B_stage_2_5.Go , \adder_32bit_0.operator_B_stage_2_4.Go , \adder_32bit_0.operator_B_stage_2_3.Go , \adder_32bit_0.operator_B_stage_2_2.Go , \adder_32bit_0.operator_C_stage_2_1.Go , \adder_32bit_0.operator_C_stage_1_0.Go };
  assign \adder_32bit_0.G3 = { \adder_32bit_0.operator_B_stage_3_15.Go , \adder_32bit_0.operator_B_stage_3_14.Go , \adder_32bit_0.operator_B_stage_3_13.Go , \adder_32bit_0.operator_B_stage_3_12.Go , \adder_32bit_0.operator_B_stage_3_11.Go , \adder_32bit_0.operator_B_stage_3_10.Go , \adder_32bit_0.operator_B_stage_3_9.Go , \adder_32bit_0.operator_B_stage_3_8.Go , \adder_32bit_0.operator_B_stage_3_7.Go , \adder_32bit_0.operator_B_stage_3_6.Go , \adder_32bit_0.operator_B_stage_3_5.Go , \adder_32bit_0.operator_B_stage_3_4.Go , \adder_32bit_0.operator_C_stage_3_3.Go , \adder_32bit_0.operator_C_stage_3_2.Go , \adder_32bit_0.operator_C_stage_2_1.Go , \adder_32bit_0.operator_C_stage_1_0.Go };
  assign \adder_32bit_0.G4 = { \adder_32bit_0.operator_B_stage_4_15.Go , \adder_32bit_0.operator_B_stage_4_14.Go , \adder_32bit_0.operator_B_stage_4_13.Go , \adder_32bit_0.operator_B_stage_4_12.Go , \adder_32bit_0.operator_B_stage_4_11.Go , \adder_32bit_0.operator_B_stage_4_10.Go , \adder_32bit_0.operator_B_stage_4_9.Go , \adder_32bit_0.operator_B_stage_4_8.Go , \adder_32bit_0.operator_C_stage_4_7.Go , \adder_32bit_0.operator_C_stage_4_6.Go , \adder_32bit_0.operator_C_stage_4_5.Go , \adder_32bit_0.operator_C_stage_4_4.Go , \adder_32bit_0.operator_C_stage_3_3.Go , \adder_32bit_0.operator_C_stage_3_2.Go , \adder_32bit_0.operator_C_stage_2_1.Go , \adder_32bit_0.operator_C_stage_1_0.Go };
  assign \adder_32bit_0.G5 = { \adder_32bit_0.operator_C_stage_5_15.Go , \adder_32bit_0.operator_C_stage_5_14.Go , \adder_32bit_0.operator_C_stage_5_13.Go , \adder_32bit_0.operator_C_stage_5_12.Go , \adder_32bit_0.operator_C_stage_5_11.Go , \adder_32bit_0.operator_C_stage_5_10.Go , \adder_32bit_0.operator_C_stage_5_9.Go , \adder_32bit_0.operator_C_stage_5_8.Go , \adder_32bit_0.operator_C_stage_4_7.Go , \adder_32bit_0.operator_C_stage_4_6.Go , \adder_32bit_0.operator_C_stage_4_5.Go , \adder_32bit_0.operator_C_stage_4_4.Go , \adder_32bit_0.operator_C_stage_3_3.Go , \adder_32bit_0.operator_C_stage_3_2.Go , \adder_32bit_0.operator_C_stage_2_1.Go , \adder_32bit_0.operator_C_stage_1_0.Go };
  assign \adder_32bit_0.G6 [30:0] = { \adder_32bit_0.operator_C_stage_5_15.Go , \adder_32bit_0.operator_C_stage_6_14.Go , \adder_32bit_0.operator_C_stage_5_14.Go , \adder_32bit_0.operator_C_stage_6_13.Go , \adder_32bit_0.operator_C_stage_5_13.Go , \adder_32bit_0.operator_C_stage_6_12.Go , \adder_32bit_0.operator_C_stage_5_12.Go , \adder_32bit_0.operator_C_stage_6_11.Go , \adder_32bit_0.operator_C_stage_5_11.Go , \adder_32bit_0.operator_C_stage_6_10.Go , \adder_32bit_0.operator_C_stage_5_10.Go , \adder_32bit_0.operator_C_stage_6_9.Go , \adder_32bit_0.operator_C_stage_5_9.Go , \adder_32bit_0.operator_C_stage_6_8.Go , \adder_32bit_0.operator_C_stage_5_8.Go , \adder_32bit_0.operator_C_stage_6_7.Go , \adder_32bit_0.operator_C_stage_4_7.Go , \adder_32bit_0.operator_C_stage_6_6.Go , \adder_32bit_0.operator_C_stage_4_6.Go , \adder_32bit_0.operator_C_stage_6_5.Go , \adder_32bit_0.operator_C_stage_4_5.Go , \adder_32bit_0.operator_C_stage_6_4.Go , \adder_32bit_0.operator_C_stage_4_4.Go , \adder_32bit_0.operator_C_stage_6_3.Go , \adder_32bit_0.operator_C_stage_3_3.Go , \adder_32bit_0.operator_C_stage_6_2.Go , \adder_32bit_0.operator_C_stage_3_2.Go , \adder_32bit_0.operator_C_stage_6_1.Go , \adder_32bit_0.operator_C_stage_2_1.Go , \adder_32bit_0.operator_C_stage_6_0.Go , \adder_32bit_0.operator_C_stage_1_0.Go };
  assign \adder_32bit_0.P0 = { \adder_32bit_0.operator_A_31.P , \adder_32bit_0.operator_A_30.P , \adder_32bit_0.operator_A_29.P , \adder_32bit_0.operator_A_28.P , \adder_32bit_0.operator_A_27.P , \adder_32bit_0.operator_A_26.P , \adder_32bit_0.operator_A_25.P , \adder_32bit_0.operator_A_24.P , \adder_32bit_0.operator_A_23.P , \adder_32bit_0.operator_A_22.P , \adder_32bit_0.operator_A_21.P , \adder_32bit_0.operator_A_20.P , \adder_32bit_0.operator_A_19.P , \adder_32bit_0.operator_A_18.P , \adder_32bit_0.operator_A_17.P , \adder_32bit_0.operator_A_16.P , \adder_32bit_0.operator_A_15.P , \adder_32bit_0.operator_A_14.P , \adder_32bit_0.operator_A_13.P , \adder_32bit_0.operator_A_12.P , \adder_32bit_0.operator_A_11.P , \adder_32bit_0.operator_A_10.P , \adder_32bit_0.operator_A_9.P , \adder_32bit_0.operator_A_8.P , \adder_32bit_0.operator_A_7.P , \adder_32bit_0.operator_A_6.P , \adder_32bit_0.operator_A_5.P , \adder_32bit_0.operator_A_4.P , \adder_32bit_0.operator_A_3.P , \adder_32bit_0.operator_A_2.P , \adder_32bit_0.operator_A_1.P , \adder_32bit_0.operator_A_0.P };
  assign \adder_32bit_0.P1 = { \adder_32bit_0.operator_B_stage_1_15.Po , \adder_32bit_0.operator_B_stage_1_14.Po , \adder_32bit_0.operator_B_stage_1_13.Po , \adder_32bit_0.operator_B_stage_1_12.Po , \adder_32bit_0.operator_B_stage_1_11.Po , \adder_32bit_0.operator_B_stage_1_10.Po , \adder_32bit_0.operator_B_stage_1_9.Po , \adder_32bit_0.operator_B_stage_1_8.Po , \adder_32bit_0.operator_B_stage_1_7.Po , \adder_32bit_0.operator_B_stage_1_6.Po , \adder_32bit_0.operator_B_stage_1_5.Po , \adder_32bit_0.operator_B_stage_1_4.Po , \adder_32bit_0.operator_B_stage_1_3.Po , \adder_32bit_0.operator_B_stage_1_2.Po , \adder_32bit_0.operator_B_stage_1_1.Po };
  assign \adder_32bit_0.P2 = { \adder_32bit_0.operator_B_stage_2_15.Po , \adder_32bit_0.operator_B_stage_2_14.Po , \adder_32bit_0.operator_B_stage_2_13.Po , \adder_32bit_0.operator_B_stage_2_12.Po , \adder_32bit_0.operator_B_stage_2_11.Po , \adder_32bit_0.operator_B_stage_2_10.Po , \adder_32bit_0.operator_B_stage_2_9.Po , \adder_32bit_0.operator_B_stage_2_8.Po , \adder_32bit_0.operator_B_stage_2_7.Po , \adder_32bit_0.operator_B_stage_2_6.Po , \adder_32bit_0.operator_B_stage_2_5.Po , \adder_32bit_0.operator_B_stage_2_4.Po , \adder_32bit_0.operator_B_stage_2_3.Po , \adder_32bit_0.operator_B_stage_2_2.Po };
  assign \adder_32bit_0.P3 = { \adder_32bit_0.operator_B_stage_3_15.Po , \adder_32bit_0.operator_B_stage_3_14.Po , \adder_32bit_0.operator_B_stage_3_13.Po , \adder_32bit_0.operator_B_stage_3_12.Po , \adder_32bit_0.operator_B_stage_3_11.Po , \adder_32bit_0.operator_B_stage_3_10.Po , \adder_32bit_0.operator_B_stage_3_9.Po , \adder_32bit_0.operator_B_stage_3_8.Po , \adder_32bit_0.operator_B_stage_3_7.Po , \adder_32bit_0.operator_B_stage_3_6.Po , \adder_32bit_0.operator_B_stage_3_5.Po , \adder_32bit_0.operator_B_stage_3_4.Po };
  assign \adder_32bit_0.P4 = { \adder_32bit_0.operator_B_stage_4_15.Po , \adder_32bit_0.operator_B_stage_4_14.Po , \adder_32bit_0.operator_B_stage_4_13.Po , \adder_32bit_0.operator_B_stage_4_12.Po , \adder_32bit_0.operator_B_stage_4_11.Po , \adder_32bit_0.operator_B_stage_4_10.Po , \adder_32bit_0.operator_B_stage_4_9.Po , \adder_32bit_0.operator_B_stage_4_8.Po };
  assign \adder_32bit_0.i_a = a;
  assign \adder_32bit_0.i_b = p;
  assign \adder_32bit_0.i_c = cout;
  assign \adder_32bit_0.operator_A_0.A = a[0];
  assign \adder_32bit_0.operator_A_0.B = p[0];
  assign \adder_32bit_0.operator_A_1.A = a[1];
  assign \adder_32bit_0.operator_A_1.B = p[1];
  assign \adder_32bit_0.operator_A_10.A = a[10];
  assign \adder_32bit_0.operator_A_10.B = p[10];
  assign \adder_32bit_0.operator_A_11.A = a[11];
  assign \adder_32bit_0.operator_A_11.B = p[11];
  assign \adder_32bit_0.operator_A_12.A = a[12];
  assign \adder_32bit_0.operator_A_12.B = p[12];
  assign \adder_32bit_0.operator_A_13.A = a[13];
  assign \adder_32bit_0.operator_A_13.B = p[13];
  assign \adder_32bit_0.operator_A_14.A = a[14];
  assign \adder_32bit_0.operator_A_14.B = p[14];
  assign \adder_32bit_0.operator_A_15.A = a[15];
  assign \adder_32bit_0.operator_A_15.B = p[15];
  assign \adder_32bit_0.operator_A_16.A = a[16];
  assign \adder_32bit_0.operator_A_16.B = p[16];
  assign \adder_32bit_0.operator_A_17.A = a[17];
  assign \adder_32bit_0.operator_A_17.B = p[17];
  assign \adder_32bit_0.operator_A_18.A = a[18];
  assign \adder_32bit_0.operator_A_18.B = p[18];
  assign \adder_32bit_0.operator_A_19.A = a[19];
  assign \adder_32bit_0.operator_A_19.B = p[19];
  assign \adder_32bit_0.operator_A_2.A = a[2];
  assign \adder_32bit_0.operator_A_2.B = p[2];
  assign \adder_32bit_0.operator_A_20.A = a[20];
  assign \adder_32bit_0.operator_A_20.B = p[20];
  assign \adder_32bit_0.operator_A_21.A = a[21];
  assign \adder_32bit_0.operator_A_21.B = p[21];
  assign \adder_32bit_0.operator_A_22.A = a[22];
  assign \adder_32bit_0.operator_A_22.B = p[22];
  assign \adder_32bit_0.operator_A_23.A = a[23];
  assign \adder_32bit_0.operator_A_23.B = p[23];
  assign \adder_32bit_0.operator_A_24.A = a[24];
  assign \adder_32bit_0.operator_A_24.B = p[24];
  assign \adder_32bit_0.operator_A_25.A = a[25];
  assign \adder_32bit_0.operator_A_25.B = p[25];
  assign \adder_32bit_0.operator_A_26.A = a[26];
  assign \adder_32bit_0.operator_A_26.B = p[26];
  assign \adder_32bit_0.operator_A_27.A = a[27];
  assign \adder_32bit_0.operator_A_27.B = p[27];
  assign \adder_32bit_0.operator_A_28.A = a[28];
  assign \adder_32bit_0.operator_A_28.B = p[28];
  assign \adder_32bit_0.operator_A_29.A = a[29];
  assign \adder_32bit_0.operator_A_29.B = p[29];
  assign \adder_32bit_0.operator_A_3.A = a[3];
  assign \adder_32bit_0.operator_A_3.B = p[3];
  assign \adder_32bit_0.operator_A_30.A = a[30];
  assign \adder_32bit_0.operator_A_30.B = p[30];
  assign \adder_32bit_0.operator_A_31.A = a[31];
  assign \adder_32bit_0.operator_A_31.B = p[31];
  assign \adder_32bit_0.operator_A_4.A = a[4];
  assign \adder_32bit_0.operator_A_4.B = p[4];
  assign \adder_32bit_0.operator_A_5.A = a[5];
  assign \adder_32bit_0.operator_A_5.B = p[5];
  assign \adder_32bit_0.operator_A_6.A = a[6];
  assign \adder_32bit_0.operator_A_6.B = p[6];
  assign \adder_32bit_0.operator_A_7.A = a[7];
  assign \adder_32bit_0.operator_A_7.B = p[7];
  assign \adder_32bit_0.operator_A_8.A = a[8];
  assign \adder_32bit_0.operator_A_8.B = p[8];
  assign \adder_32bit_0.operator_A_9.A = a[9];
  assign \adder_32bit_0.operator_A_9.B = p[9];
  assign \adder_32bit_0.operator_B_stage_1_1.G = \adder_32bit_0.operator_A_2.G ;
  assign \adder_32bit_0.operator_B_stage_1_1.G1 = \adder_32bit_0.operator_A_1.G ;
  assign \adder_32bit_0.operator_B_stage_1_1.P = \adder_32bit_0.operator_A_2.P ;
  assign \adder_32bit_0.operator_B_stage_1_1.P1 = \adder_32bit_0.operator_A_1.P ;
  assign \adder_32bit_0.operator_B_stage_1_10.G = \adder_32bit_0.operator_A_20.G ;
  assign \adder_32bit_0.operator_B_stage_1_10.G1 = \adder_32bit_0.operator_A_19.G ;
  assign \adder_32bit_0.operator_B_stage_1_10.P = \adder_32bit_0.operator_A_20.P ;
  assign \adder_32bit_0.operator_B_stage_1_10.P1 = \adder_32bit_0.operator_A_19.P ;
  assign \adder_32bit_0.operator_B_stage_1_11.G = \adder_32bit_0.operator_A_22.G ;
  assign \adder_32bit_0.operator_B_stage_1_11.G1 = \adder_32bit_0.operator_A_21.G ;
  assign \adder_32bit_0.operator_B_stage_1_11.P = \adder_32bit_0.operator_A_22.P ;
  assign \adder_32bit_0.operator_B_stage_1_11.P1 = \adder_32bit_0.operator_A_21.P ;
  assign \adder_32bit_0.operator_B_stage_1_12.G = \adder_32bit_0.operator_A_24.G ;
  assign \adder_32bit_0.operator_B_stage_1_12.G1 = \adder_32bit_0.operator_A_23.G ;
  assign \adder_32bit_0.operator_B_stage_1_12.P = \adder_32bit_0.operator_A_24.P ;
  assign \adder_32bit_0.operator_B_stage_1_12.P1 = \adder_32bit_0.operator_A_23.P ;
  assign \adder_32bit_0.operator_B_stage_1_13.G = \adder_32bit_0.operator_A_26.G ;
  assign \adder_32bit_0.operator_B_stage_1_13.G1 = \adder_32bit_0.operator_A_25.G ;
  assign \adder_32bit_0.operator_B_stage_1_13.P = \adder_32bit_0.operator_A_26.P ;
  assign \adder_32bit_0.operator_B_stage_1_13.P1 = \adder_32bit_0.operator_A_25.P ;
  assign \adder_32bit_0.operator_B_stage_1_14.G = \adder_32bit_0.operator_A_28.G ;
  assign \adder_32bit_0.operator_B_stage_1_14.G1 = \adder_32bit_0.operator_A_27.G ;
  assign \adder_32bit_0.operator_B_stage_1_14.P = \adder_32bit_0.operator_A_28.P ;
  assign \adder_32bit_0.operator_B_stage_1_14.P1 = \adder_32bit_0.operator_A_27.P ;
  assign \adder_32bit_0.operator_B_stage_1_15.G = \adder_32bit_0.operator_A_30.G ;
  assign \adder_32bit_0.operator_B_stage_1_15.G1 = \adder_32bit_0.operator_A_29.G ;
  assign \adder_32bit_0.operator_B_stage_1_15.P = \adder_32bit_0.operator_A_30.P ;
  assign \adder_32bit_0.operator_B_stage_1_15.P1 = \adder_32bit_0.operator_A_29.P ;
  assign \adder_32bit_0.operator_B_stage_1_2.G = \adder_32bit_0.operator_A_4.G ;
  assign \adder_32bit_0.operator_B_stage_1_2.G1 = \adder_32bit_0.operator_A_3.G ;
  assign \adder_32bit_0.operator_B_stage_1_2.P = \adder_32bit_0.operator_A_4.P ;
  assign \adder_32bit_0.operator_B_stage_1_2.P1 = \adder_32bit_0.operator_A_3.P ;
  assign \adder_32bit_0.operator_B_stage_1_3.G = \adder_32bit_0.operator_A_6.G ;
  assign \adder_32bit_0.operator_B_stage_1_3.G1 = \adder_32bit_0.operator_A_5.G ;
  assign \adder_32bit_0.operator_B_stage_1_3.P = \adder_32bit_0.operator_A_6.P ;
  assign \adder_32bit_0.operator_B_stage_1_3.P1 = \adder_32bit_0.operator_A_5.P ;
  assign \adder_32bit_0.operator_B_stage_1_4.G = \adder_32bit_0.operator_A_8.G ;
  assign \adder_32bit_0.operator_B_stage_1_4.G1 = \adder_32bit_0.operator_A_7.G ;
  assign \adder_32bit_0.operator_B_stage_1_4.P = \adder_32bit_0.operator_A_8.P ;
  assign \adder_32bit_0.operator_B_stage_1_4.P1 = \adder_32bit_0.operator_A_7.P ;
  assign \adder_32bit_0.operator_B_stage_1_5.G = \adder_32bit_0.operator_A_10.G ;
  assign \adder_32bit_0.operator_B_stage_1_5.G1 = \adder_32bit_0.operator_A_9.G ;
  assign \adder_32bit_0.operator_B_stage_1_5.P = \adder_32bit_0.operator_A_10.P ;
  assign \adder_32bit_0.operator_B_stage_1_5.P1 = \adder_32bit_0.operator_A_9.P ;
  assign \adder_32bit_0.operator_B_stage_1_6.G = \adder_32bit_0.operator_A_12.G ;
  assign \adder_32bit_0.operator_B_stage_1_6.G1 = \adder_32bit_0.operator_A_11.G ;
  assign \adder_32bit_0.operator_B_stage_1_6.P = \adder_32bit_0.operator_A_12.P ;
  assign \adder_32bit_0.operator_B_stage_1_6.P1 = \adder_32bit_0.operator_A_11.P ;
  assign \adder_32bit_0.operator_B_stage_1_7.G = \adder_32bit_0.operator_A_14.G ;
  assign \adder_32bit_0.operator_B_stage_1_7.G1 = \adder_32bit_0.operator_A_13.G ;
  assign \adder_32bit_0.operator_B_stage_1_7.P = \adder_32bit_0.operator_A_14.P ;
  assign \adder_32bit_0.operator_B_stage_1_7.P1 = \adder_32bit_0.operator_A_13.P ;
  assign \adder_32bit_0.operator_B_stage_1_8.G = \adder_32bit_0.operator_A_16.G ;
  assign \adder_32bit_0.operator_B_stage_1_8.G1 = \adder_32bit_0.operator_A_15.G ;
  assign \adder_32bit_0.operator_B_stage_1_8.P = \adder_32bit_0.operator_A_16.P ;
  assign \adder_32bit_0.operator_B_stage_1_8.P1 = \adder_32bit_0.operator_A_15.P ;
  assign \adder_32bit_0.operator_B_stage_1_9.G = \adder_32bit_0.operator_A_18.G ;
  assign \adder_32bit_0.operator_B_stage_1_9.G1 = \adder_32bit_0.operator_A_17.G ;
  assign \adder_32bit_0.operator_B_stage_1_9.P = \adder_32bit_0.operator_A_18.P ;
  assign \adder_32bit_0.operator_B_stage_1_9.P1 = \adder_32bit_0.operator_A_17.P ;
  assign \adder_32bit_0.operator_B_stage_2_10.G = \adder_32bit_0.operator_B_stage_1_10.Go ;
  assign \adder_32bit_0.operator_B_stage_2_10.G1 = \adder_32bit_0.operator_B_stage_1_9.Go ;
  assign \adder_32bit_0.operator_B_stage_2_10.P = \adder_32bit_0.operator_B_stage_1_10.Po ;
  assign \adder_32bit_0.operator_B_stage_2_10.P1 = \adder_32bit_0.operator_B_stage_1_9.Po ;
  assign \adder_32bit_0.operator_B_stage_2_11.G = \adder_32bit_0.operator_B_stage_1_11.Go ;
  assign \adder_32bit_0.operator_B_stage_2_11.G1 = \adder_32bit_0.operator_B_stage_1_10.Go ;
  assign \adder_32bit_0.operator_B_stage_2_11.P = \adder_32bit_0.operator_B_stage_1_11.Po ;
  assign \adder_32bit_0.operator_B_stage_2_11.P1 = \adder_32bit_0.operator_B_stage_1_10.Po ;
  assign \adder_32bit_0.operator_B_stage_2_12.G = \adder_32bit_0.operator_B_stage_1_12.Go ;
  assign \adder_32bit_0.operator_B_stage_2_12.G1 = \adder_32bit_0.operator_B_stage_1_11.Go ;
  assign \adder_32bit_0.operator_B_stage_2_12.P = \adder_32bit_0.operator_B_stage_1_12.Po ;
  assign \adder_32bit_0.operator_B_stage_2_12.P1 = \adder_32bit_0.operator_B_stage_1_11.Po ;
  assign \adder_32bit_0.operator_B_stage_2_13.G = \adder_32bit_0.operator_B_stage_1_13.Go ;
  assign \adder_32bit_0.operator_B_stage_2_13.G1 = \adder_32bit_0.operator_B_stage_1_12.Go ;
  assign \adder_32bit_0.operator_B_stage_2_13.P = \adder_32bit_0.operator_B_stage_1_13.Po ;
  assign \adder_32bit_0.operator_B_stage_2_13.P1 = \adder_32bit_0.operator_B_stage_1_12.Po ;
  assign \adder_32bit_0.operator_B_stage_2_14.G = \adder_32bit_0.operator_B_stage_1_14.Go ;
  assign \adder_32bit_0.operator_B_stage_2_14.G1 = \adder_32bit_0.operator_B_stage_1_13.Go ;
  assign \adder_32bit_0.operator_B_stage_2_14.P = \adder_32bit_0.operator_B_stage_1_14.Po ;
  assign \adder_32bit_0.operator_B_stage_2_14.P1 = \adder_32bit_0.operator_B_stage_1_13.Po ;
  assign \adder_32bit_0.operator_B_stage_2_15.G = \adder_32bit_0.operator_B_stage_1_15.Go ;
  assign \adder_32bit_0.operator_B_stage_2_15.G1 = \adder_32bit_0.operator_B_stage_1_14.Go ;
  assign \adder_32bit_0.operator_B_stage_2_15.P = \adder_32bit_0.operator_B_stage_1_15.Po ;
  assign \adder_32bit_0.operator_B_stage_2_15.P1 = \adder_32bit_0.operator_B_stage_1_14.Po ;
  assign \adder_32bit_0.operator_B_stage_2_2.G = \adder_32bit_0.operator_B_stage_1_2.Go ;
  assign \adder_32bit_0.operator_B_stage_2_2.G1 = \adder_32bit_0.operator_B_stage_1_1.Go ;
  assign \adder_32bit_0.operator_B_stage_2_2.P = \adder_32bit_0.operator_B_stage_1_2.Po ;
  assign \adder_32bit_0.operator_B_stage_2_2.P1 = \adder_32bit_0.operator_B_stage_1_1.Po ;
  assign \adder_32bit_0.operator_B_stage_2_3.G = \adder_32bit_0.operator_B_stage_1_3.Go ;
  assign \adder_32bit_0.operator_B_stage_2_3.G1 = \adder_32bit_0.operator_B_stage_1_2.Go ;
  assign \adder_32bit_0.operator_B_stage_2_3.P = \adder_32bit_0.operator_B_stage_1_3.Po ;
  assign \adder_32bit_0.operator_B_stage_2_3.P1 = \adder_32bit_0.operator_B_stage_1_2.Po ;
  assign \adder_32bit_0.operator_B_stage_2_4.G = \adder_32bit_0.operator_B_stage_1_4.Go ;
  assign \adder_32bit_0.operator_B_stage_2_4.G1 = \adder_32bit_0.operator_B_stage_1_3.Go ;
  assign \adder_32bit_0.operator_B_stage_2_4.P = \adder_32bit_0.operator_B_stage_1_4.Po ;
  assign \adder_32bit_0.operator_B_stage_2_4.P1 = \adder_32bit_0.operator_B_stage_1_3.Po ;
  assign \adder_32bit_0.operator_B_stage_2_5.G = \adder_32bit_0.operator_B_stage_1_5.Go ;
  assign \adder_32bit_0.operator_B_stage_2_5.G1 = \adder_32bit_0.operator_B_stage_1_4.Go ;
  assign \adder_32bit_0.operator_B_stage_2_5.P = \adder_32bit_0.operator_B_stage_1_5.Po ;
  assign \adder_32bit_0.operator_B_stage_2_5.P1 = \adder_32bit_0.operator_B_stage_1_4.Po ;
  assign \adder_32bit_0.operator_B_stage_2_6.G = \adder_32bit_0.operator_B_stage_1_6.Go ;
  assign \adder_32bit_0.operator_B_stage_2_6.G1 = \adder_32bit_0.operator_B_stage_1_5.Go ;
  assign \adder_32bit_0.operator_B_stage_2_6.P = \adder_32bit_0.operator_B_stage_1_6.Po ;
  assign \adder_32bit_0.operator_B_stage_2_6.P1 = \adder_32bit_0.operator_B_stage_1_5.Po ;
  assign \adder_32bit_0.operator_B_stage_2_7.G = \adder_32bit_0.operator_B_stage_1_7.Go ;
  assign \adder_32bit_0.operator_B_stage_2_7.G1 = \adder_32bit_0.operator_B_stage_1_6.Go ;
  assign \adder_32bit_0.operator_B_stage_2_7.P = \adder_32bit_0.operator_B_stage_1_7.Po ;
  assign \adder_32bit_0.operator_B_stage_2_7.P1 = \adder_32bit_0.operator_B_stage_1_6.Po ;
  assign \adder_32bit_0.operator_B_stage_2_8.G = \adder_32bit_0.operator_B_stage_1_8.Go ;
  assign \adder_32bit_0.operator_B_stage_2_8.G1 = \adder_32bit_0.operator_B_stage_1_7.Go ;
  assign \adder_32bit_0.operator_B_stage_2_8.P = \adder_32bit_0.operator_B_stage_1_8.Po ;
  assign \adder_32bit_0.operator_B_stage_2_8.P1 = \adder_32bit_0.operator_B_stage_1_7.Po ;
  assign \adder_32bit_0.operator_B_stage_2_9.G = \adder_32bit_0.operator_B_stage_1_9.Go ;
  assign \adder_32bit_0.operator_B_stage_2_9.G1 = \adder_32bit_0.operator_B_stage_1_8.Go ;
  assign \adder_32bit_0.operator_B_stage_2_9.P = \adder_32bit_0.operator_B_stage_1_9.Po ;
  assign \adder_32bit_0.operator_B_stage_2_9.P1 = \adder_32bit_0.operator_B_stage_1_8.Po ;
  assign \adder_32bit_0.operator_B_stage_3_10.G = \adder_32bit_0.operator_B_stage_2_10.Go ;
  assign \adder_32bit_0.operator_B_stage_3_10.G1 = \adder_32bit_0.operator_B_stage_2_8.Go ;
  assign \adder_32bit_0.operator_B_stage_3_10.P = \adder_32bit_0.operator_B_stage_2_10.Po ;
  assign \adder_32bit_0.operator_B_stage_3_10.P1 = \adder_32bit_0.operator_B_stage_2_8.Po ;
  assign \adder_32bit_0.operator_B_stage_3_11.G = \adder_32bit_0.operator_B_stage_2_11.Go ;
  assign \adder_32bit_0.operator_B_stage_3_11.G1 = \adder_32bit_0.operator_B_stage_2_9.Go ;
  assign \adder_32bit_0.operator_B_stage_3_11.P = \adder_32bit_0.operator_B_stage_2_11.Po ;
  assign \adder_32bit_0.operator_B_stage_3_11.P1 = \adder_32bit_0.operator_B_stage_2_9.Po ;
  assign \adder_32bit_0.operator_B_stage_3_12.G = \adder_32bit_0.operator_B_stage_2_12.Go ;
  assign \adder_32bit_0.operator_B_stage_3_12.G1 = \adder_32bit_0.operator_B_stage_2_10.Go ;
  assign \adder_32bit_0.operator_B_stage_3_12.P = \adder_32bit_0.operator_B_stage_2_12.Po ;
  assign \adder_32bit_0.operator_B_stage_3_12.P1 = \adder_32bit_0.operator_B_stage_2_10.Po ;
  assign \adder_32bit_0.operator_B_stage_3_13.G = \adder_32bit_0.operator_B_stage_2_13.Go ;
  assign \adder_32bit_0.operator_B_stage_3_13.G1 = \adder_32bit_0.operator_B_stage_2_11.Go ;
  assign \adder_32bit_0.operator_B_stage_3_13.P = \adder_32bit_0.operator_B_stage_2_13.Po ;
  assign \adder_32bit_0.operator_B_stage_3_13.P1 = \adder_32bit_0.operator_B_stage_2_11.Po ;
  assign \adder_32bit_0.operator_B_stage_3_14.G = \adder_32bit_0.operator_B_stage_2_14.Go ;
  assign \adder_32bit_0.operator_B_stage_3_14.G1 = \adder_32bit_0.operator_B_stage_2_12.Go ;
  assign \adder_32bit_0.operator_B_stage_3_14.P = \adder_32bit_0.operator_B_stage_2_14.Po ;
  assign \adder_32bit_0.operator_B_stage_3_14.P1 = \adder_32bit_0.operator_B_stage_2_12.Po ;
  assign \adder_32bit_0.operator_B_stage_3_15.G = \adder_32bit_0.operator_B_stage_2_15.Go ;
  assign \adder_32bit_0.operator_B_stage_3_15.G1 = \adder_32bit_0.operator_B_stage_2_13.Go ;
  assign \adder_32bit_0.operator_B_stage_3_15.P = \adder_32bit_0.operator_B_stage_2_15.Po ;
  assign \adder_32bit_0.operator_B_stage_3_15.P1 = \adder_32bit_0.operator_B_stage_2_13.Po ;
  assign \adder_32bit_0.operator_B_stage_3_4.G = \adder_32bit_0.operator_B_stage_2_4.Go ;
  assign \adder_32bit_0.operator_B_stage_3_4.G1 = \adder_32bit_0.operator_B_stage_2_2.Go ;
  assign \adder_32bit_0.operator_B_stage_3_4.P = \adder_32bit_0.operator_B_stage_2_4.Po ;
  assign \adder_32bit_0.operator_B_stage_3_4.P1 = \adder_32bit_0.operator_B_stage_2_2.Po ;
  assign \adder_32bit_0.operator_B_stage_3_5.G = \adder_32bit_0.operator_B_stage_2_5.Go ;
  assign \adder_32bit_0.operator_B_stage_3_5.G1 = \adder_32bit_0.operator_B_stage_2_3.Go ;
  assign \adder_32bit_0.operator_B_stage_3_5.P = \adder_32bit_0.operator_B_stage_2_5.Po ;
  assign \adder_32bit_0.operator_B_stage_3_5.P1 = \adder_32bit_0.operator_B_stage_2_3.Po ;
  assign \adder_32bit_0.operator_B_stage_3_6.G = \adder_32bit_0.operator_B_stage_2_6.Go ;
  assign \adder_32bit_0.operator_B_stage_3_6.G1 = \adder_32bit_0.operator_B_stage_2_4.Go ;
  assign \adder_32bit_0.operator_B_stage_3_6.P = \adder_32bit_0.operator_B_stage_2_6.Po ;
  assign \adder_32bit_0.operator_B_stage_3_6.P1 = \adder_32bit_0.operator_B_stage_2_4.Po ;
  assign \adder_32bit_0.operator_B_stage_3_7.G = \adder_32bit_0.operator_B_stage_2_7.Go ;
  assign \adder_32bit_0.operator_B_stage_3_7.G1 = \adder_32bit_0.operator_B_stage_2_5.Go ;
  assign \adder_32bit_0.operator_B_stage_3_7.P = \adder_32bit_0.operator_B_stage_2_7.Po ;
  assign \adder_32bit_0.operator_B_stage_3_7.P1 = \adder_32bit_0.operator_B_stage_2_5.Po ;
  assign \adder_32bit_0.operator_B_stage_3_8.G = \adder_32bit_0.operator_B_stage_2_8.Go ;
  assign \adder_32bit_0.operator_B_stage_3_8.G1 = \adder_32bit_0.operator_B_stage_2_6.Go ;
  assign \adder_32bit_0.operator_B_stage_3_8.P = \adder_32bit_0.operator_B_stage_2_8.Po ;
  assign \adder_32bit_0.operator_B_stage_3_8.P1 = \adder_32bit_0.operator_B_stage_2_6.Po ;
  assign \adder_32bit_0.operator_B_stage_3_9.G = \adder_32bit_0.operator_B_stage_2_9.Go ;
  assign \adder_32bit_0.operator_B_stage_3_9.G1 = \adder_32bit_0.operator_B_stage_2_7.Go ;
  assign \adder_32bit_0.operator_B_stage_3_9.P = \adder_32bit_0.operator_B_stage_2_9.Po ;
  assign \adder_32bit_0.operator_B_stage_3_9.P1 = \adder_32bit_0.operator_B_stage_2_7.Po ;
  assign \adder_32bit_0.operator_B_stage_4_10.G = \adder_32bit_0.operator_B_stage_3_10.Go ;
  assign \adder_32bit_0.operator_B_stage_4_10.G1 = \adder_32bit_0.operator_B_stage_3_6.Go ;
  assign \adder_32bit_0.operator_B_stage_4_10.P = \adder_32bit_0.operator_B_stage_3_10.Po ;
  assign \adder_32bit_0.operator_B_stage_4_10.P1 = \adder_32bit_0.operator_B_stage_3_6.Po ;
  assign \adder_32bit_0.operator_B_stage_4_11.G = \adder_32bit_0.operator_B_stage_3_11.Go ;
  assign \adder_32bit_0.operator_B_stage_4_11.G1 = \adder_32bit_0.operator_B_stage_3_7.Go ;
  assign \adder_32bit_0.operator_B_stage_4_11.P = \adder_32bit_0.operator_B_stage_3_11.Po ;
  assign \adder_32bit_0.operator_B_stage_4_11.P1 = \adder_32bit_0.operator_B_stage_3_7.Po ;
  assign \adder_32bit_0.operator_B_stage_4_12.G = \adder_32bit_0.operator_B_stage_3_12.Go ;
  assign \adder_32bit_0.operator_B_stage_4_12.G1 = \adder_32bit_0.operator_B_stage_3_8.Go ;
  assign \adder_32bit_0.operator_B_stage_4_12.P = \adder_32bit_0.operator_B_stage_3_12.Po ;
  assign \adder_32bit_0.operator_B_stage_4_12.P1 = \adder_32bit_0.operator_B_stage_3_8.Po ;
  assign \adder_32bit_0.operator_B_stage_4_13.G = \adder_32bit_0.operator_B_stage_3_13.Go ;
  assign \adder_32bit_0.operator_B_stage_4_13.G1 = \adder_32bit_0.operator_B_stage_3_9.Go ;
  assign \adder_32bit_0.operator_B_stage_4_13.P = \adder_32bit_0.operator_B_stage_3_13.Po ;
  assign \adder_32bit_0.operator_B_stage_4_13.P1 = \adder_32bit_0.operator_B_stage_3_9.Po ;
  assign \adder_32bit_0.operator_B_stage_4_14.G = \adder_32bit_0.operator_B_stage_3_14.Go ;
  assign \adder_32bit_0.operator_B_stage_4_14.G1 = \adder_32bit_0.operator_B_stage_3_10.Go ;
  assign \adder_32bit_0.operator_B_stage_4_14.P = \adder_32bit_0.operator_B_stage_3_14.Po ;
  assign \adder_32bit_0.operator_B_stage_4_14.P1 = \adder_32bit_0.operator_B_stage_3_10.Po ;
  assign \adder_32bit_0.operator_B_stage_4_15.G = \adder_32bit_0.operator_B_stage_3_15.Go ;
  assign \adder_32bit_0.operator_B_stage_4_15.G1 = \adder_32bit_0.operator_B_stage_3_11.Go ;
  assign \adder_32bit_0.operator_B_stage_4_15.P = \adder_32bit_0.operator_B_stage_3_15.Po ;
  assign \adder_32bit_0.operator_B_stage_4_15.P1 = \adder_32bit_0.operator_B_stage_3_11.Po ;
  assign \adder_32bit_0.operator_B_stage_4_8.G = \adder_32bit_0.operator_B_stage_3_8.Go ;
  assign \adder_32bit_0.operator_B_stage_4_8.G1 = \adder_32bit_0.operator_B_stage_3_4.Go ;
  assign \adder_32bit_0.operator_B_stage_4_8.P = \adder_32bit_0.operator_B_stage_3_8.Po ;
  assign \adder_32bit_0.operator_B_stage_4_8.P1 = \adder_32bit_0.operator_B_stage_3_4.Po ;
  assign \adder_32bit_0.operator_B_stage_4_9.G = \adder_32bit_0.operator_B_stage_3_9.Go ;
  assign \adder_32bit_0.operator_B_stage_4_9.G1 = \adder_32bit_0.operator_B_stage_3_5.Go ;
  assign \adder_32bit_0.operator_B_stage_4_9.P = \adder_32bit_0.operator_B_stage_3_9.Po ;
  assign \adder_32bit_0.operator_B_stage_4_9.P1 = \adder_32bit_0.operator_B_stage_3_5.Po ;
  assign \adder_32bit_0.operator_C_stage_1_0.G = \adder_32bit_0.operator_A_0.G ;
  assign \adder_32bit_0.operator_C_stage_1_0.G1 = cout;
  assign \adder_32bit_0.operator_C_stage_1_0.P = \adder_32bit_0.operator_A_0.P ;
  assign \adder_32bit_0.operator_C_stage_2_1.G = \adder_32bit_0.operator_B_stage_1_1.Go ;
  assign \adder_32bit_0.operator_C_stage_2_1.G1 = \adder_32bit_0.operator_C_stage_1_0.Go ;
  assign \adder_32bit_0.operator_C_stage_2_1.P = \adder_32bit_0.operator_B_stage_1_1.Po ;
  assign \adder_32bit_0.operator_C_stage_3_2.G = \adder_32bit_0.operator_B_stage_2_2.Go ;
  assign \adder_32bit_0.operator_C_stage_3_2.G1 = \adder_32bit_0.operator_C_stage_1_0.Go ;
  assign \adder_32bit_0.operator_C_stage_3_2.P = \adder_32bit_0.operator_B_stage_2_2.Po ;
  assign \adder_32bit_0.operator_C_stage_3_3.G = \adder_32bit_0.operator_B_stage_2_3.Go ;
  assign \adder_32bit_0.operator_C_stage_3_3.G1 = \adder_32bit_0.operator_C_stage_2_1.Go ;
  assign \adder_32bit_0.operator_C_stage_3_3.P = \adder_32bit_0.operator_B_stage_2_3.Po ;
  assign \adder_32bit_0.operator_C_stage_4_4.G = \adder_32bit_0.operator_B_stage_3_4.Go ;
  assign \adder_32bit_0.operator_C_stage_4_4.G1 = \adder_32bit_0.operator_C_stage_1_0.Go ;
  assign \adder_32bit_0.operator_C_stage_4_4.P = \adder_32bit_0.operator_B_stage_3_4.Po ;
  assign \adder_32bit_0.operator_C_stage_4_5.G = \adder_32bit_0.operator_B_stage_3_5.Go ;
  assign \adder_32bit_0.operator_C_stage_4_5.G1 = \adder_32bit_0.operator_C_stage_2_1.Go ;
  assign \adder_32bit_0.operator_C_stage_4_5.P = \adder_32bit_0.operator_B_stage_3_5.Po ;
  assign \adder_32bit_0.operator_C_stage_4_6.G = \adder_32bit_0.operator_B_stage_3_6.Go ;
  assign \adder_32bit_0.operator_C_stage_4_6.G1 = \adder_32bit_0.operator_C_stage_3_2.Go ;
  assign \adder_32bit_0.operator_C_stage_4_6.P = \adder_32bit_0.operator_B_stage_3_6.Po ;
  assign \adder_32bit_0.operator_C_stage_4_7.G = \adder_32bit_0.operator_B_stage_3_7.Go ;
  assign \adder_32bit_0.operator_C_stage_4_7.G1 = \adder_32bit_0.operator_C_stage_3_3.Go ;
  assign \adder_32bit_0.operator_C_stage_4_7.P = \adder_32bit_0.operator_B_stage_3_7.Po ;
  assign \adder_32bit_0.operator_C_stage_5_10.G = \adder_32bit_0.operator_B_stage_4_10.Go ;
  assign \adder_32bit_0.operator_C_stage_5_10.G1 = \adder_32bit_0.operator_C_stage_3_2.Go ;
  assign \adder_32bit_0.operator_C_stage_5_10.P = \adder_32bit_0.operator_B_stage_4_10.Po ;
  assign \adder_32bit_0.operator_C_stage_5_11.G = \adder_32bit_0.operator_B_stage_4_11.Go ;
  assign \adder_32bit_0.operator_C_stage_5_11.G1 = \adder_32bit_0.operator_C_stage_3_3.Go ;
  assign \adder_32bit_0.operator_C_stage_5_11.P = \adder_32bit_0.operator_B_stage_4_11.Po ;
  assign \adder_32bit_0.operator_C_stage_5_12.G = \adder_32bit_0.operator_B_stage_4_12.Go ;
  assign \adder_32bit_0.operator_C_stage_5_12.G1 = \adder_32bit_0.operator_C_stage_4_4.Go ;
  assign \adder_32bit_0.operator_C_stage_5_12.P = \adder_32bit_0.operator_B_stage_4_12.Po ;
  assign \adder_32bit_0.operator_C_stage_5_13.G = \adder_32bit_0.operator_B_stage_4_13.Go ;
  assign \adder_32bit_0.operator_C_stage_5_13.G1 = \adder_32bit_0.operator_C_stage_4_5.Go ;
  assign \adder_32bit_0.operator_C_stage_5_13.P = \adder_32bit_0.operator_B_stage_4_13.Po ;
  assign \adder_32bit_0.operator_C_stage_5_14.G = \adder_32bit_0.operator_B_stage_4_14.Go ;
  assign \adder_32bit_0.operator_C_stage_5_14.G1 = \adder_32bit_0.operator_C_stage_4_6.Go ;
  assign \adder_32bit_0.operator_C_stage_5_14.P = \adder_32bit_0.operator_B_stage_4_14.Po ;
  assign \adder_32bit_0.operator_C_stage_5_15.G = \adder_32bit_0.operator_B_stage_4_15.Go ;
  assign \adder_32bit_0.operator_C_stage_5_15.G1 = \adder_32bit_0.operator_C_stage_4_7.Go ;
  assign \adder_32bit_0.operator_C_stage_5_15.P = \adder_32bit_0.operator_B_stage_4_15.Po ;
  assign \adder_32bit_0.operator_C_stage_5_8.G = \adder_32bit_0.operator_B_stage_4_8.Go ;
  assign \adder_32bit_0.operator_C_stage_5_8.G1 = \adder_32bit_0.operator_C_stage_1_0.Go ;
  assign \adder_32bit_0.operator_C_stage_5_8.P = \adder_32bit_0.operator_B_stage_4_8.Po ;
  assign \adder_32bit_0.operator_C_stage_5_9.G = \adder_32bit_0.operator_B_stage_4_9.Go ;
  assign \adder_32bit_0.operator_C_stage_5_9.G1 = \adder_32bit_0.operator_C_stage_2_1.Go ;
  assign \adder_32bit_0.operator_C_stage_5_9.P = \adder_32bit_0.operator_B_stage_4_9.Po ;
  assign \adder_32bit_0.operator_C_stage_6_0.G = \adder_32bit_0.operator_A_1.G ;
  assign \adder_32bit_0.operator_C_stage_6_0.G1 = \adder_32bit_0.operator_C_stage_1_0.Go ;
  assign \adder_32bit_0.operator_C_stage_6_0.P = \adder_32bit_0.operator_A_1.P ;
  assign \adder_32bit_0.operator_C_stage_6_1.G = \adder_32bit_0.operator_A_3.G ;
  assign \adder_32bit_0.operator_C_stage_6_1.G1 = \adder_32bit_0.operator_C_stage_2_1.Go ;
  assign \adder_32bit_0.operator_C_stage_6_1.P = \adder_32bit_0.operator_A_3.P ;
  assign \adder_32bit_0.operator_C_stage_6_10.G = \adder_32bit_0.operator_A_21.G ;
  assign \adder_32bit_0.operator_C_stage_6_10.G1 = \adder_32bit_0.operator_C_stage_5_10.Go ;
  assign \adder_32bit_0.operator_C_stage_6_10.P = \adder_32bit_0.operator_A_21.P ;
  assign \adder_32bit_0.operator_C_stage_6_11.G = \adder_32bit_0.operator_A_23.G ;
  assign \adder_32bit_0.operator_C_stage_6_11.G1 = \adder_32bit_0.operator_C_stage_5_11.Go ;
  assign \adder_32bit_0.operator_C_stage_6_11.P = \adder_32bit_0.operator_A_23.P ;
  assign \adder_32bit_0.operator_C_stage_6_12.G = \adder_32bit_0.operator_A_25.G ;
  assign \adder_32bit_0.operator_C_stage_6_12.G1 = \adder_32bit_0.operator_C_stage_5_12.Go ;
  assign \adder_32bit_0.operator_C_stage_6_12.P = \adder_32bit_0.operator_A_25.P ;
  assign \adder_32bit_0.operator_C_stage_6_13.G = \adder_32bit_0.operator_A_27.G ;
  assign \adder_32bit_0.operator_C_stage_6_13.G1 = \adder_32bit_0.operator_C_stage_5_13.Go ;
  assign \adder_32bit_0.operator_C_stage_6_13.P = \adder_32bit_0.operator_A_27.P ;
  assign \adder_32bit_0.operator_C_stage_6_14.G = \adder_32bit_0.operator_A_29.G ;
  assign \adder_32bit_0.operator_C_stage_6_14.G1 = \adder_32bit_0.operator_C_stage_5_14.Go ;
  assign \adder_32bit_0.operator_C_stage_6_14.P = \adder_32bit_0.operator_A_29.P ;
  assign \adder_32bit_0.operator_C_stage_6_15.G1 = \adder_32bit_0.operator_C_stage_5_15.Go ;
  assign \adder_32bit_0.operator_C_stage_6_15.P = \adder_32bit_0.operator_A_31.P ;
  assign \adder_32bit_0.operator_C_stage_6_2.G = \adder_32bit_0.operator_A_5.G ;
  assign \adder_32bit_0.operator_C_stage_6_2.G1 = \adder_32bit_0.operator_C_stage_3_2.Go ;
  assign \adder_32bit_0.operator_C_stage_6_2.P = \adder_32bit_0.operator_A_5.P ;
  assign \adder_32bit_0.operator_C_stage_6_3.G = \adder_32bit_0.operator_A_7.G ;
  assign \adder_32bit_0.operator_C_stage_6_3.G1 = \adder_32bit_0.operator_C_stage_3_3.Go ;
  assign \adder_32bit_0.operator_C_stage_6_3.P = \adder_32bit_0.operator_A_7.P ;
  assign \adder_32bit_0.operator_C_stage_6_4.G = \adder_32bit_0.operator_A_9.G ;
  assign \adder_32bit_0.operator_C_stage_6_4.G1 = \adder_32bit_0.operator_C_stage_4_4.Go ;
  assign \adder_32bit_0.operator_C_stage_6_4.P = \adder_32bit_0.operator_A_9.P ;
  assign \adder_32bit_0.operator_C_stage_6_5.G = \adder_32bit_0.operator_A_11.G ;
  assign \adder_32bit_0.operator_C_stage_6_5.G1 = \adder_32bit_0.operator_C_stage_4_5.Go ;
  assign \adder_32bit_0.operator_C_stage_6_5.P = \adder_32bit_0.operator_A_11.P ;
  assign \adder_32bit_0.operator_C_stage_6_6.G = \adder_32bit_0.operator_A_13.G ;
  assign \adder_32bit_0.operator_C_stage_6_6.G1 = \adder_32bit_0.operator_C_stage_4_6.Go ;
  assign \adder_32bit_0.operator_C_stage_6_6.P = \adder_32bit_0.operator_A_13.P ;
  assign \adder_32bit_0.operator_C_stage_6_7.G = \adder_32bit_0.operator_A_15.G ;
  assign \adder_32bit_0.operator_C_stage_6_7.G1 = \adder_32bit_0.operator_C_stage_4_7.Go ;
  assign \adder_32bit_0.operator_C_stage_6_7.P = \adder_32bit_0.operator_A_15.P ;
  assign \adder_32bit_0.operator_C_stage_6_8.G = \adder_32bit_0.operator_A_17.G ;
  assign \adder_32bit_0.operator_C_stage_6_8.G1 = \adder_32bit_0.operator_C_stage_5_8.Go ;
  assign \adder_32bit_0.operator_C_stage_6_8.P = \adder_32bit_0.operator_A_17.P ;
  assign \adder_32bit_0.operator_C_stage_6_9.G = \adder_32bit_0.operator_A_19.G ;
  assign \adder_32bit_0.operator_C_stage_6_9.G1 = \adder_32bit_0.operator_C_stage_5_9.Go ;
  assign \adder_32bit_0.operator_C_stage_6_9.P = \adder_32bit_0.operator_A_19.P ;
  assign adr = i_wb_adr[4:2];
  assign adr_1 = i_wb_adr[5:2];
  assign \multiplier_16x16bit_pipelined.A = { \multiplier_16x16bit_pipelined.reg_layer_2_w31 , \multiplier_16x16bit_pipelined.adder_32bit.operator_A_30.A , \multiplier_16x16bit_pipelined.adder_32bit.operator_A_29.A , \multiplier_16x16bit_pipelined.adder_32bit.operator_A_28.A , \multiplier_16x16bit_pipelined.adder_32bit.operator_A_27.A , \multiplier_16x16bit_pipelined.adder_32bit.operator_A_26.A , \multiplier_16x16bit_pipelined.adder_32bit.operator_A_25.A , \multiplier_16x16bit_pipelined.adder_32bit.operator_A_24.A , \multiplier_16x16bit_pipelined.adder_32bit.operator_A_23.A , \multiplier_16x16bit_pipelined.adder_32bit.operator_A_22.A , \multiplier_16x16bit_pipelined.adder_32bit.operator_A_21.A , \multiplier_16x16bit_pipelined.adder_32bit.operator_A_20.A , \multiplier_16x16bit_pipelined.adder_32bit.operator_A_19.A , \multiplier_16x16bit_pipelined.adder_32bit.operator_A_18.A , \multiplier_16x16bit_pipelined.adder_32bit.operator_A_17.A , \multiplier_16x16bit_pipelined.adder_32bit.operator_A_16.A , \multiplier_16x16bit_pipelined.adder_32bit.operator_A_15.A , \multiplier_16x16bit_pipelined.adder_32bit.operator_A_14.A , \multiplier_16x16bit_pipelined.adder_32bit.operator_A_13.A , \multiplier_16x16bit_pipelined.adder_32bit.operator_A_12.A , \multiplier_16x16bit_pipelined.adder_32bit.operator_A_11.A , \multiplier_16x16bit_pipelined.adder_32bit.operator_A_10.A , \multiplier_16x16bit_pipelined.adder_32bit.operator_A_9.A , \multiplier_16x16bit_pipelined.adder_32bit.operator_A_8.A , \multiplier_16x16bit_pipelined.adder_32bit.operator_A_7.A , \multiplier_16x16bit_pipelined.adder_32bit.operator_A_6.A , \multiplier_16x16bit_pipelined.adder_32bit.operator_A_5.A , \multiplier_16x16bit_pipelined.adder_32bit.operator_A_4.A , \multiplier_16x16bit_pipelined.adder_32bit.operator_A_3.A , \multiplier_16x16bit_pipelined.adder_32bit.operator_A_2.A , \multiplier_16x16bit_pipelined.reg_layer_2_w1 , \multiplier_16x16bit_pipelined.reg_layer_2_w0 [0] };
  assign \multiplier_16x16bit_pipelined.B = { \multiplier_16x16bit_pipelined.reg_layer_2_w30 , 1'b0, \multiplier_16x16bit_pipelined.reg_layer_2_w28 , 1'b0, \multiplier_16x16bit_pipelined.adder_32bit.operator_A_26.B , 1'b0, \multiplier_16x16bit_pipelined.adder_32bit.operator_A_24.B , \multiplier_16x16bit_pipelined.adder_32bit.operator_A_23.B , \multiplier_16x16bit_pipelined.adder_32bit.operator_A_22.B , \multiplier_16x16bit_pipelined.adder_32bit.operator_A_21.B , \multiplier_16x16bit_pipelined.adder_32bit.operator_A_20.B , \multiplier_16x16bit_pipelined.adder_32bit.operator_A_19.B , \multiplier_16x16bit_pipelined.adder_32bit.operator_A_18.B , \multiplier_16x16bit_pipelined.adder_32bit.operator_A_17.B , \multiplier_16x16bit_pipelined.adder_32bit.operator_A_16.B , \multiplier_16x16bit_pipelined.adder_32bit.operator_A_15.B , \multiplier_16x16bit_pipelined.adder_32bit.operator_A_14.B , \multiplier_16x16bit_pipelined.adder_32bit.operator_A_13.B , \multiplier_16x16bit_pipelined.adder_32bit.operator_A_12.B , \multiplier_16x16bit_pipelined.adder_32bit.operator_A_11.B , \multiplier_16x16bit_pipelined.adder_32bit.operator_A_10.B , \multiplier_16x16bit_pipelined.adder_32bit.operator_A_9.B , \multiplier_16x16bit_pipelined.adder_32bit.operator_A_8.B , \multiplier_16x16bit_pipelined.adder_32bit.operator_A_7.B , \multiplier_16x16bit_pipelined.adder_32bit.operator_A_6.B , \multiplier_16x16bit_pipelined.adder_32bit.operator_A_5.B , \multiplier_16x16bit_pipelined.adder_32bit.operator_A_4.B , \multiplier_16x16bit_pipelined.adder_32bit.operator_A_3.B , 2'b00, \multiplier_16x16bit_pipelined.reg_layer_2_w0 [1] };
  assign \multiplier_16x16bit_pipelined.adder_32bit.G0 [30:0] = { \multiplier_16x16bit_pipelined.adder_32bit.operator_A_30.G , 1'b0, \multiplier_16x16bit_pipelined.adder_32bit.operator_A_28.G , 1'b0, \multiplier_16x16bit_pipelined.adder_32bit.operator_A_26.G , 1'b0, \multiplier_16x16bit_pipelined.adder_32bit.operator_A_24.G , \multiplier_16x16bit_pipelined.adder_32bit.operator_A_23.G , \multiplier_16x16bit_pipelined.adder_32bit.operator_A_22.G , \multiplier_16x16bit_pipelined.adder_32bit.operator_A_21.G , \multiplier_16x16bit_pipelined.adder_32bit.operator_A_20.G , \multiplier_16x16bit_pipelined.adder_32bit.operator_A_19.G , \multiplier_16x16bit_pipelined.adder_32bit.operator_A_18.G , \multiplier_16x16bit_pipelined.adder_32bit.operator_A_17.G , \multiplier_16x16bit_pipelined.adder_32bit.operator_A_16.G , \multiplier_16x16bit_pipelined.adder_32bit.operator_A_15.G , \multiplier_16x16bit_pipelined.adder_32bit.operator_A_14.G , \multiplier_16x16bit_pipelined.adder_32bit.operator_A_13.G , \multiplier_16x16bit_pipelined.adder_32bit.operator_A_12.G , \multiplier_16x16bit_pipelined.adder_32bit.operator_A_11.G , \multiplier_16x16bit_pipelined.adder_32bit.operator_A_10.G , \multiplier_16x16bit_pipelined.adder_32bit.operator_A_9.G , \multiplier_16x16bit_pipelined.adder_32bit.operator_A_8.G , \multiplier_16x16bit_pipelined.adder_32bit.operator_A_7.G , \multiplier_16x16bit_pipelined.adder_32bit.operator_A_6.G , \multiplier_16x16bit_pipelined.adder_32bit.operator_A_5.G , \multiplier_16x16bit_pipelined.adder_32bit.operator_A_4.G , \multiplier_16x16bit_pipelined.adder_32bit.operator_A_3.G , 2'b00, \multiplier_16x16bit_pipelined.adder_32bit.operator_A_0.G };
  assign \multiplier_16x16bit_pipelined.adder_32bit.G1 = { \multiplier_16x16bit_pipelined.adder_32bit.operator_A_30.G , \multiplier_16x16bit_pipelined.adder_32bit.operator_A_28.G , \multiplier_16x16bit_pipelined.adder_32bit.operator_A_26.G , \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_12.Go , \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_11.Go , \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_10.Go , \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_9.Go , \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_8.Go , \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_7.Go , \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_6.Go , \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_5.Go , \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_4.Go , \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_3.Go , \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_2.Go , 1'b0, \multiplier_16x16bit_pipelined.adder_32bit.operator_A_0.G };
  assign \multiplier_16x16bit_pipelined.adder_32bit.G2 = { \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_15.Go , \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_14.Go , \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_13.Go , \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_12.Go , \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_11.Go , \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_10.Go , \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_9.Go , \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_8.Go , \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_7.Go , \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_6.Go , \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_5.Go , \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_4.Go , \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_3.Go , \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_2.Go , \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_2_1.Go , \multiplier_16x16bit_pipelined.adder_32bit.operator_A_0.G };
  assign \multiplier_16x16bit_pipelined.adder_32bit.G3 = { \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_15.Go , \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_14.Go , \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_13.Go , \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_12.Go , \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_11.Go , \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_10.Go , \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_9.Go , \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_8.Go , \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_7.Go , \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_6.Go , \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_5.Go , \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_4.Go , \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_3_3.Go , \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_3_2.Go , \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_2_1.Go , \multiplier_16x16bit_pipelined.adder_32bit.operator_A_0.G };
  assign \multiplier_16x16bit_pipelined.adder_32bit.G4 = { \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_4_15.Go , \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_4_14.Go , \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_4_13.Go , \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_4_12.Go , \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_4_11.Go , \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_4_10.Go , \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_4_9.Go , \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_4_8.Go , \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_4_7.Go , \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_4_6.Go , \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_4_5.Go , \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_4_4.Go , \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_3_3.Go , \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_3_2.Go , \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_2_1.Go , \multiplier_16x16bit_pipelined.adder_32bit.operator_A_0.G };
  assign \multiplier_16x16bit_pipelined.adder_32bit.G5 = { \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_5_15.Go , \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_5_14.Go , \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_5_13.Go , \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_5_12.Go , \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_5_11.Go , \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_5_10.Go , \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_5_9.Go , \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_5_8.Go , \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_4_7.Go , \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_4_6.Go , \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_4_5.Go , \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_4_4.Go , \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_3_3.Go , \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_3_2.Go , \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_2_1.Go , \multiplier_16x16bit_pipelined.adder_32bit.operator_A_0.G };
  assign \multiplier_16x16bit_pipelined.adder_32bit.G6 [30:0] = { \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_5_15.Go , \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_6_14.Go , \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_5_14.Go , \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_6_13.Go , \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_5_13.Go , \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_6_12.Go , \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_5_12.Go , \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_6_11.Go , \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_5_11.Go , \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_6_10.Go , \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_5_10.Go , \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_6_9.Go , \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_5_9.Go , \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_6_8.Go , \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_5_8.Go , \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_6_7.Go , \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_4_7.Go , \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_6_6.Go , \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_4_6.Go , \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_6_5.Go , \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_4_5.Go , \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_6_4.Go , \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_4_4.Go , \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_6_3.Go , \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_3_3.Go , \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_6_2.Go , \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_3_2.Go , \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_6_1.Go , \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_2_1.Go , \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_6_0.Go , \multiplier_16x16bit_pipelined.adder_32bit.operator_A_0.G };
  assign \multiplier_16x16bit_pipelined.adder_32bit.P0 = { \multiplier_16x16bit_pipelined.reg_layer_2_w31 , \multiplier_16x16bit_pipelined.adder_32bit.operator_A_30.P , \multiplier_16x16bit_pipelined.adder_32bit.operator_A_29.A , \multiplier_16x16bit_pipelined.adder_32bit.operator_A_28.P , \multiplier_16x16bit_pipelined.adder_32bit.operator_A_27.A , \multiplier_16x16bit_pipelined.adder_32bit.operator_A_26.P , \multiplier_16x16bit_pipelined.adder_32bit.operator_A_25.A , \multiplier_16x16bit_pipelined.adder_32bit.operator_A_24.P , \multiplier_16x16bit_pipelined.adder_32bit.operator_A_23.P , \multiplier_16x16bit_pipelined.adder_32bit.operator_A_22.P , \multiplier_16x16bit_pipelined.adder_32bit.operator_A_21.P , \multiplier_16x16bit_pipelined.adder_32bit.operator_A_20.P , \multiplier_16x16bit_pipelined.adder_32bit.operator_A_19.P , \multiplier_16x16bit_pipelined.adder_32bit.operator_A_18.P , \multiplier_16x16bit_pipelined.adder_32bit.operator_A_17.P , \multiplier_16x16bit_pipelined.adder_32bit.operator_A_16.P , \multiplier_16x16bit_pipelined.adder_32bit.operator_A_15.P , \multiplier_16x16bit_pipelined.adder_32bit.operator_A_14.P , \multiplier_16x16bit_pipelined.adder_32bit.operator_A_13.P , \multiplier_16x16bit_pipelined.adder_32bit.operator_A_12.P , \multiplier_16x16bit_pipelined.adder_32bit.operator_A_11.P , \multiplier_16x16bit_pipelined.adder_32bit.operator_A_10.P , \multiplier_16x16bit_pipelined.adder_32bit.operator_A_9.P , \multiplier_16x16bit_pipelined.adder_32bit.operator_A_8.P , \multiplier_16x16bit_pipelined.adder_32bit.operator_A_7.P , \multiplier_16x16bit_pipelined.adder_32bit.operator_A_6.P , \multiplier_16x16bit_pipelined.adder_32bit.operator_A_5.P , \multiplier_16x16bit_pipelined.adder_32bit.operator_A_4.P , \multiplier_16x16bit_pipelined.adder_32bit.operator_A_3.P , \multiplier_16x16bit_pipelined.adder_32bit.operator_A_2.A , \multiplier_16x16bit_pipelined.reg_layer_2_w1 , \multiplier_16x16bit_pipelined.adder_32bit.operator_A_0.P };
  assign \multiplier_16x16bit_pipelined.adder_32bit.P1 = { \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_15.Po , \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_14.Po , \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_13.Po , \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_12.Po , \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_11.Po , \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_10.Po , \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_9.Po , \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_8.Po , \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_7.Po , \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_6.Po , \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_5.Po , \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_4.Po , \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_3.Po , \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_2.Po , \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_1.Po };
  assign \multiplier_16x16bit_pipelined.adder_32bit.P2 = { \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_15.Po , \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_14.Po , \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_13.Po , \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_12.Po , \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_11.Po , \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_10.Po , \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_9.Po , \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_8.Po , \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_7.Po , \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_6.Po , \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_5.Po , \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_4.Po , \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_3.Po , \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_2.Po };
  assign \multiplier_16x16bit_pipelined.adder_32bit.P3 = { \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_15.Po , \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_14.Po , \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_13.Po , \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_12.Po , \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_11.Po , \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_10.Po , \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_9.Po , \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_8.Po , \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_7.Po , \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_6.Po , \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_5.Po , \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_4.Po };
  assign \multiplier_16x16bit_pipelined.adder_32bit.P4 = { \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_4_15.Po , \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_4_14.Po , \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_4_13.Po , \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_4_12.Po , \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_4_11.Po , \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_4_10.Po , \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_4_9.Po , \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_4_8.Po };
  assign \multiplier_16x16bit_pipelined.adder_32bit.i_a = { \multiplier_16x16bit_pipelined.reg_layer_2_w31 , \multiplier_16x16bit_pipelined.adder_32bit.operator_A_30.A , \multiplier_16x16bit_pipelined.adder_32bit.operator_A_29.A , \multiplier_16x16bit_pipelined.adder_32bit.operator_A_28.A , \multiplier_16x16bit_pipelined.adder_32bit.operator_A_27.A , \multiplier_16x16bit_pipelined.adder_32bit.operator_A_26.A , \multiplier_16x16bit_pipelined.adder_32bit.operator_A_25.A , \multiplier_16x16bit_pipelined.adder_32bit.operator_A_24.A , \multiplier_16x16bit_pipelined.adder_32bit.operator_A_23.A , \multiplier_16x16bit_pipelined.adder_32bit.operator_A_22.A , \multiplier_16x16bit_pipelined.adder_32bit.operator_A_21.A , \multiplier_16x16bit_pipelined.adder_32bit.operator_A_20.A , \multiplier_16x16bit_pipelined.adder_32bit.operator_A_19.A , \multiplier_16x16bit_pipelined.adder_32bit.operator_A_18.A , \multiplier_16x16bit_pipelined.adder_32bit.operator_A_17.A , \multiplier_16x16bit_pipelined.adder_32bit.operator_A_16.A , \multiplier_16x16bit_pipelined.adder_32bit.operator_A_15.A , \multiplier_16x16bit_pipelined.adder_32bit.operator_A_14.A , \multiplier_16x16bit_pipelined.adder_32bit.operator_A_13.A , \multiplier_16x16bit_pipelined.adder_32bit.operator_A_12.A , \multiplier_16x16bit_pipelined.adder_32bit.operator_A_11.A , \multiplier_16x16bit_pipelined.adder_32bit.operator_A_10.A , \multiplier_16x16bit_pipelined.adder_32bit.operator_A_9.A , \multiplier_16x16bit_pipelined.adder_32bit.operator_A_8.A , \multiplier_16x16bit_pipelined.adder_32bit.operator_A_7.A , \multiplier_16x16bit_pipelined.adder_32bit.operator_A_6.A , \multiplier_16x16bit_pipelined.adder_32bit.operator_A_5.A , \multiplier_16x16bit_pipelined.adder_32bit.operator_A_4.A , \multiplier_16x16bit_pipelined.adder_32bit.operator_A_3.A , \multiplier_16x16bit_pipelined.adder_32bit.operator_A_2.A , \multiplier_16x16bit_pipelined.reg_layer_2_w1 , \multiplier_16x16bit_pipelined.reg_layer_2_w0 [0] };
  assign \multiplier_16x16bit_pipelined.adder_32bit.i_b = { 1'b0, \multiplier_16x16bit_pipelined.reg_layer_2_w30 , 1'b0, \multiplier_16x16bit_pipelined.reg_layer_2_w28 , 1'b0, \multiplier_16x16bit_pipelined.adder_32bit.operator_A_26.B , 1'b0, \multiplier_16x16bit_pipelined.adder_32bit.operator_A_24.B , \multiplier_16x16bit_pipelined.adder_32bit.operator_A_23.B , \multiplier_16x16bit_pipelined.adder_32bit.operator_A_22.B , \multiplier_16x16bit_pipelined.adder_32bit.operator_A_21.B , \multiplier_16x16bit_pipelined.adder_32bit.operator_A_20.B , \multiplier_16x16bit_pipelined.adder_32bit.operator_A_19.B , \multiplier_16x16bit_pipelined.adder_32bit.operator_A_18.B , \multiplier_16x16bit_pipelined.adder_32bit.operator_A_17.B , \multiplier_16x16bit_pipelined.adder_32bit.operator_A_16.B , \multiplier_16x16bit_pipelined.adder_32bit.operator_A_15.B , \multiplier_16x16bit_pipelined.adder_32bit.operator_A_14.B , \multiplier_16x16bit_pipelined.adder_32bit.operator_A_13.B , \multiplier_16x16bit_pipelined.adder_32bit.operator_A_12.B , \multiplier_16x16bit_pipelined.adder_32bit.operator_A_11.B , \multiplier_16x16bit_pipelined.adder_32bit.operator_A_10.B , \multiplier_16x16bit_pipelined.adder_32bit.operator_A_9.B , \multiplier_16x16bit_pipelined.adder_32bit.operator_A_8.B , \multiplier_16x16bit_pipelined.adder_32bit.operator_A_7.B , \multiplier_16x16bit_pipelined.adder_32bit.operator_A_6.B , \multiplier_16x16bit_pipelined.adder_32bit.operator_A_5.B , \multiplier_16x16bit_pipelined.adder_32bit.operator_A_4.B , \multiplier_16x16bit_pipelined.adder_32bit.operator_A_3.B , 2'b00, \multiplier_16x16bit_pipelined.reg_layer_2_w0 [1] };
  assign \multiplier_16x16bit_pipelined.adder_32bit.o_s [0] = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_0.P ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_A_0.A = \multiplier_16x16bit_pipelined.reg_layer_2_w0 [0];
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_A_0.B = \multiplier_16x16bit_pipelined.reg_layer_2_w0 [1];
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_A_1.A = \multiplier_16x16bit_pipelined.reg_layer_2_w1 ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_A_1.P = \multiplier_16x16bit_pipelined.reg_layer_2_w1 ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_A_2.P = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_2.A ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_A_25.P = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_25.A ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_A_27.P = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_27.A ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_A_28.B = \multiplier_16x16bit_pipelined.reg_layer_2_w28 ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_A_29.P = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_29.A ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_A_30.B = \multiplier_16x16bit_pipelined.reg_layer_2_w30 ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_A_31.A = \multiplier_16x16bit_pipelined.reg_layer_2_w31 ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_A_31.P = \multiplier_16x16bit_pipelined.reg_layer_2_w31 ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_1.P = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_2.A ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_1.P1 = \multiplier_16x16bit_pipelined.reg_layer_2_w1 ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_10.G = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_20.G ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_10.G1 = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_19.G ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_10.P = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_20.P ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_10.P1 = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_19.P ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_11.G = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_22.G ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_11.G1 = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_21.G ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_11.P = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_22.P ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_11.P1 = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_21.P ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_12.G = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_24.G ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_12.G1 = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_23.G ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_12.P = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_24.P ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_12.P1 = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_23.P ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_13.G = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_26.G ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_13.Go = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_26.G ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_13.P = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_26.P ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_13.P1 = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_25.A ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_14.G = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_28.G ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_14.Go = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_28.G ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_14.P = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_28.P ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_14.P1 = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_27.A ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_15.G = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_30.G ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_15.Go = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_30.G ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_15.P = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_30.P ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_15.P1 = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_29.A ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_2.G = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_4.G ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_2.G1 = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_3.G ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_2.P = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_4.P ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_2.P1 = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_3.P ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_3.G = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_6.G ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_3.G1 = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_5.G ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_3.P = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_6.P ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_3.P1 = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_5.P ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_4.G = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_8.G ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_4.G1 = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_7.G ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_4.P = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_8.P ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_4.P1 = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_7.P ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_5.G = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_10.G ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_5.G1 = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_9.G ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_5.P = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_10.P ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_5.P1 = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_9.P ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_6.G = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_12.G ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_6.G1 = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_11.G ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_6.P = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_12.P ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_6.P1 = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_11.P ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_7.G = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_14.G ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_7.G1 = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_13.G ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_7.P = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_14.P ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_7.P1 = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_13.P ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_8.G = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_16.G ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_8.G1 = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_15.G ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_8.P = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_16.P ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_8.P1 = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_15.P ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_9.G = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_18.G ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_9.G1 = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_17.G ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_9.P = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_18.P ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_9.P1 = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_17.P ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_10.G = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_10.Go ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_10.G1 = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_9.Go ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_10.P = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_10.Po ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_10.P1 = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_9.Po ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_11.G = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_11.Go ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_11.G1 = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_10.Go ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_11.P = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_11.Po ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_11.P1 = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_10.Po ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_12.G = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_12.Go ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_12.G1 = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_11.Go ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_12.P = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_12.Po ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_12.P1 = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_11.Po ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_13.G = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_26.G ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_13.G1 = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_12.Go ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_13.P = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_13.Po ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_13.P1 = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_12.Po ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_14.G = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_28.G ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_14.G1 = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_26.G ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_14.P = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_14.Po ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_14.P1 = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_13.Po ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_15.G = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_30.G ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_15.G1 = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_28.G ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_15.P = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_15.Po ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_15.P1 = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_14.Po ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_2.G = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_2.Go ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_2.Go = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_2.Go ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_2.P = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_2.Po ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_2.P1 = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_1.Po ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_3.G = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_3.Go ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_3.G1 = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_2.Go ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_3.P = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_3.Po ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_3.P1 = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_2.Po ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_4.G = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_4.Go ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_4.G1 = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_3.Go ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_4.P = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_4.Po ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_4.P1 = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_3.Po ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_5.G = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_5.Go ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_5.G1 = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_4.Go ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_5.P = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_5.Po ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_5.P1 = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_4.Po ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_6.G = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_6.Go ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_6.G1 = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_5.Go ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_6.P = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_6.Po ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_6.P1 = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_5.Po ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_7.G = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_7.Go ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_7.G1 = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_6.Go ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_7.P = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_7.Po ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_7.P1 = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_6.Po ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_8.G = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_8.Go ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_8.G1 = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_7.Go ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_8.P = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_8.Po ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_8.P1 = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_7.Po ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_9.G = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_9.Go ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_9.G1 = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_8.Go ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_9.P = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_9.Po ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_9.P1 = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_8.Po ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_10.G = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_10.Go ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_10.G1 = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_8.Go ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_10.P = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_10.Po ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_10.P1 = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_8.Po ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_11.G = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_11.Go ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_11.G1 = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_9.Go ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_11.P = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_11.Po ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_11.P1 = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_9.Po ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_12.G = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_12.Go ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_12.G1 = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_10.Go ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_12.P = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_12.Po ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_12.P1 = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_10.Po ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_13.G = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_13.Go ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_13.G1 = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_11.Go ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_13.P = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_13.Po ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_13.P1 = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_11.Po ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_14.G = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_14.Go ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_14.G1 = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_12.Go ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_14.P = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_14.Po ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_14.P1 = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_12.Po ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_15.G = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_15.Go ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_15.G1 = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_13.Go ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_15.P = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_15.Po ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_15.P1 = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_13.Po ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_4.G = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_4.Go ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_4.G1 = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_2.Go ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_4.P = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_4.Po ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_4.P1 = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_2.Po ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_5.G = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_5.Go ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_5.G1 = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_3.Go ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_5.P = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_5.Po ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_5.P1 = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_3.Po ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_6.G = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_6.Go ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_6.G1 = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_4.Go ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_6.P = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_6.Po ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_6.P1 = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_4.Po ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_7.G = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_7.Go ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_7.G1 = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_5.Go ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_7.P = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_7.Po ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_7.P1 = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_5.Po ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_8.G = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_8.Go ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_8.G1 = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_6.Go ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_8.P = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_8.Po ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_8.P1 = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_6.Po ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_9.G = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_9.Go ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_9.G1 = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_7.Go ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_9.P = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_9.Po ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_9.P1 = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_7.Po ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_4_10.G = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_10.Go ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_4_10.G1 = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_6.Go ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_4_10.P = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_10.Po ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_4_10.P1 = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_6.Po ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_4_11.G = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_11.Go ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_4_11.G1 = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_7.Go ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_4_11.P = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_11.Po ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_4_11.P1 = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_7.Po ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_4_12.G = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_12.Go ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_4_12.G1 = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_8.Go ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_4_12.P = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_12.Po ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_4_12.P1 = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_8.Po ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_4_13.G = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_13.Go ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_4_13.G1 = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_9.Go ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_4_13.P = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_13.Po ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_4_13.P1 = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_9.Po ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_4_14.G = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_14.Go ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_4_14.G1 = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_10.Go ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_4_14.P = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_14.Po ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_4_14.P1 = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_10.Po ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_4_15.G = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_15.Go ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_4_15.G1 = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_11.Go ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_4_15.P = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_15.Po ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_4_15.P1 = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_11.Po ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_4_8.G = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_8.Go ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_4_8.G1 = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_4.Go ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_4_8.P = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_8.Po ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_4_8.P1 = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_4.Po ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_4_9.G = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_9.Go ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_4_9.G1 = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_5.Go ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_4_9.P = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_9.Po ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_4_9.P1 = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_5.Po ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_1_0.G = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_0.G ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_1_0.Go = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_0.G ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_1_0.P = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_0.P ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_2_1.G1 = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_0.G ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_2_1.P = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_1.Po ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_3_2.G = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_1_2.Go ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_3_2.G1 = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_0.G ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_3_2.P = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_2.Po ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_3_3.G = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_3.Go ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_3_3.G1 = \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_2_1.Go ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_3_3.P = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_2_3.Po ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_4_4.G = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_4.Go ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_4_4.G1 = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_0.G ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_4_4.P = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_4.Po ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_4_5.G = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_5.Go ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_4_5.G1 = \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_2_1.Go ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_4_5.P = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_5.Po ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_4_6.G = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_6.Go ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_4_6.G1 = \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_3_2.Go ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_4_6.P = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_6.Po ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_4_7.G = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_7.Go ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_4_7.G1 = \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_3_3.Go ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_4_7.P = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_3_7.Po ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_5_10.G = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_4_10.Go ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_5_10.G1 = \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_3_2.Go ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_5_10.P = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_4_10.Po ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_5_11.G = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_4_11.Go ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_5_11.G1 = \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_3_3.Go ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_5_11.P = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_4_11.Po ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_5_12.G = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_4_12.Go ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_5_12.G1 = \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_4_4.Go ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_5_12.P = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_4_12.Po ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_5_13.G = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_4_13.Go ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_5_13.G1 = \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_4_5.Go ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_5_13.P = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_4_13.Po ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_5_14.G = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_4_14.Go ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_5_14.G1 = \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_4_6.Go ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_5_14.P = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_4_14.Po ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_5_15.G = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_4_15.Go ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_5_15.G1 = \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_4_7.Go ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_5_15.P = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_4_15.Po ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_5_8.G = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_4_8.Go ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_5_8.G1 = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_0.G ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_5_8.P = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_4_8.Po ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_5_9.G = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_4_9.Go ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_5_9.G1 = \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_2_1.Go ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_5_9.P = \multiplier_16x16bit_pipelined.adder_32bit.operator_B_stage_4_9.Po ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_6_0.G1 = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_0.G ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_6_0.P = \multiplier_16x16bit_pipelined.reg_layer_2_w1 ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_6_1.G = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_3.G ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_6_1.G1 = \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_2_1.Go ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_6_1.P = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_3.P ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_6_10.G = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_21.G ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_6_10.G1 = \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_5_10.Go ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_6_10.P = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_21.P ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_6_11.G = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_23.G ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_6_11.G1 = \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_5_11.Go ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_6_11.P = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_23.P ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_6_12.G1 = \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_5_12.Go ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_6_12.P = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_25.A ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_6_13.G1 = \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_5_13.Go ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_6_13.P = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_27.A ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_6_14.G1 = \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_5_14.Go ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_6_14.P = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_29.A ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_6_15.G1 = \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_5_15.Go ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_6_15.P = \multiplier_16x16bit_pipelined.reg_layer_2_w31 ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_6_2.G = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_5.G ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_6_2.G1 = \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_3_2.Go ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_6_2.P = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_5.P ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_6_3.G = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_7.G ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_6_3.G1 = \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_3_3.Go ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_6_3.P = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_7.P ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_6_4.G = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_9.G ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_6_4.G1 = \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_4_4.Go ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_6_4.P = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_9.P ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_6_5.G = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_11.G ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_6_5.G1 = \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_4_5.Go ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_6_5.P = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_11.P ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_6_6.G = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_13.G ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_6_6.G1 = \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_4_6.Go ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_6_6.P = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_13.P ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_6_7.G = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_15.G ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_6_7.G1 = \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_4_7.Go ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_6_7.P = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_15.P ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_6_8.G = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_17.G ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_6_8.G1 = \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_5_8.Go ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_6_8.P = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_17.P ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_6_9.G = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_19.G ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_6_9.G1 = \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_5_9.Go ;
  assign \multiplier_16x16bit_pipelined.adder_32bit.operator_C_stage_6_9.P = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_19.P ;
  assign \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_0.A = \multiplier_16x16bit_pipelined.mr [1];
  assign \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_0.B = \multiplier_16x16bit_pipelined.mr [0];
  assign \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_0.codes = { \multiplier_16x16bit_pipelined.mr [1:0], 1'b0 };
  assign \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_0.nBnC = \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_0.nB ;
  assign \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_0.negation = \multiplier_16x16bit_pipelined.mr [1];
  assign \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_1.A = \multiplier_16x16bit_pipelined.mr [3];
  assign \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_1.B = \multiplier_16x16bit_pipelined.mr [2];
  assign \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_1.C = \multiplier_16x16bit_pipelined.mr [1];
  assign \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_1.codes = \multiplier_16x16bit_pipelined.mr [3:1];
  assign \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_1.nC = \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_0.nA ;
  assign \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_2.A = \multiplier_16x16bit_pipelined.mr [5];
  assign \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_2.B = \multiplier_16x16bit_pipelined.mr [4];
  assign \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_2.C = \multiplier_16x16bit_pipelined.mr [3];
  assign \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_2.codes = \multiplier_16x16bit_pipelined.mr [5:3];
  assign \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_2.nC = \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_1.nA ;
  assign \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_3.A = \multiplier_16x16bit_pipelined.mr [7];
  assign \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_3.B = \multiplier_16x16bit_pipelined.mr [6];
  assign \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_3.C = \multiplier_16x16bit_pipelined.mr [5];
  assign \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_3.codes = \multiplier_16x16bit_pipelined.mr [7:5];
  assign \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_3.nC = \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_2.nA ;
  assign \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_4.A = \multiplier_16x16bit_pipelined.mr [9];
  assign \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_4.B = \multiplier_16x16bit_pipelined.mr [8];
  assign \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_4.C = \multiplier_16x16bit_pipelined.mr [7];
  assign \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_4.codes = \multiplier_16x16bit_pipelined.mr [9:7];
  assign \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_4.nC = \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_3.nA ;
  assign \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_5.A = \multiplier_16x16bit_pipelined.mr [11];
  assign \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_5.B = \multiplier_16x16bit_pipelined.mr [10];
  assign \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_5.C = \multiplier_16x16bit_pipelined.mr [9];
  assign \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_5.codes = \multiplier_16x16bit_pipelined.mr [11:9];
  assign \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_5.nC = \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_4.nA ;
  assign \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_6.A = \multiplier_16x16bit_pipelined.mr [13];
  assign \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_6.B = \multiplier_16x16bit_pipelined.mr [12];
  assign \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_6.C = \multiplier_16x16bit_pipelined.mr [11];
  assign \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_6.codes = \multiplier_16x16bit_pipelined.mr [13:11];
  assign \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_6.nC = \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_5.nA ;
  assign \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_7.A = \multiplier_16x16bit_pipelined.mr [15];
  assign \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_7.B = \multiplier_16x16bit_pipelined.mr [14];
  assign \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_7.C = \multiplier_16x16bit_pipelined.mr [13];
  assign \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_7.codes = \multiplier_16x16bit_pipelined.mr [15:13];
  assign \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_7.nC = \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_6.nA ;
  assign \multiplier_16x16bit_pipelined.booth_array_0.double = { \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_7.double , \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_6.double , \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_5.double , \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_4.double , \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_3.double , \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_2.double , \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_1.double , \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_0.double };
  assign \multiplier_16x16bit_pipelined.booth_array_0.multiplier = \multiplier_16x16bit_pipelined.mr ;
  assign \multiplier_16x16bit_pipelined.booth_array_0.negation = { \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_7.negation , \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_6.negation , \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_5.negation , \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_4.negation , \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_3.negation , \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_2.negation , \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_1.negation , \multiplier_16x16bit_pipelined.mr [1] };
  assign \multiplier_16x16bit_pipelined.booth_array_0.zero = { \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_7.zero , \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_6.zero , \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_5.zero , \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_4.zero , \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_3.zero , \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_2.zero , \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_1.zero , \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_0.zero };
  assign \multiplier_16x16bit_pipelined.double = { \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_7.double , \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_6.double , \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_5.double , \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_4.double , \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_3.double , \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_2.double , \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_1.double , \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_0.double };
  assign \multiplier_16x16bit_pipelined.i_clk = i_clk;
  assign \multiplier_16x16bit_pipelined.i_md = md;
  assign \multiplier_16x16bit_pipelined.i_mr = mr;
  assign \multiplier_16x16bit_pipelined.i_start = start;
  assign \multiplier_16x16bit_pipelined.layer_0_w0[1] = \multiplier_16x16bit_pipelined.mr [1];
  assign \multiplier_16x16bit_pipelined.layer_0_w10[0] = \multiplier_16x16bit_pipelined.layer_1_compressor42_3.A ;
  assign \multiplier_16x16bit_pipelined.layer_0_w10[1] = \multiplier_16x16bit_pipelined.layer_1_compressor42_3.B ;
  assign \multiplier_16x16bit_pipelined.layer_0_w10[2] = \multiplier_16x16bit_pipelined.layer_1_compressor42_3.C ;
  assign \multiplier_16x16bit_pipelined.layer_0_w10[3] = \multiplier_16x16bit_pipelined.layer_1_compressor42_3.D ;
  assign \multiplier_16x16bit_pipelined.layer_0_w10[4] = \multiplier_16x16bit_pipelined.layer_1_compressor42_3.cin ;
  assign \multiplier_16x16bit_pipelined.layer_0_w10[5] = \multiplier_16x16bit_pipelined.layer_2_compressor42_0.D ;
  assign \multiplier_16x16bit_pipelined.layer_0_w10[6] = \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_5.negation ;
  assign \multiplier_16x16bit_pipelined.layer_0_w11[0] = \multiplier_16x16bit_pipelined.layer_1_compressor42_4.A ;
  assign \multiplier_16x16bit_pipelined.layer_0_w11[1] = \multiplier_16x16bit_pipelined.layer_1_compressor42_4.B ;
  assign \multiplier_16x16bit_pipelined.layer_0_w11[2] = \multiplier_16x16bit_pipelined.layer_1_compressor42_4.C ;
  assign \multiplier_16x16bit_pipelined.layer_0_w11[3] = \multiplier_16x16bit_pipelined.layer_1_compressor42_4.D ;
  assign \multiplier_16x16bit_pipelined.layer_0_w11[4] = \multiplier_16x16bit_pipelined.layer_1_compressor42_4.cin ;
  assign \multiplier_16x16bit_pipelined.layer_0_w12[0] = \multiplier_16x16bit_pipelined.layer_1_compressor42_5.A ;
  assign \multiplier_16x16bit_pipelined.layer_0_w12[1] = \multiplier_16x16bit_pipelined.layer_1_compressor42_5.B ;
  assign \multiplier_16x16bit_pipelined.layer_0_w12[2] = \multiplier_16x16bit_pipelined.layer_1_compressor42_5.C ;
  assign \multiplier_16x16bit_pipelined.layer_0_w12[3] = \multiplier_16x16bit_pipelined.layer_1_compressor42_5.D ;
  assign \multiplier_16x16bit_pipelined.layer_0_w12[4] = \multiplier_16x16bit_pipelined.layer_1_compressor42_5.cin ;
  assign \multiplier_16x16bit_pipelined.layer_0_w12[5] = \multiplier_16x16bit_pipelined.layer_1_full_adder_3.A ;
  assign \multiplier_16x16bit_pipelined.layer_0_w12[6] = \multiplier_16x16bit_pipelined.layer_1_full_adder_3.B ;
  assign \multiplier_16x16bit_pipelined.layer_0_w12[7] = \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_6.negation ;
  assign \multiplier_16x16bit_pipelined.layer_0_w13[0] = \multiplier_16x16bit_pipelined.layer_1_compressor42_6.A ;
  assign \multiplier_16x16bit_pipelined.layer_0_w13[1] = \multiplier_16x16bit_pipelined.layer_1_compressor42_6.B ;
  assign \multiplier_16x16bit_pipelined.layer_0_w13[2] = \multiplier_16x16bit_pipelined.layer_1_compressor42_6.C ;
  assign \multiplier_16x16bit_pipelined.layer_0_w13[3] = \multiplier_16x16bit_pipelined.layer_1_compressor42_6.D ;
  assign \multiplier_16x16bit_pipelined.layer_0_w13[4] = \multiplier_16x16bit_pipelined.layer_1_compressor42_6.cin ;
  assign \multiplier_16x16bit_pipelined.layer_0_w13[5] = \multiplier_16x16bit_pipelined.layer_2_compressor42_1.cin ;
  assign \multiplier_16x16bit_pipelined.layer_0_w14[0] = \multiplier_16x16bit_pipelined.layer_1_compressor42_7.A ;
  assign \multiplier_16x16bit_pipelined.layer_0_w14[1] = \multiplier_16x16bit_pipelined.layer_1_compressor42_7.B ;
  assign \multiplier_16x16bit_pipelined.layer_0_w14[2] = \multiplier_16x16bit_pipelined.layer_1_compressor42_7.C ;
  assign \multiplier_16x16bit_pipelined.layer_0_w14[3] = \multiplier_16x16bit_pipelined.layer_1_compressor42_7.D ;
  assign \multiplier_16x16bit_pipelined.layer_0_w14[4] = \multiplier_16x16bit_pipelined.layer_1_compressor42_7.cin ;
  assign \multiplier_16x16bit_pipelined.layer_0_w14[5] = \multiplier_16x16bit_pipelined.layer_1_full_adder_4.A ;
  assign \multiplier_16x16bit_pipelined.layer_0_w14[6] = \multiplier_16x16bit_pipelined.layer_1_full_adder_4.B ;
  assign \multiplier_16x16bit_pipelined.layer_0_w14[7] = \multiplier_16x16bit_pipelined.layer_1_full_adder_4.cin ;
  assign \multiplier_16x16bit_pipelined.layer_0_w14[8] = \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_7.negation ;
  assign \multiplier_16x16bit_pipelined.layer_0_w15[0] = \multiplier_16x16bit_pipelined.layer_1_compressor42_8.A ;
  assign \multiplier_16x16bit_pipelined.layer_0_w15[1] = \multiplier_16x16bit_pipelined.layer_1_compressor42_8.B ;
  assign \multiplier_16x16bit_pipelined.layer_0_w15[2] = \multiplier_16x16bit_pipelined.layer_1_compressor42_8.C ;
  assign \multiplier_16x16bit_pipelined.layer_0_w15[3] = \multiplier_16x16bit_pipelined.layer_1_compressor42_8.D ;
  assign \multiplier_16x16bit_pipelined.layer_0_w15[4] = \multiplier_16x16bit_pipelined.layer_1_compressor42_8.cin ;
  assign \multiplier_16x16bit_pipelined.layer_0_w15[5] = \multiplier_16x16bit_pipelined.layer_1_full_adder_5.A ;
  assign \multiplier_16x16bit_pipelined.layer_0_w15[6] = \multiplier_16x16bit_pipelined.layer_1_full_adder_5.B ;
  assign \multiplier_16x16bit_pipelined.layer_0_w15[7] = \multiplier_16x16bit_pipelined.layer_1_full_adder_5.cin ;
  assign \multiplier_16x16bit_pipelined.layer_0_w16[0] = \multiplier_16x16bit_pipelined.layer_1_compressor42_9.A ;
  assign \multiplier_16x16bit_pipelined.layer_0_w16[1] = \multiplier_16x16bit_pipelined.layer_1_compressor42_9.B ;
  assign \multiplier_16x16bit_pipelined.layer_0_w16[2] = \multiplier_16x16bit_pipelined.layer_1_compressor42_9.C ;
  assign \multiplier_16x16bit_pipelined.layer_0_w16[3] = \multiplier_16x16bit_pipelined.layer_1_compressor42_9.D ;
  assign \multiplier_16x16bit_pipelined.layer_0_w16[4] = \multiplier_16x16bit_pipelined.layer_1_compressor42_9.cin ;
  assign \multiplier_16x16bit_pipelined.layer_0_w16[5] = \multiplier_16x16bit_pipelined.layer_1_full_adder_6.A ;
  assign \multiplier_16x16bit_pipelined.layer_0_w16[6] = \multiplier_16x16bit_pipelined.layer_1_full_adder_6.B ;
  assign \multiplier_16x16bit_pipelined.layer_0_w16[7] = \multiplier_16x16bit_pipelined.layer_1_full_adder_6.cin ;
  assign \multiplier_16x16bit_pipelined.layer_0_w17[0] = \multiplier_16x16bit_pipelined.layer_1_compressor42_10.A ;
  assign \multiplier_16x16bit_pipelined.layer_0_w17[1] = \multiplier_16x16bit_pipelined.layer_1_compressor42_10.B ;
  assign \multiplier_16x16bit_pipelined.layer_0_w17[2] = \multiplier_16x16bit_pipelined.layer_1_compressor42_10.C ;
  assign \multiplier_16x16bit_pipelined.layer_0_w17[3] = \multiplier_16x16bit_pipelined.layer_1_compressor42_10.D ;
  assign \multiplier_16x16bit_pipelined.layer_0_w17[4] = \multiplier_16x16bit_pipelined.layer_1_compressor42_10.cin ;
  assign \multiplier_16x16bit_pipelined.layer_0_w17[5] = \multiplier_16x16bit_pipelined.layer_1_full_adder_7.A ;
  assign \multiplier_16x16bit_pipelined.layer_0_w17[6] = \multiplier_16x16bit_pipelined.layer_1_full_adder_7.B ;
  assign \multiplier_16x16bit_pipelined.layer_0_w18[0] = \multiplier_16x16bit_pipelined.layer_1_compressor42_11.A ;
  assign \multiplier_16x16bit_pipelined.layer_0_w18[1] = \multiplier_16x16bit_pipelined.layer_1_compressor42_11.B ;
  assign \multiplier_16x16bit_pipelined.layer_0_w18[2] = \multiplier_16x16bit_pipelined.layer_1_compressor42_11.C ;
  assign \multiplier_16x16bit_pipelined.layer_0_w18[3] = \multiplier_16x16bit_pipelined.layer_1_compressor42_11.D ;
  assign \multiplier_16x16bit_pipelined.layer_0_w18[4] = \multiplier_16x16bit_pipelined.layer_1_compressor42_11.cin ;
  assign \multiplier_16x16bit_pipelined.layer_0_w18[5] = \multiplier_16x16bit_pipelined.layer_2_compressor42_6.cin ;
  assign \multiplier_16x16bit_pipelined.layer_0_w19[0] = \multiplier_16x16bit_pipelined.layer_1_compressor42_12.A ;
  assign \multiplier_16x16bit_pipelined.layer_0_w19[1] = \multiplier_16x16bit_pipelined.layer_1_compressor42_12.B ;
  assign \multiplier_16x16bit_pipelined.layer_0_w19[2] = \multiplier_16x16bit_pipelined.layer_1_compressor42_12.C ;
  assign \multiplier_16x16bit_pipelined.layer_0_w19[3] = \multiplier_16x16bit_pipelined.layer_1_compressor42_12.D ;
  assign \multiplier_16x16bit_pipelined.layer_0_w19[4] = \multiplier_16x16bit_pipelined.layer_1_compressor42_12.cin ;
  assign \multiplier_16x16bit_pipelined.layer_0_w19[5] = \multiplier_16x16bit_pipelined.layer_2_compressor42_7.D ;
  assign \multiplier_16x16bit_pipelined.layer_0_w20[0] = \multiplier_16x16bit_pipelined.layer_1_compressor42_13.A ;
  assign \multiplier_16x16bit_pipelined.layer_0_w20[1] = \multiplier_16x16bit_pipelined.layer_1_compressor42_13.B ;
  assign \multiplier_16x16bit_pipelined.layer_0_w20[2] = \multiplier_16x16bit_pipelined.layer_1_compressor42_13.C ;
  assign \multiplier_16x16bit_pipelined.layer_0_w20[3] = \multiplier_16x16bit_pipelined.layer_1_compressor42_13.D ;
  assign \multiplier_16x16bit_pipelined.layer_0_w20[4] = \multiplier_16x16bit_pipelined.layer_1_compressor42_13.cin ;
  assign \multiplier_16x16bit_pipelined.layer_0_w21[0] = \multiplier_16x16bit_pipelined.layer_1_compressor42_14.A ;
  assign \multiplier_16x16bit_pipelined.layer_0_w21[1] = \multiplier_16x16bit_pipelined.layer_1_compressor42_14.B ;
  assign \multiplier_16x16bit_pipelined.layer_0_w21[2] = \multiplier_16x16bit_pipelined.layer_1_compressor42_14.C ;
  assign \multiplier_16x16bit_pipelined.layer_0_w21[3] = \multiplier_16x16bit_pipelined.layer_1_compressor42_14.D ;
  assign \multiplier_16x16bit_pipelined.layer_0_w21[4] = \multiplier_16x16bit_pipelined.layer_1_compressor42_14.cin ;
  assign \multiplier_16x16bit_pipelined.layer_0_w22[0] = \multiplier_16x16bit_pipelined.layer_1_compressor42_15.A ;
  assign \multiplier_16x16bit_pipelined.layer_0_w22[1] = \multiplier_16x16bit_pipelined.layer_1_compressor42_15.B ;
  assign \multiplier_16x16bit_pipelined.layer_0_w22[2] = \multiplier_16x16bit_pipelined.layer_1_compressor42_15.C ;
  assign \multiplier_16x16bit_pipelined.layer_0_w22[3] = \multiplier_16x16bit_pipelined.layer_1_compressor42_15.D ;
  assign \multiplier_16x16bit_pipelined.layer_0_w22[4] = \multiplier_16x16bit_pipelined.layer_1_compressor42_15.cin ;
  assign \multiplier_16x16bit_pipelined.layer_0_w23[0] = \multiplier_16x16bit_pipelined.layer_1_compressor42_16.A ;
  assign \multiplier_16x16bit_pipelined.layer_0_w23[1] = \multiplier_16x16bit_pipelined.layer_1_compressor42_16.B ;
  assign \multiplier_16x16bit_pipelined.layer_0_w23[2] = \multiplier_16x16bit_pipelined.layer_1_compressor42_16.C ;
  assign \multiplier_16x16bit_pipelined.layer_0_w23[3] = \multiplier_16x16bit_pipelined.layer_1_compressor42_16.D ;
  assign \multiplier_16x16bit_pipelined.layer_0_w24[0] = \multiplier_16x16bit_pipelined.layer_1_full_adder_8.A ;
  assign \multiplier_16x16bit_pipelined.layer_0_w24[1] = \multiplier_16x16bit_pipelined.layer_1_full_adder_8.B ;
  assign \multiplier_16x16bit_pipelined.layer_0_w24[2] = \multiplier_16x16bit_pipelined.layer_1_full_adder_8.cin ;
  assign \multiplier_16x16bit_pipelined.layer_0_w25[0] = \multiplier_16x16bit_pipelined.layer_1_full_adder_9.A ;
  assign \multiplier_16x16bit_pipelined.layer_0_w25[1] = \multiplier_16x16bit_pipelined.layer_1_full_adder_9.B ;
  assign \multiplier_16x16bit_pipelined.layer_0_w25[2] = \multiplier_16x16bit_pipelined.layer_1_full_adder_9.cin ;
  assign \multiplier_16x16bit_pipelined.layer_0_w26[0] = \multiplier_16x16bit_pipelined.layer_1_full_adder_10.A ;
  assign \multiplier_16x16bit_pipelined.layer_0_w26[1] = \multiplier_16x16bit_pipelined.layer_1_full_adder_10.B ;
  assign \multiplier_16x16bit_pipelined.layer_0_w26[2] = \multiplier_16x16bit_pipelined.layer_1_full_adder_10.cin ;
  assign \multiplier_16x16bit_pipelined.layer_0_w27[0] = \multiplier_16x16bit_pipelined.layer_1_full_adder_11.A ;
  assign \multiplier_16x16bit_pipelined.layer_0_w27[1] = \multiplier_16x16bit_pipelined.layer_1_full_adder_11.B ;
  assign \multiplier_16x16bit_pipelined.layer_0_w28[0] = \multiplier_16x16bit_pipelined.layer_2_full_adder_11.B ;
  assign \multiplier_16x16bit_pipelined.layer_0_w28[1] = \multiplier_16x16bit_pipelined.layer_2_full_adder_11.cin ;
  assign \multiplier_16x16bit_pipelined.layer_0_w2[2] = \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_1.negation ;
  assign \multiplier_16x16bit_pipelined.layer_0_w4[0] = \multiplier_16x16bit_pipelined.layer_1_full_adder_0.A ;
  assign \multiplier_16x16bit_pipelined.layer_0_w4[1] = \multiplier_16x16bit_pipelined.layer_1_full_adder_0.B ;
  assign \multiplier_16x16bit_pipelined.layer_0_w4[2] = \multiplier_16x16bit_pipelined.layer_1_full_adder_0.cin ;
  assign \multiplier_16x16bit_pipelined.layer_0_w4[3] = \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_2.negation ;
  assign \multiplier_16x16bit_pipelined.layer_0_w5[0] = \multiplier_16x16bit_pipelined.layer_1_full_adder_1.A ;
  assign \multiplier_16x16bit_pipelined.layer_0_w5[1] = \multiplier_16x16bit_pipelined.layer_1_full_adder_1.B ;
  assign \multiplier_16x16bit_pipelined.layer_0_w5[2] = \multiplier_16x16bit_pipelined.layer_1_full_adder_1.cin ;
  assign \multiplier_16x16bit_pipelined.layer_0_w6[0] = \multiplier_16x16bit_pipelined.layer_1_compressor42_0.A ;
  assign \multiplier_16x16bit_pipelined.layer_0_w6[1] = \multiplier_16x16bit_pipelined.layer_1_compressor42_0.B ;
  assign \multiplier_16x16bit_pipelined.layer_0_w6[2] = \multiplier_16x16bit_pipelined.layer_1_compressor42_0.C ;
  assign \multiplier_16x16bit_pipelined.layer_0_w6[3] = \multiplier_16x16bit_pipelined.layer_1_compressor42_0.D ;
  assign \multiplier_16x16bit_pipelined.layer_0_w6[4] = \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_3.negation ;
  assign \multiplier_16x16bit_pipelined.layer_0_w7[0] = \multiplier_16x16bit_pipelined.layer_1_full_adder_2.A ;
  assign \multiplier_16x16bit_pipelined.layer_0_w7[1] = \multiplier_16x16bit_pipelined.layer_1_full_adder_2.B ;
  assign \multiplier_16x16bit_pipelined.layer_0_w7[2] = \multiplier_16x16bit_pipelined.layer_1_full_adder_2.cin ;
  assign \multiplier_16x16bit_pipelined.layer_0_w8[0] = \multiplier_16x16bit_pipelined.layer_1_compressor42_1.A ;
  assign \multiplier_16x16bit_pipelined.layer_0_w8[1] = \multiplier_16x16bit_pipelined.layer_1_compressor42_1.B ;
  assign \multiplier_16x16bit_pipelined.layer_0_w8[2] = \multiplier_16x16bit_pipelined.layer_1_compressor42_1.C ;
  assign \multiplier_16x16bit_pipelined.layer_0_w8[3] = \multiplier_16x16bit_pipelined.layer_1_compressor42_1.D ;
  assign \multiplier_16x16bit_pipelined.layer_0_w8[4] = \multiplier_16x16bit_pipelined.layer_1_compressor42_1.cin ;
  assign \multiplier_16x16bit_pipelined.layer_0_w8[5] = \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_4.negation ;
  assign \multiplier_16x16bit_pipelined.layer_0_w9[0] = \multiplier_16x16bit_pipelined.layer_1_compressor42_2.A ;
  assign \multiplier_16x16bit_pipelined.layer_0_w9[1] = \multiplier_16x16bit_pipelined.layer_1_compressor42_2.B ;
  assign \multiplier_16x16bit_pipelined.layer_0_w9[2] = \multiplier_16x16bit_pipelined.layer_1_compressor42_2.C ;
  assign \multiplier_16x16bit_pipelined.layer_0_w9[3] = \multiplier_16x16bit_pipelined.layer_1_compressor42_2.D ;
  assign \multiplier_16x16bit_pipelined.layer_0_w9[4] = \multiplier_16x16bit_pipelined.layer_1_compressor42_2.cin ;
  assign \multiplier_16x16bit_pipelined.layer_1_compressor42_0.cin = \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_3.negation ;
  assign \multiplier_16x16bit_pipelined.layer_1_full_adder_3.cin = \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_6.negation ;
  assign \multiplier_16x16bit_pipelined.layer_1_w0[0] = \multiplier_16x16bit_pipelined.layer_0_w0[0] ;
  assign \multiplier_16x16bit_pipelined.layer_1_w0[1] = \multiplier_16x16bit_pipelined.mr [1];
  assign \multiplier_16x16bit_pipelined.layer_1_w1 = \multiplier_16x16bit_pipelined.layer_0_w1 ;
  assign \multiplier_16x16bit_pipelined.layer_1_w10[0] = \multiplier_16x16bit_pipelined.layer_1_compressor42_2.carry ;
  assign \multiplier_16x16bit_pipelined.layer_1_w10[1] = \multiplier_16x16bit_pipelined.layer_1_compressor42_2.cout ;
  assign \multiplier_16x16bit_pipelined.layer_1_w10[2] = \multiplier_16x16bit_pipelined.layer_1_compressor42_3.S ;
  assign \multiplier_16x16bit_pipelined.layer_1_w10[3] = \multiplier_16x16bit_pipelined.layer_2_compressor42_0.D ;
  assign \multiplier_16x16bit_pipelined.layer_1_w10[4] = \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_5.negation ;
  assign \multiplier_16x16bit_pipelined.layer_1_w11[0] = \multiplier_16x16bit_pipelined.layer_1_compressor42_3.carry ;
  assign \multiplier_16x16bit_pipelined.layer_1_w11[1] = \multiplier_16x16bit_pipelined.layer_1_compressor42_3.cout ;
  assign \multiplier_16x16bit_pipelined.layer_1_w11[2] = \multiplier_16x16bit_pipelined.layer_1_compressor42_4.S ;
  assign \multiplier_16x16bit_pipelined.layer_1_w11[3] = \multiplier_16x16bit_pipelined.layer_0_w11[5] ;
  assign \multiplier_16x16bit_pipelined.layer_1_w12[0] = \multiplier_16x16bit_pipelined.layer_1_compressor42_4.carry ;
  assign \multiplier_16x16bit_pipelined.layer_1_w12[1] = \multiplier_16x16bit_pipelined.layer_1_compressor42_4.cout ;
  assign \multiplier_16x16bit_pipelined.layer_1_w12[2] = \multiplier_16x16bit_pipelined.layer_1_compressor42_5.S ;
  assign \multiplier_16x16bit_pipelined.layer_1_w12[3] = \multiplier_16x16bit_pipelined.layer_1_full_adder_3.S ;
  assign \multiplier_16x16bit_pipelined.layer_1_w13[0] = \multiplier_16x16bit_pipelined.layer_1_compressor42_5.carry ;
  assign \multiplier_16x16bit_pipelined.layer_1_w13[1] = \multiplier_16x16bit_pipelined.layer_1_compressor42_5.cout ;
  assign \multiplier_16x16bit_pipelined.layer_1_w13[2] = \multiplier_16x16bit_pipelined.layer_1_full_adder_3.cout ;
  assign \multiplier_16x16bit_pipelined.layer_1_w13[3] = \multiplier_16x16bit_pipelined.layer_1_compressor42_6.S ;
  assign \multiplier_16x16bit_pipelined.layer_1_w13[4] = \multiplier_16x16bit_pipelined.layer_2_compressor42_1.cin ;
  assign \multiplier_16x16bit_pipelined.layer_1_w13[5] = \multiplier_16x16bit_pipelined.layer_0_w13[6] ;
  assign \multiplier_16x16bit_pipelined.layer_1_w14[0] = \multiplier_16x16bit_pipelined.layer_1_compressor42_6.carry ;
  assign \multiplier_16x16bit_pipelined.layer_1_w14[1] = \multiplier_16x16bit_pipelined.layer_1_compressor42_6.cout ;
  assign \multiplier_16x16bit_pipelined.layer_1_w14[2] = \multiplier_16x16bit_pipelined.layer_1_compressor42_7.S ;
  assign \multiplier_16x16bit_pipelined.layer_1_w14[3] = \multiplier_16x16bit_pipelined.layer_1_full_adder_4.S ;
  assign \multiplier_16x16bit_pipelined.layer_1_w14[4] = \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_7.negation ;
  assign \multiplier_16x16bit_pipelined.layer_1_w15[0] = \multiplier_16x16bit_pipelined.layer_1_compressor42_7.carry ;
  assign \multiplier_16x16bit_pipelined.layer_1_w15[1] = \multiplier_16x16bit_pipelined.layer_1_compressor42_7.cout ;
  assign \multiplier_16x16bit_pipelined.layer_1_w15[2] = \multiplier_16x16bit_pipelined.layer_1_full_adder_4.cout ;
  assign \multiplier_16x16bit_pipelined.layer_1_w15[3] = \multiplier_16x16bit_pipelined.layer_1_compressor42_8.S ;
  assign \multiplier_16x16bit_pipelined.layer_1_w15[4] = \multiplier_16x16bit_pipelined.layer_1_full_adder_5.S ;
  assign \multiplier_16x16bit_pipelined.layer_1_w16[0] = \multiplier_16x16bit_pipelined.layer_1_compressor42_8.carry ;
  assign \multiplier_16x16bit_pipelined.layer_1_w16[1] = \multiplier_16x16bit_pipelined.layer_1_compressor42_8.cout ;
  assign \multiplier_16x16bit_pipelined.layer_1_w16[2] = \multiplier_16x16bit_pipelined.layer_1_full_adder_5.cout ;
  assign \multiplier_16x16bit_pipelined.layer_1_w16[3] = \multiplier_16x16bit_pipelined.layer_1_compressor42_9.S ;
  assign \multiplier_16x16bit_pipelined.layer_1_w16[4] = \multiplier_16x16bit_pipelined.layer_1_full_adder_6.S ;
  assign \multiplier_16x16bit_pipelined.layer_1_w17[0] = \multiplier_16x16bit_pipelined.layer_1_compressor42_9.carry ;
  assign \multiplier_16x16bit_pipelined.layer_1_w17[1] = \multiplier_16x16bit_pipelined.layer_1_compressor42_9.cout ;
  assign \multiplier_16x16bit_pipelined.layer_1_w17[2] = \multiplier_16x16bit_pipelined.layer_1_full_adder_6.cout ;
  assign \multiplier_16x16bit_pipelined.layer_1_w17[3] = \multiplier_16x16bit_pipelined.layer_1_compressor42_10.S ;
  assign \multiplier_16x16bit_pipelined.layer_1_w17[4] = \multiplier_16x16bit_pipelined.layer_1_full_adder_7.S ;
  assign \multiplier_16x16bit_pipelined.layer_1_w18[0] = \multiplier_16x16bit_pipelined.layer_1_compressor42_10.carry ;
  assign \multiplier_16x16bit_pipelined.layer_1_w18[1] = \multiplier_16x16bit_pipelined.layer_1_compressor42_10.cout ;
  assign \multiplier_16x16bit_pipelined.layer_1_w18[2] = \multiplier_16x16bit_pipelined.layer_1_full_adder_7.cout ;
  assign \multiplier_16x16bit_pipelined.layer_1_w18[3] = \multiplier_16x16bit_pipelined.layer_1_compressor42_11.S ;
  assign \multiplier_16x16bit_pipelined.layer_1_w18[4] = \multiplier_16x16bit_pipelined.layer_2_compressor42_6.cin ;
  assign \multiplier_16x16bit_pipelined.layer_1_w18[5] = \multiplier_16x16bit_pipelined.layer_0_w18[6] ;
  assign \multiplier_16x16bit_pipelined.layer_1_w19[0] = \multiplier_16x16bit_pipelined.layer_1_compressor42_11.carry ;
  assign \multiplier_16x16bit_pipelined.layer_1_w19[1] = \multiplier_16x16bit_pipelined.layer_1_compressor42_11.cout ;
  assign \multiplier_16x16bit_pipelined.layer_1_w19[2] = \multiplier_16x16bit_pipelined.layer_1_compressor42_12.S ;
  assign \multiplier_16x16bit_pipelined.layer_1_w19[3] = \multiplier_16x16bit_pipelined.layer_2_compressor42_7.D ;
  assign \multiplier_16x16bit_pipelined.layer_1_w20[0] = \multiplier_16x16bit_pipelined.layer_1_compressor42_12.carry ;
  assign \multiplier_16x16bit_pipelined.layer_1_w20[1] = \multiplier_16x16bit_pipelined.layer_1_compressor42_12.cout ;
  assign \multiplier_16x16bit_pipelined.layer_1_w20[2] = \multiplier_16x16bit_pipelined.layer_1_compressor42_13.S ;
  assign \multiplier_16x16bit_pipelined.layer_1_w20[3] = \multiplier_16x16bit_pipelined.layer_0_w20[5] ;
  assign \multiplier_16x16bit_pipelined.layer_1_w21[0] = \multiplier_16x16bit_pipelined.layer_1_compressor42_13.carry ;
  assign \multiplier_16x16bit_pipelined.layer_1_w21[1] = \multiplier_16x16bit_pipelined.layer_1_compressor42_13.cout ;
  assign \multiplier_16x16bit_pipelined.layer_1_w21[2] = \multiplier_16x16bit_pipelined.layer_1_compressor42_14.S ;
  assign \multiplier_16x16bit_pipelined.layer_1_w22[0] = \multiplier_16x16bit_pipelined.layer_1_compressor42_14.carry ;
  assign \multiplier_16x16bit_pipelined.layer_1_w22[1] = \multiplier_16x16bit_pipelined.layer_1_compressor42_14.cout ;
  assign \multiplier_16x16bit_pipelined.layer_1_w22[2] = \multiplier_16x16bit_pipelined.layer_1_compressor42_15.S ;
  assign \multiplier_16x16bit_pipelined.layer_1_w23[0] = \multiplier_16x16bit_pipelined.layer_1_compressor42_15.carry ;
  assign \multiplier_16x16bit_pipelined.layer_1_w23[1] = \multiplier_16x16bit_pipelined.layer_1_compressor42_15.cout ;
  assign \multiplier_16x16bit_pipelined.layer_1_w23[2] = \multiplier_16x16bit_pipelined.layer_1_compressor42_16.S ;
  assign \multiplier_16x16bit_pipelined.layer_1_w24[0] = \multiplier_16x16bit_pipelined.layer_1_compressor42_16.carry ;
  assign \multiplier_16x16bit_pipelined.layer_1_w24[1] = \multiplier_16x16bit_pipelined.layer_1_compressor42_16.cout ;
  assign \multiplier_16x16bit_pipelined.layer_1_w24[2] = \multiplier_16x16bit_pipelined.layer_1_full_adder_8.S ;
  assign \multiplier_16x16bit_pipelined.layer_1_w24[3] = \multiplier_16x16bit_pipelined.layer_0_w24[3] ;
  assign \multiplier_16x16bit_pipelined.layer_1_w25[0] = \multiplier_16x16bit_pipelined.layer_1_full_adder_8.cout ;
  assign \multiplier_16x16bit_pipelined.layer_1_w25[1] = \multiplier_16x16bit_pipelined.layer_1_full_adder_9.S ;
  assign \multiplier_16x16bit_pipelined.layer_1_w26[0] = \multiplier_16x16bit_pipelined.layer_1_full_adder_9.cout ;
  assign \multiplier_16x16bit_pipelined.layer_1_w26[1] = \multiplier_16x16bit_pipelined.layer_1_full_adder_10.S ;
  assign \multiplier_16x16bit_pipelined.layer_1_w27[0] = \multiplier_16x16bit_pipelined.layer_1_full_adder_10.cout ;
  assign \multiplier_16x16bit_pipelined.layer_1_w27[1] = \multiplier_16x16bit_pipelined.layer_1_full_adder_11.S ;
  assign \multiplier_16x16bit_pipelined.layer_1_w28[0] = \multiplier_16x16bit_pipelined.layer_1_full_adder_11.cout ;
  assign \multiplier_16x16bit_pipelined.layer_1_w28[1] = \multiplier_16x16bit_pipelined.layer_2_full_adder_11.B ;
  assign \multiplier_16x16bit_pipelined.layer_1_w28[2] = \multiplier_16x16bit_pipelined.layer_2_full_adder_11.cin ;
  assign \multiplier_16x16bit_pipelined.layer_1_w29[0] = \multiplier_16x16bit_pipelined.layer_0_w29[0] ;
  assign \multiplier_16x16bit_pipelined.layer_1_w2[0] = \multiplier_16x16bit_pipelined.layer_0_w2[0] ;
  assign \multiplier_16x16bit_pipelined.layer_1_w2[1] = \multiplier_16x16bit_pipelined.layer_0_w2[1] ;
  assign \multiplier_16x16bit_pipelined.layer_1_w2[2] = \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_1.negation ;
  assign \multiplier_16x16bit_pipelined.layer_1_w30 = \multiplier_16x16bit_pipelined.layer_0_w30 ;
  assign \multiplier_16x16bit_pipelined.layer_1_w3[0] = \multiplier_16x16bit_pipelined.layer_0_w3[0] ;
  assign \multiplier_16x16bit_pipelined.layer_1_w3[1] = \multiplier_16x16bit_pipelined.layer_0_w3[1] ;
  assign \multiplier_16x16bit_pipelined.layer_1_w4[0] = \multiplier_16x16bit_pipelined.layer_1_full_adder_0.S ;
  assign \multiplier_16x16bit_pipelined.layer_1_w4[1] = \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_2.negation ;
  assign \multiplier_16x16bit_pipelined.layer_1_w5[0] = \multiplier_16x16bit_pipelined.layer_1_full_adder_0.cout ;
  assign \multiplier_16x16bit_pipelined.layer_1_w5[1] = \multiplier_16x16bit_pipelined.layer_1_full_adder_1.S ;
  assign \multiplier_16x16bit_pipelined.layer_1_w6[0] = \multiplier_16x16bit_pipelined.layer_1_full_adder_1.cout ;
  assign \multiplier_16x16bit_pipelined.layer_1_w6[1] = \multiplier_16x16bit_pipelined.layer_1_compressor42_0.S ;
  assign \multiplier_16x16bit_pipelined.layer_1_w7[0] = \multiplier_16x16bit_pipelined.layer_1_compressor42_0.carry ;
  assign \multiplier_16x16bit_pipelined.layer_1_w7[1] = \multiplier_16x16bit_pipelined.layer_1_compressor42_0.cout ;
  assign \multiplier_16x16bit_pipelined.layer_1_w7[2] = \multiplier_16x16bit_pipelined.layer_1_full_adder_2.S ;
  assign \multiplier_16x16bit_pipelined.layer_1_w7[3] = \multiplier_16x16bit_pipelined.layer_0_w7[3] ;
  assign \multiplier_16x16bit_pipelined.layer_1_w8[0] = \multiplier_16x16bit_pipelined.layer_1_full_adder_2.cout ;
  assign \multiplier_16x16bit_pipelined.layer_1_w8[1] = \multiplier_16x16bit_pipelined.layer_1_compressor42_1.S ;
  assign \multiplier_16x16bit_pipelined.layer_1_w8[2] = \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_4.negation ;
  assign \multiplier_16x16bit_pipelined.layer_1_w9[0] = \multiplier_16x16bit_pipelined.layer_1_compressor42_1.carry ;
  assign \multiplier_16x16bit_pipelined.layer_1_w9[1] = \multiplier_16x16bit_pipelined.layer_1_compressor42_1.cout ;
  assign \multiplier_16x16bit_pipelined.layer_1_w9[2] = \multiplier_16x16bit_pipelined.layer_1_compressor42_2.S ;
  assign \multiplier_16x16bit_pipelined.layer_2_compressor42_0.A = \multiplier_16x16bit_pipelined.layer_1_compressor42_2.carry ;
  assign \multiplier_16x16bit_pipelined.layer_2_compressor42_0.B = \multiplier_16x16bit_pipelined.layer_1_compressor42_2.cout ;
  assign \multiplier_16x16bit_pipelined.layer_2_compressor42_0.C = \multiplier_16x16bit_pipelined.layer_1_compressor42_3.S ;
  assign \multiplier_16x16bit_pipelined.layer_2_compressor42_0.cin = \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_5.negation ;
  assign \multiplier_16x16bit_pipelined.layer_2_compressor42_1.A = \multiplier_16x16bit_pipelined.layer_1_compressor42_5.carry ;
  assign \multiplier_16x16bit_pipelined.layer_2_compressor42_1.B = \multiplier_16x16bit_pipelined.layer_1_compressor42_5.cout ;
  assign \multiplier_16x16bit_pipelined.layer_2_compressor42_1.C = \multiplier_16x16bit_pipelined.layer_1_full_adder_3.cout ;
  assign \multiplier_16x16bit_pipelined.layer_2_compressor42_1.D = \multiplier_16x16bit_pipelined.layer_1_compressor42_6.S ;
  assign \multiplier_16x16bit_pipelined.layer_2_compressor42_2.A = \multiplier_16x16bit_pipelined.layer_1_compressor42_6.carry ;
  assign \multiplier_16x16bit_pipelined.layer_2_compressor42_2.B = \multiplier_16x16bit_pipelined.layer_1_compressor42_6.cout ;
  assign \multiplier_16x16bit_pipelined.layer_2_compressor42_2.C = \multiplier_16x16bit_pipelined.layer_1_compressor42_7.S ;
  assign \multiplier_16x16bit_pipelined.layer_2_compressor42_2.D = \multiplier_16x16bit_pipelined.layer_1_full_adder_4.S ;
  assign \multiplier_16x16bit_pipelined.layer_2_compressor42_2.cin = \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_7.negation ;
  assign \multiplier_16x16bit_pipelined.layer_2_compressor42_3.A = \multiplier_16x16bit_pipelined.layer_1_compressor42_7.carry ;
  assign \multiplier_16x16bit_pipelined.layer_2_compressor42_3.B = \multiplier_16x16bit_pipelined.layer_1_compressor42_7.cout ;
  assign \multiplier_16x16bit_pipelined.layer_2_compressor42_3.C = \multiplier_16x16bit_pipelined.layer_1_full_adder_4.cout ;
  assign \multiplier_16x16bit_pipelined.layer_2_compressor42_3.D = \multiplier_16x16bit_pipelined.layer_1_compressor42_8.S ;
  assign \multiplier_16x16bit_pipelined.layer_2_compressor42_3.cin = \multiplier_16x16bit_pipelined.layer_1_full_adder_5.S ;
  assign \multiplier_16x16bit_pipelined.layer_2_compressor42_4.A = \multiplier_16x16bit_pipelined.layer_1_compressor42_8.carry ;
  assign \multiplier_16x16bit_pipelined.layer_2_compressor42_4.B = \multiplier_16x16bit_pipelined.layer_1_compressor42_8.cout ;
  assign \multiplier_16x16bit_pipelined.layer_2_compressor42_4.C = \multiplier_16x16bit_pipelined.layer_1_full_adder_5.cout ;
  assign \multiplier_16x16bit_pipelined.layer_2_compressor42_4.D = \multiplier_16x16bit_pipelined.layer_1_compressor42_9.S ;
  assign \multiplier_16x16bit_pipelined.layer_2_compressor42_4.cin = \multiplier_16x16bit_pipelined.layer_1_full_adder_6.S ;
  assign \multiplier_16x16bit_pipelined.layer_2_compressor42_5.A = \multiplier_16x16bit_pipelined.layer_1_compressor42_9.carry ;
  assign \multiplier_16x16bit_pipelined.layer_2_compressor42_5.B = \multiplier_16x16bit_pipelined.layer_1_compressor42_9.cout ;
  assign \multiplier_16x16bit_pipelined.layer_2_compressor42_5.C = \multiplier_16x16bit_pipelined.layer_1_full_adder_6.cout ;
  assign \multiplier_16x16bit_pipelined.layer_2_compressor42_5.D = \multiplier_16x16bit_pipelined.layer_1_compressor42_10.S ;
  assign \multiplier_16x16bit_pipelined.layer_2_compressor42_5.cin = \multiplier_16x16bit_pipelined.layer_1_full_adder_7.S ;
  assign \multiplier_16x16bit_pipelined.layer_2_compressor42_6.A = \multiplier_16x16bit_pipelined.layer_1_compressor42_10.carry ;
  assign \multiplier_16x16bit_pipelined.layer_2_compressor42_6.B = \multiplier_16x16bit_pipelined.layer_1_compressor42_10.cout ;
  assign \multiplier_16x16bit_pipelined.layer_2_compressor42_6.C = \multiplier_16x16bit_pipelined.layer_1_full_adder_7.cout ;
  assign \multiplier_16x16bit_pipelined.layer_2_compressor42_6.D = \multiplier_16x16bit_pipelined.layer_1_compressor42_11.S ;
  assign \multiplier_16x16bit_pipelined.layer_2_compressor42_7.A = \multiplier_16x16bit_pipelined.layer_1_compressor42_11.carry ;
  assign \multiplier_16x16bit_pipelined.layer_2_compressor42_7.B = \multiplier_16x16bit_pipelined.layer_1_compressor42_11.cout ;
  assign \multiplier_16x16bit_pipelined.layer_2_compressor42_7.C = \multiplier_16x16bit_pipelined.layer_1_compressor42_12.S ;
  assign \multiplier_16x16bit_pipelined.layer_2_full_adder_0.A = \multiplier_16x16bit_pipelined.layer_1_compressor42_0.carry ;
  assign \multiplier_16x16bit_pipelined.layer_2_full_adder_0.B = \multiplier_16x16bit_pipelined.layer_1_compressor42_0.cout ;
  assign \multiplier_16x16bit_pipelined.layer_2_full_adder_0.cin = \multiplier_16x16bit_pipelined.layer_1_full_adder_2.S ;
  assign \multiplier_16x16bit_pipelined.layer_2_full_adder_1.A = \multiplier_16x16bit_pipelined.layer_1_full_adder_2.cout ;
  assign \multiplier_16x16bit_pipelined.layer_2_full_adder_1.B = \multiplier_16x16bit_pipelined.layer_1_compressor42_1.S ;
  assign \multiplier_16x16bit_pipelined.layer_2_full_adder_1.cin = \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_4.negation ;
  assign \multiplier_16x16bit_pipelined.layer_2_full_adder_10.A = \multiplier_16x16bit_pipelined.layer_1_full_adder_8.cout ;
  assign \multiplier_16x16bit_pipelined.layer_2_full_adder_10.B = \multiplier_16x16bit_pipelined.layer_1_full_adder_9.S ;
  assign \multiplier_16x16bit_pipelined.layer_2_full_adder_11.A = \multiplier_16x16bit_pipelined.layer_1_full_adder_11.cout ;
  assign \multiplier_16x16bit_pipelined.layer_2_full_adder_2.A = \multiplier_16x16bit_pipelined.layer_1_compressor42_1.carry ;
  assign \multiplier_16x16bit_pipelined.layer_2_full_adder_2.B = \multiplier_16x16bit_pipelined.layer_1_compressor42_1.cout ;
  assign \multiplier_16x16bit_pipelined.layer_2_full_adder_2.cin = \multiplier_16x16bit_pipelined.layer_1_compressor42_2.S ;
  assign \multiplier_16x16bit_pipelined.layer_2_full_adder_3.A = \multiplier_16x16bit_pipelined.layer_1_compressor42_3.carry ;
  assign \multiplier_16x16bit_pipelined.layer_2_full_adder_3.B = \multiplier_16x16bit_pipelined.layer_1_compressor42_3.cout ;
  assign \multiplier_16x16bit_pipelined.layer_2_full_adder_3.cin = \multiplier_16x16bit_pipelined.layer_1_compressor42_4.S ;
  assign \multiplier_16x16bit_pipelined.layer_2_full_adder_4.A = \multiplier_16x16bit_pipelined.layer_1_compressor42_4.carry ;
  assign \multiplier_16x16bit_pipelined.layer_2_full_adder_4.B = \multiplier_16x16bit_pipelined.layer_1_compressor42_4.cout ;
  assign \multiplier_16x16bit_pipelined.layer_2_full_adder_4.cin = \multiplier_16x16bit_pipelined.layer_1_compressor42_5.S ;
  assign \multiplier_16x16bit_pipelined.layer_2_full_adder_5.A = \multiplier_16x16bit_pipelined.layer_1_compressor42_12.carry ;
  assign \multiplier_16x16bit_pipelined.layer_2_full_adder_5.B = \multiplier_16x16bit_pipelined.layer_1_compressor42_12.cout ;
  assign \multiplier_16x16bit_pipelined.layer_2_full_adder_5.cin = \multiplier_16x16bit_pipelined.layer_1_compressor42_13.S ;
  assign \multiplier_16x16bit_pipelined.layer_2_full_adder_6.A = \multiplier_16x16bit_pipelined.layer_1_compressor42_13.carry ;
  assign \multiplier_16x16bit_pipelined.layer_2_full_adder_6.B = \multiplier_16x16bit_pipelined.layer_1_compressor42_13.cout ;
  assign \multiplier_16x16bit_pipelined.layer_2_full_adder_6.cin = \multiplier_16x16bit_pipelined.layer_1_compressor42_14.S ;
  assign \multiplier_16x16bit_pipelined.layer_2_full_adder_7.A = \multiplier_16x16bit_pipelined.layer_1_compressor42_14.carry ;
  assign \multiplier_16x16bit_pipelined.layer_2_full_adder_7.B = \multiplier_16x16bit_pipelined.layer_1_compressor42_14.cout ;
  assign \multiplier_16x16bit_pipelined.layer_2_full_adder_7.cin = \multiplier_16x16bit_pipelined.layer_1_compressor42_15.S ;
  assign \multiplier_16x16bit_pipelined.layer_2_full_adder_8.A = \multiplier_16x16bit_pipelined.layer_1_compressor42_15.carry ;
  assign \multiplier_16x16bit_pipelined.layer_2_full_adder_8.B = \multiplier_16x16bit_pipelined.layer_1_compressor42_15.cout ;
  assign \multiplier_16x16bit_pipelined.layer_2_full_adder_8.cin = \multiplier_16x16bit_pipelined.layer_1_compressor42_16.S ;
  assign \multiplier_16x16bit_pipelined.layer_2_full_adder_9.A = \multiplier_16x16bit_pipelined.layer_1_compressor42_16.carry ;
  assign \multiplier_16x16bit_pipelined.layer_2_full_adder_9.B = \multiplier_16x16bit_pipelined.layer_1_compressor42_16.cout ;
  assign \multiplier_16x16bit_pipelined.layer_2_full_adder_9.cin = \multiplier_16x16bit_pipelined.layer_1_full_adder_8.S ;
  assign \multiplier_16x16bit_pipelined.layer_2_w0 = { \multiplier_16x16bit_pipelined.mr [1], \multiplier_16x16bit_pipelined.layer_0_w0[0] };
  assign \multiplier_16x16bit_pipelined.layer_2_w1 = \multiplier_16x16bit_pipelined.layer_0_w1 ;
  assign \multiplier_16x16bit_pipelined.layer_2_w10 = { \multiplier_16x16bit_pipelined.layer_2_compressor42_0.S , \multiplier_16x16bit_pipelined.layer_2_full_adder_2.cout };
  assign \multiplier_16x16bit_pipelined.layer_2_w11 = { \multiplier_16x16bit_pipelined.layer_0_w11[5] , \multiplier_16x16bit_pipelined.layer_2_full_adder_3.S , \multiplier_16x16bit_pipelined.layer_2_compressor42_0.cout , \multiplier_16x16bit_pipelined.layer_2_compressor42_0.carry };
  assign \multiplier_16x16bit_pipelined.layer_2_w12 = { \multiplier_16x16bit_pipelined.layer_1_full_adder_3.S , \multiplier_16x16bit_pipelined.layer_2_full_adder_4.S , \multiplier_16x16bit_pipelined.layer_2_full_adder_3.cout };
  assign \multiplier_16x16bit_pipelined.layer_2_w13 = { \multiplier_16x16bit_pipelined.layer_0_w13[6] , \multiplier_16x16bit_pipelined.layer_2_compressor42_1.S , \multiplier_16x16bit_pipelined.layer_2_full_adder_4.cout };
  assign \multiplier_16x16bit_pipelined.layer_2_w14 = { \multiplier_16x16bit_pipelined.layer_2_compressor42_2.S , \multiplier_16x16bit_pipelined.layer_2_compressor42_1.cout , \multiplier_16x16bit_pipelined.layer_2_compressor42_1.carry };
  assign \multiplier_16x16bit_pipelined.layer_2_w15 = { \multiplier_16x16bit_pipelined.layer_2_compressor42_3.S , \multiplier_16x16bit_pipelined.layer_2_compressor42_2.cout , \multiplier_16x16bit_pipelined.layer_2_compressor42_2.carry };
  assign \multiplier_16x16bit_pipelined.layer_2_w16 = { \multiplier_16x16bit_pipelined.layer_2_compressor42_4.S , \multiplier_16x16bit_pipelined.layer_2_compressor42_3.cout , \multiplier_16x16bit_pipelined.layer_2_compressor42_3.carry };
  assign \multiplier_16x16bit_pipelined.layer_2_w17 = { \multiplier_16x16bit_pipelined.layer_2_compressor42_5.S , \multiplier_16x16bit_pipelined.layer_2_compressor42_4.cout , \multiplier_16x16bit_pipelined.layer_2_compressor42_4.carry };
  assign \multiplier_16x16bit_pipelined.layer_2_w18 = { \multiplier_16x16bit_pipelined.layer_0_w18[6] , \multiplier_16x16bit_pipelined.layer_2_compressor42_6.S , \multiplier_16x16bit_pipelined.layer_2_compressor42_5.cout , \multiplier_16x16bit_pipelined.layer_2_compressor42_5.carry };
  assign \multiplier_16x16bit_pipelined.layer_2_w19 = { \multiplier_16x16bit_pipelined.layer_2_compressor42_7.S , \multiplier_16x16bit_pipelined.layer_2_compressor42_6.cout , \multiplier_16x16bit_pipelined.layer_2_compressor42_6.carry };
  assign \multiplier_16x16bit_pipelined.layer_2_w2 = { \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_1.negation , \multiplier_16x16bit_pipelined.layer_0_w2[1] , \multiplier_16x16bit_pipelined.layer_0_w2[0] };
  assign \multiplier_16x16bit_pipelined.layer_2_w20 = { \multiplier_16x16bit_pipelined.layer_0_w20[5] , \multiplier_16x16bit_pipelined.layer_2_full_adder_5.S , \multiplier_16x16bit_pipelined.layer_2_compressor42_7.cout , \multiplier_16x16bit_pipelined.layer_2_compressor42_7.carry };
  assign \multiplier_16x16bit_pipelined.layer_2_w21 = { \multiplier_16x16bit_pipelined.layer_2_full_adder_6.S , \multiplier_16x16bit_pipelined.layer_2_full_adder_5.cout };
  assign \multiplier_16x16bit_pipelined.layer_2_w22 = { \multiplier_16x16bit_pipelined.layer_2_full_adder_7.S , \multiplier_16x16bit_pipelined.layer_2_full_adder_6.cout };
  assign \multiplier_16x16bit_pipelined.layer_2_w23 = { \multiplier_16x16bit_pipelined.layer_2_full_adder_8.S , \multiplier_16x16bit_pipelined.layer_2_full_adder_7.cout };
  assign \multiplier_16x16bit_pipelined.layer_2_w24 = { \multiplier_16x16bit_pipelined.layer_0_w24[3] , \multiplier_16x16bit_pipelined.layer_2_full_adder_9.S , \multiplier_16x16bit_pipelined.layer_2_full_adder_8.cout };
  assign \multiplier_16x16bit_pipelined.layer_2_w25 = { \multiplier_16x16bit_pipelined.layer_2_full_adder_10.S , \multiplier_16x16bit_pipelined.layer_2_full_adder_9.cout };
  assign \multiplier_16x16bit_pipelined.layer_2_w26 = { \multiplier_16x16bit_pipelined.layer_1_full_adder_10.S , \multiplier_16x16bit_pipelined.layer_1_full_adder_9.cout , \multiplier_16x16bit_pipelined.layer_2_full_adder_10.cout };
  assign \multiplier_16x16bit_pipelined.layer_2_w27 = { \multiplier_16x16bit_pipelined.layer_1_full_adder_11.S , \multiplier_16x16bit_pipelined.layer_1_full_adder_10.cout };
  assign \multiplier_16x16bit_pipelined.layer_2_w28 = \multiplier_16x16bit_pipelined.layer_2_full_adder_11.S ;
  assign \multiplier_16x16bit_pipelined.layer_2_w29 = { \multiplier_16x16bit_pipelined.layer_0_w29[0] , \multiplier_16x16bit_pipelined.layer_2_full_adder_11.cout };
  assign \multiplier_16x16bit_pipelined.layer_2_w3 = { \multiplier_16x16bit_pipelined.layer_0_w3[1] , \multiplier_16x16bit_pipelined.layer_0_w3[0] };
  assign \multiplier_16x16bit_pipelined.layer_2_w30 = \multiplier_16x16bit_pipelined.layer_0_w30 ;
  assign \multiplier_16x16bit_pipelined.layer_2_w4 = { \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_2.negation , \multiplier_16x16bit_pipelined.layer_1_full_adder_0.S };
  assign \multiplier_16x16bit_pipelined.layer_2_w5 = { \multiplier_16x16bit_pipelined.layer_1_full_adder_1.S , \multiplier_16x16bit_pipelined.layer_1_full_adder_0.cout };
  assign \multiplier_16x16bit_pipelined.layer_2_w6 = { \multiplier_16x16bit_pipelined.layer_1_compressor42_0.S , \multiplier_16x16bit_pipelined.layer_1_full_adder_1.cout };
  assign \multiplier_16x16bit_pipelined.layer_2_w7 = { \multiplier_16x16bit_pipelined.layer_0_w7[3] , \multiplier_16x16bit_pipelined.layer_2_full_adder_0.S };
  assign \multiplier_16x16bit_pipelined.layer_2_w8 = { \multiplier_16x16bit_pipelined.layer_2_full_adder_1.S , \multiplier_16x16bit_pipelined.layer_2_full_adder_0.cout };
  assign \multiplier_16x16bit_pipelined.layer_2_w9 = { \multiplier_16x16bit_pipelined.layer_2_full_adder_2.S , \multiplier_16x16bit_pipelined.layer_2_full_adder_1.cout };
  assign \multiplier_16x16bit_pipelined.layer_3_full_adder_0.A = \multiplier_16x16bit_pipelined.reg_layer_2_w11 [0];
  assign \multiplier_16x16bit_pipelined.layer_3_full_adder_0.B = \multiplier_16x16bit_pipelined.reg_layer_2_w11 [1];
  assign \multiplier_16x16bit_pipelined.layer_3_full_adder_0.cin = \multiplier_16x16bit_pipelined.reg_layer_2_w11 [2];
  assign \multiplier_16x16bit_pipelined.layer_3_full_adder_1.A = \multiplier_16x16bit_pipelined.reg_layer_2_w12 [0];
  assign \multiplier_16x16bit_pipelined.layer_3_full_adder_1.B = \multiplier_16x16bit_pipelined.reg_layer_2_w12 [1];
  assign \multiplier_16x16bit_pipelined.layer_3_full_adder_1.cin = \multiplier_16x16bit_pipelined.reg_layer_2_w12 [2];
  assign \multiplier_16x16bit_pipelined.layer_3_full_adder_10.A = \multiplier_16x16bit_pipelined.reg_layer_2_w21 [0];
  assign \multiplier_16x16bit_pipelined.layer_3_full_adder_10.B = \multiplier_16x16bit_pipelined.reg_layer_2_w21 [1];
  assign \multiplier_16x16bit_pipelined.layer_3_full_adder_10.cin = \multiplier_16x16bit_pipelined.reg_layer_2_w21 [2];
  assign \multiplier_16x16bit_pipelined.layer_3_full_adder_11.A = \multiplier_16x16bit_pipelined.reg_layer_2_w24 [0];
  assign \multiplier_16x16bit_pipelined.layer_3_full_adder_11.B = \multiplier_16x16bit_pipelined.reg_layer_2_w24 [1];
  assign \multiplier_16x16bit_pipelined.layer_3_full_adder_11.S = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_24.B ;
  assign \multiplier_16x16bit_pipelined.layer_3_full_adder_11.cin = \multiplier_16x16bit_pipelined.reg_layer_2_w24 [2];
  assign \multiplier_16x16bit_pipelined.layer_3_full_adder_12.A = \multiplier_16x16bit_pipelined.reg_layer_2_w26 [0];
  assign \multiplier_16x16bit_pipelined.layer_3_full_adder_12.B = \multiplier_16x16bit_pipelined.reg_layer_2_w26 [1];
  assign \multiplier_16x16bit_pipelined.layer_3_full_adder_12.S = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_26.B ;
  assign \multiplier_16x16bit_pipelined.layer_3_full_adder_12.cin = \multiplier_16x16bit_pipelined.reg_layer_2_w26 [2];
  assign \multiplier_16x16bit_pipelined.layer_3_full_adder_13.A = \multiplier_16x16bit_pipelined.reg_layer_2_w29 [0];
  assign \multiplier_16x16bit_pipelined.layer_3_full_adder_13.B = \multiplier_16x16bit_pipelined.reg_layer_2_w29 [1];
  assign \multiplier_16x16bit_pipelined.layer_3_full_adder_13.S = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_29.A ;
  assign \multiplier_16x16bit_pipelined.layer_3_full_adder_13.cin = \multiplier_16x16bit_pipelined.reg_layer_2_w29 [2];
  assign \multiplier_16x16bit_pipelined.layer_3_full_adder_13.cout = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_30.A ;
  assign \multiplier_16x16bit_pipelined.layer_3_full_adder_2.A = \multiplier_16x16bit_pipelined.reg_layer_2_w13 [0];
  assign \multiplier_16x16bit_pipelined.layer_3_full_adder_2.B = \multiplier_16x16bit_pipelined.reg_layer_2_w13 [1];
  assign \multiplier_16x16bit_pipelined.layer_3_full_adder_2.cin = \multiplier_16x16bit_pipelined.reg_layer_2_w13 [2];
  assign \multiplier_16x16bit_pipelined.layer_3_full_adder_3.A = \multiplier_16x16bit_pipelined.reg_layer_2_w14 [0];
  assign \multiplier_16x16bit_pipelined.layer_3_full_adder_3.B = \multiplier_16x16bit_pipelined.reg_layer_2_w14 [1];
  assign \multiplier_16x16bit_pipelined.layer_3_full_adder_3.cin = \multiplier_16x16bit_pipelined.reg_layer_2_w14 [2];
  assign \multiplier_16x16bit_pipelined.layer_3_full_adder_4.A = \multiplier_16x16bit_pipelined.reg_layer_2_w15 [0];
  assign \multiplier_16x16bit_pipelined.layer_3_full_adder_4.B = \multiplier_16x16bit_pipelined.reg_layer_2_w15 [1];
  assign \multiplier_16x16bit_pipelined.layer_3_full_adder_4.cin = \multiplier_16x16bit_pipelined.reg_layer_2_w15 [2];
  assign \multiplier_16x16bit_pipelined.layer_3_full_adder_5.A = \multiplier_16x16bit_pipelined.reg_layer_2_w16 [0];
  assign \multiplier_16x16bit_pipelined.layer_3_full_adder_5.B = \multiplier_16x16bit_pipelined.reg_layer_2_w16 [1];
  assign \multiplier_16x16bit_pipelined.layer_3_full_adder_5.cin = \multiplier_16x16bit_pipelined.reg_layer_2_w16 [2];
  assign \multiplier_16x16bit_pipelined.layer_3_full_adder_6.A = \multiplier_16x16bit_pipelined.reg_layer_2_w17 [0];
  assign \multiplier_16x16bit_pipelined.layer_3_full_adder_6.B = \multiplier_16x16bit_pipelined.reg_layer_2_w17 [1];
  assign \multiplier_16x16bit_pipelined.layer_3_full_adder_6.cin = \multiplier_16x16bit_pipelined.reg_layer_2_w17 [2];
  assign \multiplier_16x16bit_pipelined.layer_3_full_adder_7.A = \multiplier_16x16bit_pipelined.reg_layer_2_w18 [0];
  assign \multiplier_16x16bit_pipelined.layer_3_full_adder_7.B = \multiplier_16x16bit_pipelined.reg_layer_2_w18 [1];
  assign \multiplier_16x16bit_pipelined.layer_3_full_adder_7.cin = \multiplier_16x16bit_pipelined.reg_layer_2_w18 [2];
  assign \multiplier_16x16bit_pipelined.layer_3_full_adder_8.A = \multiplier_16x16bit_pipelined.reg_layer_2_w19 [0];
  assign \multiplier_16x16bit_pipelined.layer_3_full_adder_8.B = \multiplier_16x16bit_pipelined.reg_layer_2_w19 [1];
  assign \multiplier_16x16bit_pipelined.layer_3_full_adder_8.cin = \multiplier_16x16bit_pipelined.reg_layer_2_w19 [2];
  assign \multiplier_16x16bit_pipelined.layer_3_full_adder_9.A = \multiplier_16x16bit_pipelined.reg_layer_2_w20 [0];
  assign \multiplier_16x16bit_pipelined.layer_3_full_adder_9.B = \multiplier_16x16bit_pipelined.reg_layer_2_w20 [1];
  assign \multiplier_16x16bit_pipelined.layer_3_full_adder_9.cin = \multiplier_16x16bit_pipelined.reg_layer_2_w20 [2];
  assign \multiplier_16x16bit_pipelined.layer_3_w0[0] = \multiplier_16x16bit_pipelined.reg_layer_2_w0 [0];
  assign \multiplier_16x16bit_pipelined.layer_3_w0[1] = \multiplier_16x16bit_pipelined.reg_layer_2_w0 [1];
  assign \multiplier_16x16bit_pipelined.layer_3_w1 = \multiplier_16x16bit_pipelined.reg_layer_2_w1 ;
  assign \multiplier_16x16bit_pipelined.layer_3_w10[0] = \multiplier_16x16bit_pipelined.reg_layer_2_w10 [0];
  assign \multiplier_16x16bit_pipelined.layer_3_w10[1] = \multiplier_16x16bit_pipelined.reg_layer_2_w10 [1];
  assign \multiplier_16x16bit_pipelined.layer_3_w11[0] = \multiplier_16x16bit_pipelined.layer_3_full_adder_0.S ;
  assign \multiplier_16x16bit_pipelined.layer_3_w11[1] = \multiplier_16x16bit_pipelined.reg_layer_2_w11 [3];
  assign \multiplier_16x16bit_pipelined.layer_3_w12[0] = \multiplier_16x16bit_pipelined.layer_3_full_adder_0.cout ;
  assign \multiplier_16x16bit_pipelined.layer_3_w12[1] = \multiplier_16x16bit_pipelined.layer_3_full_adder_1.S ;
  assign \multiplier_16x16bit_pipelined.layer_3_w13[0] = \multiplier_16x16bit_pipelined.layer_3_full_adder_1.cout ;
  assign \multiplier_16x16bit_pipelined.layer_3_w13[1] = \multiplier_16x16bit_pipelined.layer_3_full_adder_2.S ;
  assign \multiplier_16x16bit_pipelined.layer_3_w14[0] = \multiplier_16x16bit_pipelined.layer_3_full_adder_2.cout ;
  assign \multiplier_16x16bit_pipelined.layer_3_w14[1] = \multiplier_16x16bit_pipelined.layer_3_full_adder_3.S ;
  assign \multiplier_16x16bit_pipelined.layer_3_w15[0] = \multiplier_16x16bit_pipelined.layer_3_full_adder_3.cout ;
  assign \multiplier_16x16bit_pipelined.layer_3_w15[1] = \multiplier_16x16bit_pipelined.layer_3_full_adder_4.S ;
  assign \multiplier_16x16bit_pipelined.layer_3_w16[0] = \multiplier_16x16bit_pipelined.layer_3_full_adder_4.cout ;
  assign \multiplier_16x16bit_pipelined.layer_3_w16[1] = \multiplier_16x16bit_pipelined.layer_3_full_adder_5.S ;
  assign \multiplier_16x16bit_pipelined.layer_3_w16[2] = \multiplier_16x16bit_pipelined.reg_layer_2_w16 [3];
  assign \multiplier_16x16bit_pipelined.layer_3_w17[0] = \multiplier_16x16bit_pipelined.layer_3_full_adder_5.cout ;
  assign \multiplier_16x16bit_pipelined.layer_3_w17[1] = \multiplier_16x16bit_pipelined.layer_3_full_adder_6.S ;
  assign \multiplier_16x16bit_pipelined.layer_3_w18[0] = \multiplier_16x16bit_pipelined.layer_3_full_adder_6.cout ;
  assign \multiplier_16x16bit_pipelined.layer_3_w18[1] = \multiplier_16x16bit_pipelined.layer_3_full_adder_7.S ;
  assign \multiplier_16x16bit_pipelined.layer_3_w18[2] = \multiplier_16x16bit_pipelined.reg_layer_2_w18 [3];
  assign \multiplier_16x16bit_pipelined.layer_3_w19[0] = \multiplier_16x16bit_pipelined.layer_3_full_adder_7.cout ;
  assign \multiplier_16x16bit_pipelined.layer_3_w19[1] = \multiplier_16x16bit_pipelined.layer_3_full_adder_8.S ;
  assign \multiplier_16x16bit_pipelined.layer_3_w20[0] = \multiplier_16x16bit_pipelined.layer_3_full_adder_8.cout ;
  assign \multiplier_16x16bit_pipelined.layer_3_w20[1] = \multiplier_16x16bit_pipelined.layer_3_full_adder_9.S ;
  assign \multiplier_16x16bit_pipelined.layer_3_w20[2] = \multiplier_16x16bit_pipelined.reg_layer_2_w20 [3];
  assign \multiplier_16x16bit_pipelined.layer_3_w21[0] = \multiplier_16x16bit_pipelined.layer_3_full_adder_9.cout ;
  assign \multiplier_16x16bit_pipelined.layer_3_w21[1] = \multiplier_16x16bit_pipelined.layer_3_full_adder_10.S ;
  assign \multiplier_16x16bit_pipelined.layer_3_w22[0] = \multiplier_16x16bit_pipelined.layer_3_full_adder_10.cout ;
  assign \multiplier_16x16bit_pipelined.layer_3_w22[1] = \multiplier_16x16bit_pipelined.reg_layer_2_w22 [0];
  assign \multiplier_16x16bit_pipelined.layer_3_w22[2] = \multiplier_16x16bit_pipelined.reg_layer_2_w22 [1];
  assign \multiplier_16x16bit_pipelined.layer_3_w23[0] = \multiplier_16x16bit_pipelined.reg_layer_2_w23 [0];
  assign \multiplier_16x16bit_pipelined.layer_3_w23[1] = \multiplier_16x16bit_pipelined.reg_layer_2_w23 [1];
  assign \multiplier_16x16bit_pipelined.layer_3_w24 = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_24.B ;
  assign \multiplier_16x16bit_pipelined.layer_3_w25[0] = \multiplier_16x16bit_pipelined.layer_3_full_adder_11.cout ;
  assign \multiplier_16x16bit_pipelined.layer_3_w25[1] = \multiplier_16x16bit_pipelined.reg_layer_2_w25 [0];
  assign \multiplier_16x16bit_pipelined.layer_3_w25[2] = \multiplier_16x16bit_pipelined.reg_layer_2_w25 [1];
  assign \multiplier_16x16bit_pipelined.layer_3_w26 = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_26.B ;
  assign \multiplier_16x16bit_pipelined.layer_3_w27[0] = \multiplier_16x16bit_pipelined.layer_3_full_adder_12.cout ;
  assign \multiplier_16x16bit_pipelined.layer_3_w27[1] = \multiplier_16x16bit_pipelined.reg_layer_2_w27 [0];
  assign \multiplier_16x16bit_pipelined.layer_3_w27[2] = \multiplier_16x16bit_pipelined.reg_layer_2_w27 [1];
  assign \multiplier_16x16bit_pipelined.layer_3_w28 = \multiplier_16x16bit_pipelined.reg_layer_2_w28 ;
  assign \multiplier_16x16bit_pipelined.layer_3_w29 = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_29.A ;
  assign \multiplier_16x16bit_pipelined.layer_3_w2[0] = \multiplier_16x16bit_pipelined.reg_layer_2_w2 [0];
  assign \multiplier_16x16bit_pipelined.layer_3_w2[1] = \multiplier_16x16bit_pipelined.reg_layer_2_w2 [1];
  assign \multiplier_16x16bit_pipelined.layer_3_w2[2] = \multiplier_16x16bit_pipelined.reg_layer_2_w2 [2];
  assign \multiplier_16x16bit_pipelined.layer_3_w30[0] = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_30.A ;
  assign \multiplier_16x16bit_pipelined.layer_3_w30[1] = \multiplier_16x16bit_pipelined.reg_layer_2_w30 ;
  assign \multiplier_16x16bit_pipelined.layer_3_w31 = \multiplier_16x16bit_pipelined.reg_layer_2_w31 ;
  assign \multiplier_16x16bit_pipelined.layer_3_w3[0] = \multiplier_16x16bit_pipelined.reg_layer_2_w3 [0];
  assign \multiplier_16x16bit_pipelined.layer_3_w3[1] = \multiplier_16x16bit_pipelined.reg_layer_2_w3 [1];
  assign \multiplier_16x16bit_pipelined.layer_3_w4[0] = \multiplier_16x16bit_pipelined.reg_layer_2_w4 [0];
  assign \multiplier_16x16bit_pipelined.layer_3_w4[1] = \multiplier_16x16bit_pipelined.reg_layer_2_w4 [1];
  assign \multiplier_16x16bit_pipelined.layer_3_w5[0] = \multiplier_16x16bit_pipelined.reg_layer_2_w5 [0];
  assign \multiplier_16x16bit_pipelined.layer_3_w5[1] = \multiplier_16x16bit_pipelined.reg_layer_2_w5 [1];
  assign \multiplier_16x16bit_pipelined.layer_3_w6[0] = \multiplier_16x16bit_pipelined.reg_layer_2_w6 [0];
  assign \multiplier_16x16bit_pipelined.layer_3_w6[1] = \multiplier_16x16bit_pipelined.reg_layer_2_w6 [1];
  assign \multiplier_16x16bit_pipelined.layer_3_w7[0] = \multiplier_16x16bit_pipelined.reg_layer_2_w7 [0];
  assign \multiplier_16x16bit_pipelined.layer_3_w7[1] = \multiplier_16x16bit_pipelined.reg_layer_2_w7 [1];
  assign \multiplier_16x16bit_pipelined.layer_3_w8[0] = \multiplier_16x16bit_pipelined.reg_layer_2_w8 [0];
  assign \multiplier_16x16bit_pipelined.layer_3_w8[1] = \multiplier_16x16bit_pipelined.reg_layer_2_w8 [1];
  assign \multiplier_16x16bit_pipelined.layer_3_w9[0] = \multiplier_16x16bit_pipelined.reg_layer_2_w9 [0];
  assign \multiplier_16x16bit_pipelined.layer_3_w9[1] = \multiplier_16x16bit_pipelined.reg_layer_2_w9 [1];
  assign \multiplier_16x16bit_pipelined.layer_4_full_adder_0.A = \multiplier_16x16bit_pipelined.reg_layer_2_w2 [0];
  assign \multiplier_16x16bit_pipelined.layer_4_full_adder_0.B = \multiplier_16x16bit_pipelined.reg_layer_2_w2 [1];
  assign \multiplier_16x16bit_pipelined.layer_4_full_adder_0.S = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_2.A ;
  assign \multiplier_16x16bit_pipelined.layer_4_full_adder_0.cin = \multiplier_16x16bit_pipelined.reg_layer_2_w2 [2];
  assign \multiplier_16x16bit_pipelined.layer_4_full_adder_0.cout = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_3.A ;
  assign \multiplier_16x16bit_pipelined.layer_4_full_adder_1.A = \multiplier_16x16bit_pipelined.layer_3_full_adder_4.cout ;
  assign \multiplier_16x16bit_pipelined.layer_4_full_adder_1.B = \multiplier_16x16bit_pipelined.layer_3_full_adder_5.S ;
  assign \multiplier_16x16bit_pipelined.layer_4_full_adder_1.S = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_16.B ;
  assign \multiplier_16x16bit_pipelined.layer_4_full_adder_1.cin = \multiplier_16x16bit_pipelined.reg_layer_2_w16 [3];
  assign \multiplier_16x16bit_pipelined.layer_4_full_adder_1.cout = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_17.A ;
  assign \multiplier_16x16bit_pipelined.layer_4_full_adder_2.A = \multiplier_16x16bit_pipelined.layer_3_full_adder_6.cout ;
  assign \multiplier_16x16bit_pipelined.layer_4_full_adder_2.B = \multiplier_16x16bit_pipelined.layer_3_full_adder_7.S ;
  assign \multiplier_16x16bit_pipelined.layer_4_full_adder_2.S = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_18.B ;
  assign \multiplier_16x16bit_pipelined.layer_4_full_adder_2.cin = \multiplier_16x16bit_pipelined.reg_layer_2_w18 [3];
  assign \multiplier_16x16bit_pipelined.layer_4_full_adder_2.cout = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_19.A ;
  assign \multiplier_16x16bit_pipelined.layer_4_full_adder_3.A = \multiplier_16x16bit_pipelined.layer_3_full_adder_8.cout ;
  assign \multiplier_16x16bit_pipelined.layer_4_full_adder_3.B = \multiplier_16x16bit_pipelined.layer_3_full_adder_9.S ;
  assign \multiplier_16x16bit_pipelined.layer_4_full_adder_3.S = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_20.B ;
  assign \multiplier_16x16bit_pipelined.layer_4_full_adder_3.cin = \multiplier_16x16bit_pipelined.reg_layer_2_w20 [3];
  assign \multiplier_16x16bit_pipelined.layer_4_full_adder_3.cout = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_21.A ;
  assign \multiplier_16x16bit_pipelined.layer_4_full_adder_4.A = \multiplier_16x16bit_pipelined.layer_3_full_adder_10.cout ;
  assign \multiplier_16x16bit_pipelined.layer_4_full_adder_4.B = \multiplier_16x16bit_pipelined.reg_layer_2_w22 [0];
  assign \multiplier_16x16bit_pipelined.layer_4_full_adder_4.S = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_22.B ;
  assign \multiplier_16x16bit_pipelined.layer_4_full_adder_4.cin = \multiplier_16x16bit_pipelined.reg_layer_2_w22 [1];
  assign \multiplier_16x16bit_pipelined.layer_4_full_adder_4.cout = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_23.A ;
  assign \multiplier_16x16bit_pipelined.layer_4_full_adder_5.A = \multiplier_16x16bit_pipelined.layer_3_full_adder_11.cout ;
  assign \multiplier_16x16bit_pipelined.layer_4_full_adder_5.B = \multiplier_16x16bit_pipelined.reg_layer_2_w25 [0];
  assign \multiplier_16x16bit_pipelined.layer_4_full_adder_5.S = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_25.A ;
  assign \multiplier_16x16bit_pipelined.layer_4_full_adder_5.cin = \multiplier_16x16bit_pipelined.reg_layer_2_w25 [1];
  assign \multiplier_16x16bit_pipelined.layer_4_full_adder_5.cout = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_26.A ;
  assign \multiplier_16x16bit_pipelined.layer_4_full_adder_6.A = \multiplier_16x16bit_pipelined.layer_3_full_adder_12.cout ;
  assign \multiplier_16x16bit_pipelined.layer_4_full_adder_6.B = \multiplier_16x16bit_pipelined.reg_layer_2_w27 [0];
  assign \multiplier_16x16bit_pipelined.layer_4_full_adder_6.S = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_27.A ;
  assign \multiplier_16x16bit_pipelined.layer_4_full_adder_6.cin = \multiplier_16x16bit_pipelined.reg_layer_2_w27 [1];
  assign \multiplier_16x16bit_pipelined.layer_4_full_adder_6.cout = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_28.A ;
  assign \multiplier_16x16bit_pipelined.layer_4_half_adder_0.A = \multiplier_16x16bit_pipelined.reg_layer_2_w3 [0];
  assign \multiplier_16x16bit_pipelined.layer_4_half_adder_0.B = \multiplier_16x16bit_pipelined.reg_layer_2_w3 [1];
  assign \multiplier_16x16bit_pipelined.layer_4_half_adder_0.S = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_3.B ;
  assign \multiplier_16x16bit_pipelined.layer_4_half_adder_0.carry = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_4.A ;
  assign \multiplier_16x16bit_pipelined.layer_4_half_adder_1.A = \multiplier_16x16bit_pipelined.reg_layer_2_w4 [0];
  assign \multiplier_16x16bit_pipelined.layer_4_half_adder_1.B = \multiplier_16x16bit_pipelined.reg_layer_2_w4 [1];
  assign \multiplier_16x16bit_pipelined.layer_4_half_adder_1.S = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_4.B ;
  assign \multiplier_16x16bit_pipelined.layer_4_half_adder_1.carry = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_5.A ;
  assign \multiplier_16x16bit_pipelined.layer_4_half_adder_10.A = \multiplier_16x16bit_pipelined.layer_3_full_adder_1.cout ;
  assign \multiplier_16x16bit_pipelined.layer_4_half_adder_10.B = \multiplier_16x16bit_pipelined.layer_3_full_adder_2.S ;
  assign \multiplier_16x16bit_pipelined.layer_4_half_adder_10.S = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_13.B ;
  assign \multiplier_16x16bit_pipelined.layer_4_half_adder_10.carry = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_14.A ;
  assign \multiplier_16x16bit_pipelined.layer_4_half_adder_11.A = \multiplier_16x16bit_pipelined.layer_3_full_adder_2.cout ;
  assign \multiplier_16x16bit_pipelined.layer_4_half_adder_11.B = \multiplier_16x16bit_pipelined.layer_3_full_adder_3.S ;
  assign \multiplier_16x16bit_pipelined.layer_4_half_adder_11.S = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_14.B ;
  assign \multiplier_16x16bit_pipelined.layer_4_half_adder_11.carry = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_15.A ;
  assign \multiplier_16x16bit_pipelined.layer_4_half_adder_12.A = \multiplier_16x16bit_pipelined.layer_3_full_adder_3.cout ;
  assign \multiplier_16x16bit_pipelined.layer_4_half_adder_12.B = \multiplier_16x16bit_pipelined.layer_3_full_adder_4.S ;
  assign \multiplier_16x16bit_pipelined.layer_4_half_adder_12.S = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_15.B ;
  assign \multiplier_16x16bit_pipelined.layer_4_half_adder_12.carry = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_16.A ;
  assign \multiplier_16x16bit_pipelined.layer_4_half_adder_13.A = \multiplier_16x16bit_pipelined.layer_3_full_adder_5.cout ;
  assign \multiplier_16x16bit_pipelined.layer_4_half_adder_13.B = \multiplier_16x16bit_pipelined.layer_3_full_adder_6.S ;
  assign \multiplier_16x16bit_pipelined.layer_4_half_adder_13.S = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_17.B ;
  assign \multiplier_16x16bit_pipelined.layer_4_half_adder_13.carry = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_18.A ;
  assign \multiplier_16x16bit_pipelined.layer_4_half_adder_14.A = \multiplier_16x16bit_pipelined.layer_3_full_adder_7.cout ;
  assign \multiplier_16x16bit_pipelined.layer_4_half_adder_14.B = \multiplier_16x16bit_pipelined.layer_3_full_adder_8.S ;
  assign \multiplier_16x16bit_pipelined.layer_4_half_adder_14.S = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_19.B ;
  assign \multiplier_16x16bit_pipelined.layer_4_half_adder_14.carry = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_20.A ;
  assign \multiplier_16x16bit_pipelined.layer_4_half_adder_15.A = \multiplier_16x16bit_pipelined.layer_3_full_adder_9.cout ;
  assign \multiplier_16x16bit_pipelined.layer_4_half_adder_15.B = \multiplier_16x16bit_pipelined.layer_3_full_adder_10.S ;
  assign \multiplier_16x16bit_pipelined.layer_4_half_adder_15.S = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_21.B ;
  assign \multiplier_16x16bit_pipelined.layer_4_half_adder_15.carry = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_22.A ;
  assign \multiplier_16x16bit_pipelined.layer_4_half_adder_16.A = \multiplier_16x16bit_pipelined.reg_layer_2_w23 [0];
  assign \multiplier_16x16bit_pipelined.layer_4_half_adder_16.B = \multiplier_16x16bit_pipelined.reg_layer_2_w23 [1];
  assign \multiplier_16x16bit_pipelined.layer_4_half_adder_16.S = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_23.B ;
  assign \multiplier_16x16bit_pipelined.layer_4_half_adder_16.carry = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_24.A ;
  assign \multiplier_16x16bit_pipelined.layer_4_half_adder_2.A = \multiplier_16x16bit_pipelined.reg_layer_2_w5 [0];
  assign \multiplier_16x16bit_pipelined.layer_4_half_adder_2.B = \multiplier_16x16bit_pipelined.reg_layer_2_w5 [1];
  assign \multiplier_16x16bit_pipelined.layer_4_half_adder_2.S = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_5.B ;
  assign \multiplier_16x16bit_pipelined.layer_4_half_adder_2.carry = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_6.A ;
  assign \multiplier_16x16bit_pipelined.layer_4_half_adder_3.A = \multiplier_16x16bit_pipelined.reg_layer_2_w6 [0];
  assign \multiplier_16x16bit_pipelined.layer_4_half_adder_3.B = \multiplier_16x16bit_pipelined.reg_layer_2_w6 [1];
  assign \multiplier_16x16bit_pipelined.layer_4_half_adder_3.S = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_6.B ;
  assign \multiplier_16x16bit_pipelined.layer_4_half_adder_3.carry = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_7.A ;
  assign \multiplier_16x16bit_pipelined.layer_4_half_adder_4.A = \multiplier_16x16bit_pipelined.reg_layer_2_w7 [0];
  assign \multiplier_16x16bit_pipelined.layer_4_half_adder_4.B = \multiplier_16x16bit_pipelined.reg_layer_2_w7 [1];
  assign \multiplier_16x16bit_pipelined.layer_4_half_adder_4.S = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_7.B ;
  assign \multiplier_16x16bit_pipelined.layer_4_half_adder_4.carry = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_8.A ;
  assign \multiplier_16x16bit_pipelined.layer_4_half_adder_5.A = \multiplier_16x16bit_pipelined.reg_layer_2_w8 [0];
  assign \multiplier_16x16bit_pipelined.layer_4_half_adder_5.B = \multiplier_16x16bit_pipelined.reg_layer_2_w8 [1];
  assign \multiplier_16x16bit_pipelined.layer_4_half_adder_5.S = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_8.B ;
  assign \multiplier_16x16bit_pipelined.layer_4_half_adder_5.carry = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_9.A ;
  assign \multiplier_16x16bit_pipelined.layer_4_half_adder_6.A = \multiplier_16x16bit_pipelined.reg_layer_2_w9 [0];
  assign \multiplier_16x16bit_pipelined.layer_4_half_adder_6.B = \multiplier_16x16bit_pipelined.reg_layer_2_w9 [1];
  assign \multiplier_16x16bit_pipelined.layer_4_half_adder_6.S = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_9.B ;
  assign \multiplier_16x16bit_pipelined.layer_4_half_adder_6.carry = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_10.A ;
  assign \multiplier_16x16bit_pipelined.layer_4_half_adder_7.A = \multiplier_16x16bit_pipelined.reg_layer_2_w10 [0];
  assign \multiplier_16x16bit_pipelined.layer_4_half_adder_7.B = \multiplier_16x16bit_pipelined.reg_layer_2_w10 [1];
  assign \multiplier_16x16bit_pipelined.layer_4_half_adder_7.S = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_10.B ;
  assign \multiplier_16x16bit_pipelined.layer_4_half_adder_7.carry = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_11.A ;
  assign \multiplier_16x16bit_pipelined.layer_4_half_adder_8.A = \multiplier_16x16bit_pipelined.layer_3_full_adder_0.S ;
  assign \multiplier_16x16bit_pipelined.layer_4_half_adder_8.B = \multiplier_16x16bit_pipelined.reg_layer_2_w11 [3];
  assign \multiplier_16x16bit_pipelined.layer_4_half_adder_8.S = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_11.B ;
  assign \multiplier_16x16bit_pipelined.layer_4_half_adder_8.carry = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_12.A ;
  assign \multiplier_16x16bit_pipelined.layer_4_half_adder_9.A = \multiplier_16x16bit_pipelined.layer_3_full_adder_0.cout ;
  assign \multiplier_16x16bit_pipelined.layer_4_half_adder_9.B = \multiplier_16x16bit_pipelined.layer_3_full_adder_1.S ;
  assign \multiplier_16x16bit_pipelined.layer_4_half_adder_9.S = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_12.B ;
  assign \multiplier_16x16bit_pipelined.layer_4_half_adder_9.carry = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_13.A ;
  assign \multiplier_16x16bit_pipelined.layer_4_w0[0] = \multiplier_16x16bit_pipelined.reg_layer_2_w0 [0];
  assign \multiplier_16x16bit_pipelined.layer_4_w0[1] = \multiplier_16x16bit_pipelined.reg_layer_2_w0 [1];
  assign \multiplier_16x16bit_pipelined.layer_4_w1 = \multiplier_16x16bit_pipelined.reg_layer_2_w1 ;
  assign \multiplier_16x16bit_pipelined.layer_4_w10[0] = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_10.A ;
  assign \multiplier_16x16bit_pipelined.layer_4_w10[1] = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_10.B ;
  assign \multiplier_16x16bit_pipelined.layer_4_w11[0] = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_11.A ;
  assign \multiplier_16x16bit_pipelined.layer_4_w11[1] = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_11.B ;
  assign \multiplier_16x16bit_pipelined.layer_4_w12[0] = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_12.A ;
  assign \multiplier_16x16bit_pipelined.layer_4_w12[1] = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_12.B ;
  assign \multiplier_16x16bit_pipelined.layer_4_w13[0] = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_13.A ;
  assign \multiplier_16x16bit_pipelined.layer_4_w13[1] = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_13.B ;
  assign \multiplier_16x16bit_pipelined.layer_4_w14[0] = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_14.A ;
  assign \multiplier_16x16bit_pipelined.layer_4_w14[1] = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_14.B ;
  assign \multiplier_16x16bit_pipelined.layer_4_w15[0] = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_15.A ;
  assign \multiplier_16x16bit_pipelined.layer_4_w15[1] = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_15.B ;
  assign \multiplier_16x16bit_pipelined.layer_4_w16[0] = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_16.A ;
  assign \multiplier_16x16bit_pipelined.layer_4_w16[1] = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_16.B ;
  assign \multiplier_16x16bit_pipelined.layer_4_w17[0] = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_17.A ;
  assign \multiplier_16x16bit_pipelined.layer_4_w17[1] = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_17.B ;
  assign \multiplier_16x16bit_pipelined.layer_4_w18[0] = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_18.A ;
  assign \multiplier_16x16bit_pipelined.layer_4_w18[1] = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_18.B ;
  assign \multiplier_16x16bit_pipelined.layer_4_w19[0] = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_19.A ;
  assign \multiplier_16x16bit_pipelined.layer_4_w19[1] = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_19.B ;
  assign \multiplier_16x16bit_pipelined.layer_4_w2 = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_2.A ;
  assign \multiplier_16x16bit_pipelined.layer_4_w20[0] = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_20.A ;
  assign \multiplier_16x16bit_pipelined.layer_4_w20[1] = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_20.B ;
  assign \multiplier_16x16bit_pipelined.layer_4_w21[0] = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_21.A ;
  assign \multiplier_16x16bit_pipelined.layer_4_w21[1] = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_21.B ;
  assign \multiplier_16x16bit_pipelined.layer_4_w22[0] = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_22.A ;
  assign \multiplier_16x16bit_pipelined.layer_4_w22[1] = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_22.B ;
  assign \multiplier_16x16bit_pipelined.layer_4_w23[0] = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_23.A ;
  assign \multiplier_16x16bit_pipelined.layer_4_w23[1] = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_23.B ;
  assign \multiplier_16x16bit_pipelined.layer_4_w24[0] = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_24.A ;
  assign \multiplier_16x16bit_pipelined.layer_4_w24[1] = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_24.B ;
  assign \multiplier_16x16bit_pipelined.layer_4_w25 = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_25.A ;
  assign \multiplier_16x16bit_pipelined.layer_4_w26[0] = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_26.A ;
  assign \multiplier_16x16bit_pipelined.layer_4_w26[1] = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_26.B ;
  assign \multiplier_16x16bit_pipelined.layer_4_w27 = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_27.A ;
  assign \multiplier_16x16bit_pipelined.layer_4_w28[0] = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_28.A ;
  assign \multiplier_16x16bit_pipelined.layer_4_w28[1] = \multiplier_16x16bit_pipelined.reg_layer_2_w28 ;
  assign \multiplier_16x16bit_pipelined.layer_4_w29 = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_29.A ;
  assign \multiplier_16x16bit_pipelined.layer_4_w30[0] = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_30.A ;
  assign \multiplier_16x16bit_pipelined.layer_4_w30[1] = \multiplier_16x16bit_pipelined.reg_layer_2_w30 ;
  assign \multiplier_16x16bit_pipelined.layer_4_w31 = \multiplier_16x16bit_pipelined.reg_layer_2_w31 ;
  assign \multiplier_16x16bit_pipelined.layer_4_w3[0] = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_3.A ;
  assign \multiplier_16x16bit_pipelined.layer_4_w3[1] = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_3.B ;
  assign \multiplier_16x16bit_pipelined.layer_4_w4[0] = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_4.A ;
  assign \multiplier_16x16bit_pipelined.layer_4_w4[1] = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_4.B ;
  assign \multiplier_16x16bit_pipelined.layer_4_w5[0] = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_5.A ;
  assign \multiplier_16x16bit_pipelined.layer_4_w5[1] = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_5.B ;
  assign \multiplier_16x16bit_pipelined.layer_4_w6[0] = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_6.A ;
  assign \multiplier_16x16bit_pipelined.layer_4_w6[1] = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_6.B ;
  assign \multiplier_16x16bit_pipelined.layer_4_w7[0] = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_7.A ;
  assign \multiplier_16x16bit_pipelined.layer_4_w7[1] = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_7.B ;
  assign \multiplier_16x16bit_pipelined.layer_4_w8[0] = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_8.A ;
  assign \multiplier_16x16bit_pipelined.layer_4_w8[1] = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_8.B ;
  assign \multiplier_16x16bit_pipelined.layer_4_w9[0] = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_9.A ;
  assign \multiplier_16x16bit_pipelined.layer_4_w9[1] = \multiplier_16x16bit_pipelined.adder_32bit.operator_A_9.B ;
  assign \multiplier_16x16bit_pipelined.negation = { \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_7.negation , \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_6.negation , \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_5.negation , \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_4.negation , \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_3.negation , \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_2.negation , \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_1.negation , \multiplier_16x16bit_pipelined.mr [1] };
  assign \multiplier_16x16bit_pipelined.o_product = { \multiplier_16x16bit_pipelined.adder_32bit.o_s [31:1], \multiplier_16x16bit_pipelined.adder_32bit.operator_A_0.P };
  assign \multiplier_16x16bit_pipelined.partial_product_gen_0.double = \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_0.double ;
  assign \multiplier_16x16bit_pipelined.partial_product_gen_0.md = \multiplier_16x16bit_pipelined.md ;
  assign \multiplier_16x16bit_pipelined.partial_product_gen_0.negation = \multiplier_16x16bit_pipelined.mr [1];
  assign \multiplier_16x16bit_pipelined.partial_product_gen_0.pp = { \multiplier_16x16bit_pipelined.layer_1_compressor42_9.A , \multiplier_16x16bit_pipelined.layer_1_compressor42_8.A , \multiplier_16x16bit_pipelined.layer_1_compressor42_7.A , \multiplier_16x16bit_pipelined.layer_1_compressor42_6.A , \multiplier_16x16bit_pipelined.layer_1_compressor42_5.A , \multiplier_16x16bit_pipelined.layer_1_compressor42_4.A , \multiplier_16x16bit_pipelined.layer_1_compressor42_3.A , \multiplier_16x16bit_pipelined.layer_1_compressor42_2.A , \multiplier_16x16bit_pipelined.layer_1_compressor42_1.A , \multiplier_16x16bit_pipelined.layer_1_full_adder_2.A , \multiplier_16x16bit_pipelined.layer_1_compressor42_0.A , \multiplier_16x16bit_pipelined.layer_1_full_adder_1.A , \multiplier_16x16bit_pipelined.layer_1_full_adder_0.A , \multiplier_16x16bit_pipelined.layer_0_w3[0] , \multiplier_16x16bit_pipelined.layer_0_w2[0] , \multiplier_16x16bit_pipelined.layer_0_w1 , \multiplier_16x16bit_pipelined.layer_0_w0[0] };
  assign \multiplier_16x16bit_pipelined.partial_product_gen_0.zero = \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_0.zero ;
  assign \multiplier_16x16bit_pipelined.partial_product_gen_1.double = \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_1.double ;
  assign \multiplier_16x16bit_pipelined.partial_product_gen_1.md = \multiplier_16x16bit_pipelined.md ;
  assign \multiplier_16x16bit_pipelined.partial_product_gen_1.negation = \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_1.negation ;
  assign \multiplier_16x16bit_pipelined.partial_product_gen_1.pp = { \multiplier_16x16bit_pipelined.layer_1_compressor42_11.A , \multiplier_16x16bit_pipelined.layer_1_compressor42_10.A , \multiplier_16x16bit_pipelined.layer_1_compressor42_9.B , \multiplier_16x16bit_pipelined.layer_1_compressor42_8.B , \multiplier_16x16bit_pipelined.layer_1_compressor42_7.B , \multiplier_16x16bit_pipelined.layer_1_compressor42_6.B , \multiplier_16x16bit_pipelined.layer_1_compressor42_5.B , \multiplier_16x16bit_pipelined.layer_1_compressor42_4.B , \multiplier_16x16bit_pipelined.layer_1_compressor42_3.B , \multiplier_16x16bit_pipelined.layer_1_compressor42_2.B , \multiplier_16x16bit_pipelined.layer_1_compressor42_1.B , \multiplier_16x16bit_pipelined.layer_1_full_adder_2.B , \multiplier_16x16bit_pipelined.layer_1_compressor42_0.B , \multiplier_16x16bit_pipelined.layer_1_full_adder_1.B , \multiplier_16x16bit_pipelined.layer_1_full_adder_0.B , \multiplier_16x16bit_pipelined.layer_0_w3[1] , \multiplier_16x16bit_pipelined.layer_0_w2[1] };
  assign \multiplier_16x16bit_pipelined.partial_product_gen_1.zero = \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_1.zero ;
  assign \multiplier_16x16bit_pipelined.partial_product_gen_2.double = \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_2.double ;
  assign \multiplier_16x16bit_pipelined.partial_product_gen_2.md = \multiplier_16x16bit_pipelined.md ;
  assign \multiplier_16x16bit_pipelined.partial_product_gen_2.negation = \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_2.negation ;
  assign \multiplier_16x16bit_pipelined.partial_product_gen_2.pp = { \multiplier_16x16bit_pipelined.layer_1_compressor42_13.A , \multiplier_16x16bit_pipelined.layer_1_compressor42_12.A , \multiplier_16x16bit_pipelined.layer_1_compressor42_11.B , \multiplier_16x16bit_pipelined.layer_1_compressor42_10.B , \multiplier_16x16bit_pipelined.layer_1_compressor42_9.C , \multiplier_16x16bit_pipelined.layer_1_compressor42_8.C , \multiplier_16x16bit_pipelined.layer_1_compressor42_7.C , \multiplier_16x16bit_pipelined.layer_1_compressor42_6.C , \multiplier_16x16bit_pipelined.layer_1_compressor42_5.C , \multiplier_16x16bit_pipelined.layer_1_compressor42_4.C , \multiplier_16x16bit_pipelined.layer_1_compressor42_3.C , \multiplier_16x16bit_pipelined.layer_1_compressor42_2.C , \multiplier_16x16bit_pipelined.layer_1_compressor42_1.C , \multiplier_16x16bit_pipelined.layer_1_full_adder_2.cin , \multiplier_16x16bit_pipelined.layer_1_compressor42_0.C , \multiplier_16x16bit_pipelined.layer_1_full_adder_1.cin , \multiplier_16x16bit_pipelined.layer_1_full_adder_0.cin };
  assign \multiplier_16x16bit_pipelined.partial_product_gen_2.zero = \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_2.zero ;
  assign \multiplier_16x16bit_pipelined.partial_product_gen_3.double = \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_3.double ;
  assign \multiplier_16x16bit_pipelined.partial_product_gen_3.md = \multiplier_16x16bit_pipelined.md ;
  assign \multiplier_16x16bit_pipelined.partial_product_gen_3.negation = \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_3.negation ;
  assign \multiplier_16x16bit_pipelined.partial_product_gen_3.pp = { \multiplier_16x16bit_pipelined.layer_1_compressor42_15.A , \multiplier_16x16bit_pipelined.layer_1_compressor42_14.A , \multiplier_16x16bit_pipelined.layer_1_compressor42_13.B , \multiplier_16x16bit_pipelined.layer_1_compressor42_12.B , \multiplier_16x16bit_pipelined.layer_1_compressor42_11.C , \multiplier_16x16bit_pipelined.layer_1_compressor42_10.C , \multiplier_16x16bit_pipelined.layer_1_compressor42_9.D , \multiplier_16x16bit_pipelined.layer_1_compressor42_8.D , \multiplier_16x16bit_pipelined.layer_1_compressor42_7.D , \multiplier_16x16bit_pipelined.layer_1_compressor42_6.D , \multiplier_16x16bit_pipelined.layer_1_compressor42_5.D , \multiplier_16x16bit_pipelined.layer_1_compressor42_4.D , \multiplier_16x16bit_pipelined.layer_1_compressor42_3.D , \multiplier_16x16bit_pipelined.layer_1_compressor42_2.D , \multiplier_16x16bit_pipelined.layer_1_compressor42_1.D , \multiplier_16x16bit_pipelined.layer_0_w7[3] , \multiplier_16x16bit_pipelined.layer_1_compressor42_0.D };
  assign \multiplier_16x16bit_pipelined.partial_product_gen_3.zero = \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_3.zero ;
  assign \multiplier_16x16bit_pipelined.partial_product_gen_4.double = \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_4.double ;
  assign \multiplier_16x16bit_pipelined.partial_product_gen_4.md = \multiplier_16x16bit_pipelined.md ;
  assign \multiplier_16x16bit_pipelined.partial_product_gen_4.negation = \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_4.negation ;
  assign \multiplier_16x16bit_pipelined.partial_product_gen_4.pp = { \multiplier_16x16bit_pipelined.layer_1_full_adder_8.A , \multiplier_16x16bit_pipelined.layer_1_compressor42_16.A , \multiplier_16x16bit_pipelined.layer_1_compressor42_15.B , \multiplier_16x16bit_pipelined.layer_1_compressor42_14.B , \multiplier_16x16bit_pipelined.layer_1_compressor42_13.C , \multiplier_16x16bit_pipelined.layer_1_compressor42_12.C , \multiplier_16x16bit_pipelined.layer_1_compressor42_11.D , \multiplier_16x16bit_pipelined.layer_1_compressor42_10.D , \multiplier_16x16bit_pipelined.layer_1_compressor42_9.cin , \multiplier_16x16bit_pipelined.layer_1_compressor42_8.cin , \multiplier_16x16bit_pipelined.layer_1_compressor42_7.cin , \multiplier_16x16bit_pipelined.layer_1_compressor42_6.cin , \multiplier_16x16bit_pipelined.layer_1_compressor42_5.cin , \multiplier_16x16bit_pipelined.layer_1_compressor42_4.cin , \multiplier_16x16bit_pipelined.layer_1_compressor42_3.cin , \multiplier_16x16bit_pipelined.layer_1_compressor42_2.cin , \multiplier_16x16bit_pipelined.layer_1_compressor42_1.cin };
  assign \multiplier_16x16bit_pipelined.partial_product_gen_4.zero = \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_4.zero ;
  assign \multiplier_16x16bit_pipelined.partial_product_gen_5.double = \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_5.double ;
  assign \multiplier_16x16bit_pipelined.partial_product_gen_5.md = \multiplier_16x16bit_pipelined.md ;
  assign \multiplier_16x16bit_pipelined.partial_product_gen_5.negation = \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_5.negation ;
  assign \multiplier_16x16bit_pipelined.partial_product_gen_5.pp = { \multiplier_16x16bit_pipelined.layer_1_full_adder_10.A , \multiplier_16x16bit_pipelined.layer_1_full_adder_9.A , \multiplier_16x16bit_pipelined.layer_1_full_adder_8.B , \multiplier_16x16bit_pipelined.layer_1_compressor42_16.B , \multiplier_16x16bit_pipelined.layer_1_compressor42_15.C , \multiplier_16x16bit_pipelined.layer_1_compressor42_14.C , \multiplier_16x16bit_pipelined.layer_1_compressor42_13.D , \multiplier_16x16bit_pipelined.layer_1_compressor42_12.D , \multiplier_16x16bit_pipelined.layer_1_compressor42_11.cin , \multiplier_16x16bit_pipelined.layer_1_compressor42_10.cin , \multiplier_16x16bit_pipelined.layer_1_full_adder_6.A , \multiplier_16x16bit_pipelined.layer_1_full_adder_5.A , \multiplier_16x16bit_pipelined.layer_1_full_adder_4.A , \multiplier_16x16bit_pipelined.layer_2_compressor42_1.cin , \multiplier_16x16bit_pipelined.layer_1_full_adder_3.A , \multiplier_16x16bit_pipelined.layer_0_w11[5] , \multiplier_16x16bit_pipelined.layer_2_compressor42_0.D };
  assign \multiplier_16x16bit_pipelined.partial_product_gen_5.zero = \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_5.zero ;
  assign \multiplier_16x16bit_pipelined.partial_product_gen_6.double = \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_6.double ;
  assign \multiplier_16x16bit_pipelined.partial_product_gen_6.md = \multiplier_16x16bit_pipelined.md ;
  assign \multiplier_16x16bit_pipelined.partial_product_gen_6.negation = \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_6.negation ;
  assign \multiplier_16x16bit_pipelined.partial_product_gen_6.pp = { \multiplier_16x16bit_pipelined.layer_2_full_adder_11.B , \multiplier_16x16bit_pipelined.layer_1_full_adder_11.A , \multiplier_16x16bit_pipelined.layer_1_full_adder_10.B , \multiplier_16x16bit_pipelined.layer_1_full_adder_9.B , \multiplier_16x16bit_pipelined.layer_1_full_adder_8.cin , \multiplier_16x16bit_pipelined.layer_1_compressor42_16.C , \multiplier_16x16bit_pipelined.layer_1_compressor42_15.D , \multiplier_16x16bit_pipelined.layer_1_compressor42_14.D , \multiplier_16x16bit_pipelined.layer_1_compressor42_13.cin , \multiplier_16x16bit_pipelined.layer_1_compressor42_12.cin , \multiplier_16x16bit_pipelined.layer_2_compressor42_6.cin , \multiplier_16x16bit_pipelined.layer_1_full_adder_7.A , \multiplier_16x16bit_pipelined.layer_1_full_adder_6.B , \multiplier_16x16bit_pipelined.layer_1_full_adder_5.B , \multiplier_16x16bit_pipelined.layer_1_full_adder_4.B , \multiplier_16x16bit_pipelined.layer_0_w13[6] , \multiplier_16x16bit_pipelined.layer_1_full_adder_3.B };
  assign \multiplier_16x16bit_pipelined.partial_product_gen_6.zero = \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_6.zero ;
  assign \multiplier_16x16bit_pipelined.partial_product_gen_7.double = \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_7.double ;
  assign \multiplier_16x16bit_pipelined.partial_product_gen_7.md = \multiplier_16x16bit_pipelined.md ;
  assign \multiplier_16x16bit_pipelined.partial_product_gen_7.negation = \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_7.negation ;
  assign \multiplier_16x16bit_pipelined.partial_product_gen_7.pp = { \multiplier_16x16bit_pipelined.layer_0_w30 , \multiplier_16x16bit_pipelined.layer_0_w29[0] , \multiplier_16x16bit_pipelined.layer_2_full_adder_11.cin , \multiplier_16x16bit_pipelined.layer_1_full_adder_11.B , \multiplier_16x16bit_pipelined.layer_1_full_adder_10.cin , \multiplier_16x16bit_pipelined.layer_1_full_adder_9.cin , \multiplier_16x16bit_pipelined.layer_0_w24[3] , \multiplier_16x16bit_pipelined.layer_1_compressor42_16.D , \multiplier_16x16bit_pipelined.layer_1_compressor42_15.cin , \multiplier_16x16bit_pipelined.layer_1_compressor42_14.cin , \multiplier_16x16bit_pipelined.layer_0_w20[5] , \multiplier_16x16bit_pipelined.layer_2_compressor42_7.D , \multiplier_16x16bit_pipelined.layer_0_w18[6] , \multiplier_16x16bit_pipelined.layer_1_full_adder_7.B , \multiplier_16x16bit_pipelined.layer_1_full_adder_6.cin , \multiplier_16x16bit_pipelined.layer_1_full_adder_5.cin , \multiplier_16x16bit_pipelined.layer_1_full_adder_4.cin };
  assign \multiplier_16x16bit_pipelined.partial_product_gen_7.zero = \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_7.zero ;
  assign \multiplier_16x16bit_pipelined.zero = { \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_7.zero , \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_6.zero , \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_5.zero , \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_4.zero , \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_3.zero , \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_2.zero , \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_1.zero , \multiplier_16x16bit_pipelined.booth_array_0.booth_radix4_0.zero };
  assign o_un = un;
  assign product = { \multiplier_16x16bit_pipelined.adder_32bit.o_s [31:1], \multiplier_16x16bit_pipelined.adder_32bit.operator_A_0.P };
  assign \rdata[0] = { kp[15], kp[15], kp[15], kp[15], kp[15], kp[15], kp[15], kp[15], kp[15], kp[15], kp[15], kp[15], kp[15], kp[15], kp[15], kp[15], kp };
  assign \rdata[10] = { 27'b000000000000000000000000000, of };
  assign \rdata[1] = { ki[15], ki[15], ki[15], ki[15], ki[15], ki[15], ki[15], ki[15], ki[15], ki[15], ki[15], ki[15], ki[15], ki[15], ki[15], ki[15], ki };
  assign \rdata[2] = { kd[15], kd[15], kd[15], kd[15], kd[15], kd[15], kd[15], kd[15], kd[15], kd[15], kd[15], kd[15], kd[15], kd[15], kd[15], kd[15], kd };
  assign \rdata[3] = { sp[15], sp[15], sp[15], sp[15], sp[15], sp[15], sp[15], sp[15], sp[15], sp[15], sp[15], sp[15], sp[15], sp[15], sp[15], sp[15], sp };
  assign \rdata[4] = { pv[15], pv[15], pv[15], pv[15], pv[15], pv[15], pv[15], pv[15], pv[15], pv[15], pv[15], pv[15], pv[15], pv[15], pv[15], pv[15], pv };
  assign \rdata[5] = { kpd[15], kpd[15], kpd[15], kpd[15], kpd[15], kpd[15], kpd[15], kpd[15], kpd[15], kpd[15], kpd[15], kpd[15], kpd[15], kpd[15], kpd[15], kpd[15], kpd };
  assign \rdata[6] = { \err[0] [15], \err[0] [15], \err[0] [15], \err[0] [15], \err[0] [15], \err[0] [15], \err[0] [15], \err[0] [15], \err[0] [15], \err[0] [15], \err[0] [15], \err[0] [15], \err[0] [15], \err[0] [15], \err[0] [15], \err[0] [15], \err[0] };
  assign \rdata[7] = { \err[1] [15], \err[1] [15], \err[1] [15], \err[1] [15], \err[1] [15], \err[1] [15], \err[1] [15], \err[1] [15], \err[1] [15], \err[1] [15], \err[1] [15], \err[1] [15], \err[1] [15], \err[1] [15], \err[1] [15], \err[1] [15], \err[1] };
  assign \rdata[8] = un;
  assign \rdata[9] = sigma;
  assign rl[10:6] = { rla, rlb, rlb, rlb, rlb };
  assign rl[4:0] = { 5'b00000 };
  assign sum = \adder_32bit_0.o_s ;
  assign wl = { wla, wla, wla, wlb, wlb, 3'b000 };
endmodule
