module NV_NVDLA_CDMA_IMG_sg2pack_fifo_flopram_rwsa_128x11(clk, clk_mgated, pwrbus_ram_pd, di, iwe, we, wa, ra, dout);
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:422" *)
  wire [10:0] _0000_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:577" *)
  wire [10:0] _0001_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:577" *)
  wire [10:0] _0002_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:577" *)
  wire [10:0] _0003_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:577" *)
  wire [10:0] _0004_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:577" *)
  wire [10:0] _0005_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:577" *)
  wire [10:0] _0006_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:577" *)
  wire [10:0] _0007_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:577" *)
  wire [10:0] _0008_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:577" *)
  wire [10:0] _0009_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:577" *)
  wire [10:0] _0010_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:577" *)
  wire [10:0] _0011_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:577" *)
  wire [10:0] _0012_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:577" *)
  wire [10:0] _0013_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:577" *)
  wire [10:0] _0014_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:577" *)
  wire [10:0] _0015_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:577" *)
  wire [10:0] _0016_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:577" *)
  wire [10:0] _0017_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:577" *)
  wire [10:0] _0018_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:577" *)
  wire [10:0] _0019_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:577" *)
  wire [10:0] _0020_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:577" *)
  wire [10:0] _0021_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:577" *)
  wire [10:0] _0022_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:577" *)
  wire [10:0] _0023_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:577" *)
  wire [10:0] _0024_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:577" *)
  wire [10:0] _0025_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:577" *)
  wire [10:0] _0026_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:577" *)
  wire [10:0] _0027_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:577" *)
  wire [10:0] _0028_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:577" *)
  wire [10:0] _0029_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:577" *)
  wire [10:0] _0030_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:577" *)
  wire [10:0] _0031_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:577" *)
  wire [10:0] _0032_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:577" *)
  wire [10:0] _0033_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:577" *)
  wire [10:0] _0034_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:577" *)
  wire [10:0] _0035_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:577" *)
  wire [10:0] _0036_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:577" *)
  wire [10:0] _0037_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:577" *)
  wire [10:0] _0038_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:577" *)
  wire [10:0] _0039_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:577" *)
  wire [10:0] _0040_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:577" *)
  wire [10:0] _0041_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:577" *)
  wire [10:0] _0042_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:577" *)
  wire [10:0] _0043_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:577" *)
  wire [10:0] _0044_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:577" *)
  wire [10:0] _0045_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:577" *)
  wire [10:0] _0046_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:577" *)
  wire [10:0] _0047_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:577" *)
  wire [10:0] _0048_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:577" *)
  wire [10:0] _0049_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:577" *)
  wire [10:0] _0050_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:577" *)
  wire [10:0] _0051_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:577" *)
  wire [10:0] _0052_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:577" *)
  wire [10:0] _0053_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:577" *)
  wire [10:0] _0054_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:577" *)
  wire [10:0] _0055_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:577" *)
  wire [10:0] _0056_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:577" *)
  wire [10:0] _0057_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:577" *)
  wire [10:0] _0058_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:577" *)
  wire [10:0] _0059_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:577" *)
  wire [10:0] _0060_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:577" *)
  wire [10:0] _0061_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:577" *)
  wire [10:0] _0062_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:577" *)
  wire [10:0] _0063_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:577" *)
  wire [10:0] _0064_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:577" *)
  wire [10:0] _0065_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:577" *)
  wire [10:0] _0066_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:577" *)
  wire [10:0] _0067_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:577" *)
  wire [10:0] _0068_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:577" *)
  wire [10:0] _0069_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:577" *)
  wire [10:0] _0070_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:577" *)
  wire [10:0] _0071_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:577" *)
  wire [10:0] _0072_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:577" *)
  wire [10:0] _0073_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:577" *)
  wire [10:0] _0074_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:577" *)
  wire [10:0] _0075_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:577" *)
  wire [10:0] _0076_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:577" *)
  wire [10:0] _0077_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:577" *)
  wire [10:0] _0078_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:577" *)
  wire [10:0] _0079_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:577" *)
  wire [10:0] _0080_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:577" *)
  wire [10:0] _0081_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:577" *)
  wire [10:0] _0082_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:577" *)
  wire [10:0] _0083_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:577" *)
  wire [10:0] _0084_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:577" *)
  wire [10:0] _0085_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:577" *)
  wire [10:0] _0086_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:577" *)
  wire [10:0] _0087_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:577" *)
  wire [10:0] _0088_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:577" *)
  wire [10:0] _0089_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:577" *)
  wire [10:0] _0090_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:577" *)
  wire [10:0] _0091_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:577" *)
  wire [10:0] _0092_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:577" *)
  wire [10:0] _0093_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:577" *)
  wire [10:0] _0094_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:577" *)
  wire [10:0] _0095_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:577" *)
  wire [10:0] _0096_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:577" *)
  wire [10:0] _0097_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:577" *)
  wire [10:0] _0098_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:577" *)
  wire [10:0] _0099_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:577" *)
  wire [10:0] _0100_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:577" *)
  wire [10:0] _0101_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:577" *)
  wire [10:0] _0102_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:577" *)
  wire [10:0] _0103_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:577" *)
  wire [10:0] _0104_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:577" *)
  wire [10:0] _0105_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:577" *)
  wire [10:0] _0106_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:577" *)
  wire [10:0] _0107_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:577" *)
  wire [10:0] _0108_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:577" *)
  wire [10:0] _0109_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:577" *)
  wire [10:0] _0110_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:577" *)
  wire [10:0] _0111_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:577" *)
  wire [10:0] _0112_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:577" *)
  wire [10:0] _0113_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:577" *)
  wire [10:0] _0114_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:577" *)
  wire [10:0] _0115_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:577" *)
  wire [10:0] _0116_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:577" *)
  wire [10:0] _0117_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:577" *)
  wire [10:0] _0118_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:577" *)
  wire [10:0] _0119_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:577" *)
  wire [10:0] _0120_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:577" *)
  wire [10:0] _0121_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:577" *)
  wire [10:0] _0122_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:577" *)
  wire [10:0] _0123_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:577" *)
  wire [10:0] _0124_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:577" *)
  wire [10:0] _0125_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:577" *)
  wire [10:0] _0126_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:577" *)
  wire [10:0] _0127_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:577" *)
  wire [10:0] _0128_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:578" *)
  wire _0129_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:581" *)
  wire _0130_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:584" *)
  wire _0131_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:587" *)
  wire _0132_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:590" *)
  wire _0133_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:593" *)
  wire _0134_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:596" *)
  wire _0135_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:599" *)
  wire _0136_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:602" *)
  wire _0137_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:605" *)
  wire _0138_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:608" *)
  wire _0139_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:611" *)
  wire _0140_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:614" *)
  wire _0141_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:617" *)
  wire _0142_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:620" *)
  wire _0143_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:623" *)
  wire _0144_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:626" *)
  wire _0145_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:629" *)
  wire _0146_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:632" *)
  wire _0147_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:635" *)
  wire _0148_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:638" *)
  wire _0149_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:641" *)
  wire _0150_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:644" *)
  wire _0151_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:647" *)
  wire _0152_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:650" *)
  wire _0153_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:653" *)
  wire _0154_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:656" *)
  wire _0155_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:659" *)
  wire _0156_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:662" *)
  wire _0157_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:665" *)
  wire _0158_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:668" *)
  wire _0159_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:671" *)
  wire _0160_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:674" *)
  wire _0161_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:677" *)
  wire _0162_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:680" *)
  wire _0163_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:683" *)
  wire _0164_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:686" *)
  wire _0165_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:689" *)
  wire _0166_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:692" *)
  wire _0167_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:695" *)
  wire _0168_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:698" *)
  wire _0169_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:701" *)
  wire _0170_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:704" *)
  wire _0171_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:707" *)
  wire _0172_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:710" *)
  wire _0173_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:713" *)
  wire _0174_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:716" *)
  wire _0175_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:719" *)
  wire _0176_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:722" *)
  wire _0177_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:725" *)
  wire _0178_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:728" *)
  wire _0179_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:731" *)
  wire _0180_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:734" *)
  wire _0181_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:737" *)
  wire _0182_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:740" *)
  wire _0183_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:743" *)
  wire _0184_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:746" *)
  wire _0185_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:749" *)
  wire _0186_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:752" *)
  wire _0187_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:755" *)
  wire _0188_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:758" *)
  wire _0189_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:761" *)
  wire _0190_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:764" *)
  wire _0191_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:767" *)
  wire _0192_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:770" *)
  wire _0193_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:773" *)
  wire _0194_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:776" *)
  wire _0195_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:779" *)
  wire _0196_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:782" *)
  wire _0197_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:785" *)
  wire _0198_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:788" *)
  wire _0199_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:791" *)
  wire _0200_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:794" *)
  wire _0201_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:797" *)
  wire _0202_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:800" *)
  wire _0203_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:803" *)
  wire _0204_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:806" *)
  wire _0205_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:809" *)
  wire _0206_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:812" *)
  wire _0207_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:815" *)
  wire _0208_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:818" *)
  wire _0209_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:821" *)
  wire _0210_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:824" *)
  wire _0211_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:827" *)
  wire _0212_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:830" *)
  wire _0213_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:833" *)
  wire _0214_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:836" *)
  wire _0215_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:839" *)
  wire _0216_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:842" *)
  wire _0217_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:845" *)
  wire _0218_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:848" *)
  wire _0219_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:851" *)
  wire _0220_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:854" *)
  wire _0221_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:857" *)
  wire _0222_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:860" *)
  wire _0223_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:863" *)
  wire _0224_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:866" *)
  wire _0225_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:869" *)
  wire _0226_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:872" *)
  wire _0227_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:875" *)
  wire _0228_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:878" *)
  wire _0229_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:881" *)
  wire _0230_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:884" *)
  wire _0231_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:887" *)
  wire _0232_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:890" *)
  wire _0233_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:893" *)
  wire _0234_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:896" *)
  wire _0235_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:899" *)
  wire _0236_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:902" *)
  wire _0237_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:905" *)
  wire _0238_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:908" *)
  wire _0239_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:911" *)
  wire _0240_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:914" *)
  wire _0241_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:917" *)
  wire _0242_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:920" *)
  wire _0243_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:923" *)
  wire _0244_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:926" *)
  wire _0245_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:929" *)
  wire _0246_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:932" *)
  wire _0247_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:935" *)
  wire _0248_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:938" *)
  wire _0249_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:941" *)
  wire _0250_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:944" *)
  wire _0251_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:947" *)
  wire _0252_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:950" *)
  wire _0253_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:953" *)
  wire _0254_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:956" *)
  wire _0255_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:959" *)
  wire _0256_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:578" *)
  wire _0257_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:581" *)
  wire _0258_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:584" *)
  wire _0259_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:587" *)
  wire _0260_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:590" *)
  wire _0261_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:593" *)
  wire _0262_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:596" *)
  wire _0263_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:599" *)
  wire _0264_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:602" *)
  wire _0265_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:605" *)
  wire _0266_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:608" *)
  wire _0267_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:611" *)
  wire _0268_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:614" *)
  wire _0269_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:617" *)
  wire _0270_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:620" *)
  wire _0271_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:623" *)
  wire _0272_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:626" *)
  wire _0273_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:629" *)
  wire _0274_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:632" *)
  wire _0275_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:635" *)
  wire _0276_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:638" *)
  wire _0277_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:641" *)
  wire _0278_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:644" *)
  wire _0279_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:647" *)
  wire _0280_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:650" *)
  wire _0281_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:653" *)
  wire _0282_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:656" *)
  wire _0283_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:659" *)
  wire _0284_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:662" *)
  wire _0285_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:665" *)
  wire _0286_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:668" *)
  wire _0287_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:671" *)
  wire _0288_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:674" *)
  wire _0289_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:677" *)
  wire _0290_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:680" *)
  wire _0291_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:683" *)
  wire _0292_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:686" *)
  wire _0293_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:689" *)
  wire _0294_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:692" *)
  wire _0295_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:695" *)
  wire _0296_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:698" *)
  wire _0297_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:701" *)
  wire _0298_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:704" *)
  wire _0299_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:707" *)
  wire _0300_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:710" *)
  wire _0301_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:713" *)
  wire _0302_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:716" *)
  wire _0303_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:719" *)
  wire _0304_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:722" *)
  wire _0305_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:725" *)
  wire _0306_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:728" *)
  wire _0307_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:731" *)
  wire _0308_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:734" *)
  wire _0309_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:737" *)
  wire _0310_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:740" *)
  wire _0311_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:743" *)
  wire _0312_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:746" *)
  wire _0313_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:749" *)
  wire _0314_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:752" *)
  wire _0315_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:755" *)
  wire _0316_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:758" *)
  wire _0317_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:761" *)
  wire _0318_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:764" *)
  wire _0319_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:767" *)
  wire _0320_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:770" *)
  wire _0321_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:773" *)
  wire _0322_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:776" *)
  wire _0323_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:779" *)
  wire _0324_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:782" *)
  wire _0325_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:785" *)
  wire _0326_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:788" *)
  wire _0327_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:791" *)
  wire _0328_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:794" *)
  wire _0329_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:797" *)
  wire _0330_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:800" *)
  wire _0331_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:803" *)
  wire _0332_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:806" *)
  wire _0333_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:809" *)
  wire _0334_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:812" *)
  wire _0335_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:815" *)
  wire _0336_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:818" *)
  wire _0337_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:821" *)
  wire _0338_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:824" *)
  wire _0339_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:827" *)
  wire _0340_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:830" *)
  wire _0341_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:833" *)
  wire _0342_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:836" *)
  wire _0343_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:839" *)
  wire _0344_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:842" *)
  wire _0345_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:845" *)
  wire _0346_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:848" *)
  wire _0347_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:851" *)
  wire _0348_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:854" *)
  wire _0349_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:857" *)
  wire _0350_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:860" *)
  wire _0351_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:863" *)
  wire _0352_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:866" *)
  wire _0353_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:869" *)
  wire _0354_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:872" *)
  wire _0355_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:875" *)
  wire _0356_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:878" *)
  wire _0357_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:881" *)
  wire _0358_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:884" *)
  wire _0359_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:887" *)
  wire _0360_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:890" *)
  wire _0361_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:893" *)
  wire _0362_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:896" *)
  wire _0363_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:899" *)
  wire _0364_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:902" *)
  wire _0365_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:905" *)
  wire _0366_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:908" *)
  wire _0367_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:911" *)
  wire _0368_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:914" *)
  wire _0369_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:917" *)
  wire _0370_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:920" *)
  wire _0371_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:923" *)
  wire _0372_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:926" *)
  wire _0373_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:929" *)
  wire _0374_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:932" *)
  wire _0375_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:935" *)
  wire _0376_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:938" *)
  wire _0377_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:941" *)
  wire _0378_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:944" *)
  wire _0379_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:947" *)
  wire _0380_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:950" *)
  wire _0381_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:953" *)
  wire _0382_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:956" *)
  wire _0383_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:959" *)
  wire _0384_;
  wire _0385_;
  wire _0386_;
  wire _0387_;
  wire _0388_;
  wire _0389_;
  wire _0390_;
  wire _0391_;
  wire _0392_;
  wire _0393_;
  wire _0394_;
  wire _0395_;
  wire _0396_;
  wire _0397_;
  wire _0398_;
  wire _0399_;
  wire _0400_;
  wire _0401_;
  wire _0402_;
  wire _0403_;
  wire _0404_;
  wire _0405_;
  wire _0406_;
  wire _0407_;
  wire _0408_;
  wire _0409_;
  wire _0410_;
  wire _0411_;
  wire _0412_;
  wire _0413_;
  wire _0414_;
  wire _0415_;
  wire _0416_;
  wire _0417_;
  wire _0418_;
  wire _0419_;
  wire _0420_;
  wire _0421_;
  wire _0422_;
  wire _0423_;
  wire _0424_;
  wire _0425_;
  wire _0426_;
  wire _0427_;
  wire _0428_;
  wire _0429_;
  wire _0430_;
  wire _0431_;
  wire _0432_;
  wire _0433_;
  wire _0434_;
  wire _0435_;
  wire _0436_;
  wire _0437_;
  wire _0438_;
  wire _0439_;
  wire _0440_;
  wire _0441_;
  wire _0442_;
  wire _0443_;
  wire _0444_;
  wire _0445_;
  wire _0446_;
  wire _0447_;
  wire _0448_;
  wire _0449_;
  wire _0450_;
  wire _0451_;
  wire _0452_;
  wire _0453_;
  wire _0454_;
  wire _0455_;
  wire _0456_;
  wire _0457_;
  wire _0458_;
  wire _0459_;
  wire _0460_;
  wire _0461_;
  wire _0462_;
  wire _0463_;
  wire _0464_;
  wire _0465_;
  wire _0466_;
  wire _0467_;
  wire _0468_;
  wire _0469_;
  wire _0470_;
  wire _0471_;
  wire _0472_;
  wire _0473_;
  wire _0474_;
  wire _0475_;
  wire _0476_;
  wire _0477_;
  wire _0478_;
  wire _0479_;
  wire _0480_;
  wire _0481_;
  wire _0482_;
  wire _0483_;
  wire _0484_;
  wire _0485_;
  wire _0486_;
  wire _0487_;
  wire _0488_;
  wire _0489_;
  wire _0490_;
  wire _0491_;
  wire _0492_;
  wire _0493_;
  wire _0494_;
  wire _0495_;
  wire _0496_;
  wire _0497_;
  wire _0498_;
  wire _0499_;
  wire _0500_;
  wire _0501_;
  wire _0502_;
  wire _0503_;
  wire _0504_;
  wire _0505_;
  wire _0506_;
  wire _0507_;
  wire _0508_;
  wire _0509_;
  wire _0510_;
  wire _0511_;
  wire _0512_;
  wire _0513_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:380" *)
  input clk;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:381" *)
  input clk_mgated;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:383" *)
  input [10:0] di;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:421" *)
  reg [10:0] di_d;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:388" *)
  output [10:0] dout;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:384" *)
  input iwe;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:382" *)
  input [31:0] pwrbus_ram_pd;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:387" *)
  input [7:0] ra;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:449" *)
  reg [10:0] ram_ff0;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:450" *)
  reg [10:0] ram_ff1;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:459" *)
  reg [10:0] ram_ff10;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:549" *)
  reg [10:0] ram_ff100;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:550" *)
  reg [10:0] ram_ff101;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:551" *)
  reg [10:0] ram_ff102;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:552" *)
  reg [10:0] ram_ff103;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:553" *)
  reg [10:0] ram_ff104;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:554" *)
  reg [10:0] ram_ff105;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:555" *)
  reg [10:0] ram_ff106;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:556" *)
  reg [10:0] ram_ff107;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:557" *)
  reg [10:0] ram_ff108;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:558" *)
  reg [10:0] ram_ff109;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:460" *)
  reg [10:0] ram_ff11;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:559" *)
  reg [10:0] ram_ff110;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:560" *)
  reg [10:0] ram_ff111;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:561" *)
  reg [10:0] ram_ff112;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:562" *)
  reg [10:0] ram_ff113;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:563" *)
  reg [10:0] ram_ff114;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:564" *)
  reg [10:0] ram_ff115;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:565" *)
  reg [10:0] ram_ff116;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:566" *)
  reg [10:0] ram_ff117;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:567" *)
  reg [10:0] ram_ff118;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:568" *)
  reg [10:0] ram_ff119;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:461" *)
  reg [10:0] ram_ff12;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:569" *)
  reg [10:0] ram_ff120;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:570" *)
  reg [10:0] ram_ff121;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:571" *)
  reg [10:0] ram_ff122;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:572" *)
  reg [10:0] ram_ff123;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:573" *)
  reg [10:0] ram_ff124;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:574" *)
  reg [10:0] ram_ff125;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:575" *)
  reg [10:0] ram_ff126;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:576" *)
  reg [10:0] ram_ff127;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:462" *)
  reg [10:0] ram_ff13;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:463" *)
  reg [10:0] ram_ff14;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:464" *)
  reg [10:0] ram_ff15;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:465" *)
  reg [10:0] ram_ff16;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:466" *)
  reg [10:0] ram_ff17;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:467" *)
  reg [10:0] ram_ff18;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:468" *)
  reg [10:0] ram_ff19;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:451" *)
  reg [10:0] ram_ff2;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:469" *)
  reg [10:0] ram_ff20;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:470" *)
  reg [10:0] ram_ff21;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:471" *)
  reg [10:0] ram_ff22;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:472" *)
  reg [10:0] ram_ff23;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:473" *)
  reg [10:0] ram_ff24;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:474" *)
  reg [10:0] ram_ff25;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:475" *)
  reg [10:0] ram_ff26;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:476" *)
  reg [10:0] ram_ff27;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:477" *)
  reg [10:0] ram_ff28;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:478" *)
  reg [10:0] ram_ff29;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:452" *)
  reg [10:0] ram_ff3;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:479" *)
  reg [10:0] ram_ff30;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:480" *)
  reg [10:0] ram_ff31;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:481" *)
  reg [10:0] ram_ff32;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:482" *)
  reg [10:0] ram_ff33;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:483" *)
  reg [10:0] ram_ff34;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:484" *)
  reg [10:0] ram_ff35;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:485" *)
  reg [10:0] ram_ff36;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:486" *)
  reg [10:0] ram_ff37;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:487" *)
  reg [10:0] ram_ff38;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:488" *)
  reg [10:0] ram_ff39;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:453" *)
  reg [10:0] ram_ff4;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:489" *)
  reg [10:0] ram_ff40;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:490" *)
  reg [10:0] ram_ff41;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:491" *)
  reg [10:0] ram_ff42;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:492" *)
  reg [10:0] ram_ff43;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:493" *)
  reg [10:0] ram_ff44;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:494" *)
  reg [10:0] ram_ff45;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:495" *)
  reg [10:0] ram_ff46;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:496" *)
  reg [10:0] ram_ff47;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:497" *)
  reg [10:0] ram_ff48;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:498" *)
  reg [10:0] ram_ff49;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:454" *)
  reg [10:0] ram_ff5;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:499" *)
  reg [10:0] ram_ff50;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:500" *)
  reg [10:0] ram_ff51;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:501" *)
  reg [10:0] ram_ff52;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:502" *)
  reg [10:0] ram_ff53;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:503" *)
  reg [10:0] ram_ff54;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:504" *)
  reg [10:0] ram_ff55;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:505" *)
  reg [10:0] ram_ff56;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:506" *)
  reg [10:0] ram_ff57;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:507" *)
  reg [10:0] ram_ff58;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:508" *)
  reg [10:0] ram_ff59;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:455" *)
  reg [10:0] ram_ff6;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:509" *)
  reg [10:0] ram_ff60;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:510" *)
  reg [10:0] ram_ff61;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:511" *)
  reg [10:0] ram_ff62;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:512" *)
  reg [10:0] ram_ff63;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:513" *)
  reg [10:0] ram_ff64;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:514" *)
  reg [10:0] ram_ff65;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:515" *)
  reg [10:0] ram_ff66;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:516" *)
  reg [10:0] ram_ff67;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:517" *)
  reg [10:0] ram_ff68;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:518" *)
  reg [10:0] ram_ff69;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:456" *)
  reg [10:0] ram_ff7;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:519" *)
  reg [10:0] ram_ff70;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:520" *)
  reg [10:0] ram_ff71;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:521" *)
  reg [10:0] ram_ff72;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:522" *)
  reg [10:0] ram_ff73;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:523" *)
  reg [10:0] ram_ff74;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:524" *)
  reg [10:0] ram_ff75;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:525" *)
  reg [10:0] ram_ff76;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:526" *)
  reg [10:0] ram_ff77;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:527" *)
  reg [10:0] ram_ff78;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:528" *)
  reg [10:0] ram_ff79;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:457" *)
  reg [10:0] ram_ff8;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:529" *)
  reg [10:0] ram_ff80;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:530" *)
  reg [10:0] ram_ff81;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:531" *)
  reg [10:0] ram_ff82;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:532" *)
  reg [10:0] ram_ff83;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:533" *)
  reg [10:0] ram_ff84;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:534" *)
  reg [10:0] ram_ff85;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:535" *)
  reg [10:0] ram_ff86;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:536" *)
  reg [10:0] ram_ff87;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:537" *)
  reg [10:0] ram_ff88;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:538" *)
  reg [10:0] ram_ff89;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:458" *)
  reg [10:0] ram_ff9;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:539" *)
  reg [10:0] ram_ff90;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:540" *)
  reg [10:0] ram_ff91;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:541" *)
  reg [10:0] ram_ff92;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:542" *)
  reg [10:0] ram_ff93;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:543" *)
  reg [10:0] ram_ff94;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:544" *)
  reg [10:0] ram_ff95;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:545" *)
  reg [10:0] ram_ff96;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:546" *)
  reg [10:0] ram_ff97;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:547" *)
  reg [10:0] ram_ff98;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:548" *)
  reg [10:0] ram_ff99;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:386" *)
  input [6:0] wa;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:385" *)
  input we;
  assign _0129_ = ! (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:578" *) wa;
  assign _0130_ = wa == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:581" *) 1'b1;
  assign _0131_ = wa == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:584" *) 2'b10;
  assign _0132_ = wa == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:587" *) 2'b11;
  assign _0133_ = wa == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:590" *) 3'b100;
  assign _0134_ = wa == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:593" *) 3'b101;
  assign _0135_ = wa == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:596" *) 3'b110;
  assign _0136_ = wa == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:599" *) 3'b111;
  assign _0137_ = wa == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:602" *) 4'b1000;
  assign _0138_ = wa == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:605" *) 4'b1001;
  assign _0139_ = wa == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:608" *) 4'b1010;
  assign _0140_ = wa == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:611" *) 4'b1011;
  assign _0141_ = wa == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:614" *) 4'b1100;
  assign _0142_ = wa == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:617" *) 4'b1101;
  assign _0143_ = wa == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:620" *) 4'b1110;
  assign _0144_ = wa == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:623" *) 4'b1111;
  assign _0145_ = wa == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:626" *) 5'b10000;
  assign _0146_ = wa == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:629" *) 5'b10001;
  assign _0147_ = wa == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:632" *) 5'b10010;
  assign _0148_ = wa == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:635" *) 5'b10011;
  assign _0149_ = wa == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:638" *) 5'b10100;
  assign _0150_ = wa == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:641" *) 5'b10101;
  assign _0151_ = wa == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:644" *) 5'b10110;
  assign _0152_ = wa == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:647" *) 5'b10111;
  assign _0153_ = wa == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:650" *) 5'b11000;
  assign _0154_ = wa == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:653" *) 5'b11001;
  assign _0155_ = wa == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:656" *) 5'b11010;
  assign _0156_ = wa == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:659" *) 5'b11011;
  assign _0157_ = wa == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:662" *) 5'b11100;
  assign _0158_ = wa == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:665" *) 5'b11101;
  assign _0159_ = wa == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:668" *) 5'b11110;
  assign _0160_ = wa == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:671" *) 5'b11111;
  assign _0161_ = wa == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:674" *) 6'b100000;
  assign _0162_ = wa == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:677" *) 6'b100001;
  assign _0163_ = wa == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:680" *) 6'b100010;
  assign _0164_ = wa == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:683" *) 6'b100011;
  assign _0165_ = wa == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:686" *) 6'b100100;
  assign _0166_ = wa == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:689" *) 6'b100101;
  assign _0167_ = wa == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:692" *) 6'b100110;
  assign _0168_ = wa == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:695" *) 6'b100111;
  assign _0169_ = wa == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:698" *) 6'b101000;
  assign _0170_ = wa == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:701" *) 6'b101001;
  assign _0171_ = wa == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:704" *) 6'b101010;
  assign _0172_ = wa == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:707" *) 6'b101011;
  assign _0173_ = wa == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:710" *) 6'b101100;
  assign _0174_ = wa == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:713" *) 6'b101101;
  assign _0175_ = wa == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:716" *) 6'b101110;
  assign _0176_ = wa == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:719" *) 6'b101111;
  assign _0177_ = wa == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:722" *) 6'b110000;
  assign _0178_ = wa == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:725" *) 6'b110001;
  assign _0179_ = wa == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:728" *) 6'b110010;
  assign _0180_ = wa == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:731" *) 6'b110011;
  assign _0181_ = wa == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:734" *) 6'b110100;
  assign _0182_ = wa == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:737" *) 6'b110101;
  assign _0183_ = wa == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:740" *) 6'b110110;
  assign _0184_ = wa == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:743" *) 6'b110111;
  assign _0185_ = wa == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:746" *) 6'b111000;
  assign _0186_ = wa == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:749" *) 6'b111001;
  assign _0187_ = wa == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:752" *) 6'b111010;
  assign _0188_ = wa == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:755" *) 6'b111011;
  assign _0189_ = wa == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:758" *) 6'b111100;
  assign _0190_ = wa == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:761" *) 6'b111101;
  assign _0191_ = wa == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:764" *) 6'b111110;
  assign _0192_ = wa == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:767" *) 6'b111111;
  assign _0193_ = wa == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:770" *) 7'b1000000;
  assign _0194_ = wa == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:773" *) 7'b1000001;
  assign _0195_ = wa == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:776" *) 7'b1000010;
  assign _0196_ = wa == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:779" *) 7'b1000011;
  assign _0197_ = wa == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:782" *) 7'b1000100;
  assign _0198_ = wa == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:785" *) 7'b1000101;
  assign _0199_ = wa == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:788" *) 7'b1000110;
  assign _0200_ = wa == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:791" *) 7'b1000111;
  assign _0201_ = wa == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:794" *) 7'b1001000;
  assign _0202_ = wa == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:797" *) 7'b1001001;
  assign _0203_ = wa == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:800" *) 7'b1001010;
  assign _0204_ = wa == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:803" *) 7'b1001011;
  assign _0205_ = wa == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:806" *) 7'b1001100;
  assign _0206_ = wa == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:809" *) 7'b1001101;
  assign _0207_ = wa == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:812" *) 7'b1001110;
  assign _0208_ = wa == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:815" *) 7'b1001111;
  assign _0209_ = wa == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:818" *) 7'b1010000;
  assign _0210_ = wa == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:821" *) 7'b1010001;
  assign _0211_ = wa == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:824" *) 7'b1010010;
  assign _0212_ = wa == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:827" *) 7'b1010011;
  assign _0213_ = wa == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:830" *) 7'b1010100;
  assign _0214_ = wa == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:833" *) 7'b1010101;
  assign _0215_ = wa == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:836" *) 7'b1010110;
  assign _0216_ = wa == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:839" *) 7'b1010111;
  assign _0217_ = wa == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:842" *) 7'b1011000;
  assign _0218_ = wa == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:845" *) 7'b1011001;
  assign _0219_ = wa == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:848" *) 7'b1011010;
  assign _0220_ = wa == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:851" *) 7'b1011011;
  assign _0221_ = wa == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:854" *) 7'b1011100;
  assign _0222_ = wa == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:857" *) 7'b1011101;
  assign _0223_ = wa == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:860" *) 7'b1011110;
  assign _0224_ = wa == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:863" *) 7'b1011111;
  assign _0225_ = wa == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:866" *) 7'b1100000;
  assign _0226_ = wa == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:869" *) 7'b1100001;
  assign _0227_ = wa == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:872" *) 7'b1100010;
  assign _0228_ = wa == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:875" *) 7'b1100011;
  assign _0229_ = wa == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:878" *) 7'b1100100;
  assign _0230_ = wa == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:881" *) 7'b1100101;
  assign _0231_ = wa == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:884" *) 7'b1100110;
  assign _0232_ = wa == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:887" *) 7'b1100111;
  assign _0233_ = wa == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:890" *) 7'b1101000;
  assign _0234_ = wa == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:893" *) 7'b1101001;
  assign _0235_ = wa == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:896" *) 7'b1101010;
  assign _0236_ = wa == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:899" *) 7'b1101011;
  assign _0237_ = wa == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:902" *) 7'b1101100;
  assign _0238_ = wa == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:905" *) 7'b1101101;
  assign _0239_ = wa == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:908" *) 7'b1101110;
  assign _0240_ = wa == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:911" *) 7'b1101111;
  assign _0241_ = wa == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:914" *) 7'b1110000;
  assign _0242_ = wa == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:917" *) 7'b1110001;
  assign _0243_ = wa == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:920" *) 7'b1110010;
  assign _0244_ = wa == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:923" *) 7'b1110011;
  assign _0245_ = wa == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:926" *) 7'b1110100;
  assign _0246_ = wa == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:929" *) 7'b1110101;
  assign _0247_ = wa == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:932" *) 7'b1110110;
  assign _0248_ = wa == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:935" *) 7'b1110111;
  assign _0249_ = wa == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:938" *) 7'b1111000;
  assign _0250_ = wa == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:941" *) 7'b1111001;
  assign _0251_ = wa == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:944" *) 7'b1111010;
  assign _0252_ = wa == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:947" *) 7'b1111011;
  assign _0253_ = wa == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:950" *) 7'b1111100;
  assign _0254_ = wa == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:953" *) 7'b1111101;
  assign _0255_ = wa == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:956" *) 7'b1111110;
  assign _0256_ = wa == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:959" *) 7'b1111111;
  assign _0257_ = we && (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:578" *) _0129_;
  assign _0258_ = we && (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:581" *) _0130_;
  assign _0259_ = we && (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:584" *) _0131_;
  assign _0260_ = we && (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:587" *) _0132_;
  assign _0261_ = we && (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:590" *) _0133_;
  assign _0262_ = we && (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:593" *) _0134_;
  assign _0263_ = we && (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:596" *) _0135_;
  assign _0264_ = we && (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:599" *) _0136_;
  assign _0265_ = we && (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:602" *) _0137_;
  assign _0266_ = we && (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:605" *) _0138_;
  assign _0267_ = we && (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:608" *) _0139_;
  assign _0268_ = we && (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:611" *) _0140_;
  assign _0269_ = we && (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:614" *) _0141_;
  assign _0270_ = we && (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:617" *) _0142_;
  assign _0271_ = we && (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:620" *) _0143_;
  assign _0272_ = we && (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:623" *) _0144_;
  assign _0273_ = we && (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:626" *) _0145_;
  assign _0274_ = we && (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:629" *) _0146_;
  assign _0275_ = we && (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:632" *) _0147_;
  assign _0276_ = we && (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:635" *) _0148_;
  assign _0277_ = we && (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:638" *) _0149_;
  assign _0278_ = we && (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:641" *) _0150_;
  assign _0279_ = we && (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:644" *) _0151_;
  assign _0280_ = we && (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:647" *) _0152_;
  assign _0281_ = we && (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:650" *) _0153_;
  assign _0282_ = we && (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:653" *) _0154_;
  assign _0283_ = we && (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:656" *) _0155_;
  assign _0284_ = we && (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:659" *) _0156_;
  assign _0285_ = we && (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:662" *) _0157_;
  assign _0286_ = we && (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:665" *) _0158_;
  assign _0287_ = we && (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:668" *) _0159_;
  assign _0288_ = we && (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:671" *) _0160_;
  assign _0289_ = we && (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:674" *) _0161_;
  assign _0290_ = we && (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:677" *) _0162_;
  assign _0291_ = we && (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:680" *) _0163_;
  assign _0292_ = we && (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:683" *) _0164_;
  assign _0293_ = we && (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:686" *) _0165_;
  assign _0294_ = we && (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:689" *) _0166_;
  assign _0295_ = we && (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:692" *) _0167_;
  assign _0296_ = we && (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:695" *) _0168_;
  assign _0297_ = we && (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:698" *) _0169_;
  assign _0298_ = we && (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:701" *) _0170_;
  assign _0299_ = we && (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:704" *) _0171_;
  assign _0300_ = we && (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:707" *) _0172_;
  assign _0301_ = we && (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:710" *) _0173_;
  assign _0302_ = we && (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:713" *) _0174_;
  assign _0303_ = we && (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:716" *) _0175_;
  assign _0304_ = we && (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:719" *) _0176_;
  assign _0305_ = we && (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:722" *) _0177_;
  assign _0306_ = we && (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:725" *) _0178_;
  assign _0307_ = we && (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:728" *) _0179_;
  assign _0308_ = we && (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:731" *) _0180_;
  assign _0309_ = we && (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:734" *) _0181_;
  assign _0310_ = we && (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:737" *) _0182_;
  assign _0311_ = we && (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:740" *) _0183_;
  assign _0312_ = we && (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:743" *) _0184_;
  assign _0313_ = we && (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:746" *) _0185_;
  assign _0314_ = we && (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:749" *) _0186_;
  assign _0315_ = we && (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:752" *) _0187_;
  assign _0316_ = we && (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:755" *) _0188_;
  assign _0317_ = we && (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:758" *) _0189_;
  assign _0318_ = we && (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:761" *) _0190_;
  assign _0319_ = we && (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:764" *) _0191_;
  assign _0320_ = we && (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:767" *) _0192_;
  assign _0321_ = we && (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:770" *) _0193_;
  assign _0322_ = we && (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:773" *) _0194_;
  assign _0323_ = we && (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:776" *) _0195_;
  assign _0324_ = we && (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:779" *) _0196_;
  assign _0325_ = we && (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:782" *) _0197_;
  assign _0326_ = we && (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:785" *) _0198_;
  assign _0327_ = we && (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:788" *) _0199_;
  assign _0328_ = we && (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:791" *) _0200_;
  assign _0329_ = we && (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:794" *) _0201_;
  assign _0330_ = we && (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:797" *) _0202_;
  assign _0331_ = we && (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:800" *) _0203_;
  assign _0332_ = we && (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:803" *) _0204_;
  assign _0333_ = we && (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:806" *) _0205_;
  assign _0334_ = we && (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:809" *) _0206_;
  assign _0335_ = we && (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:812" *) _0207_;
  assign _0336_ = we && (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:815" *) _0208_;
  assign _0337_ = we && (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:818" *) _0209_;
  assign _0338_ = we && (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:821" *) _0210_;
  assign _0339_ = we && (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:824" *) _0211_;
  assign _0340_ = we && (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:827" *) _0212_;
  assign _0341_ = we && (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:830" *) _0213_;
  assign _0342_ = we && (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:833" *) _0214_;
  assign _0343_ = we && (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:836" *) _0215_;
  assign _0344_ = we && (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:839" *) _0216_;
  assign _0345_ = we && (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:842" *) _0217_;
  assign _0346_ = we && (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:845" *) _0218_;
  assign _0347_ = we && (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:848" *) _0219_;
  assign _0348_ = we && (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:851" *) _0220_;
  assign _0349_ = we && (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:854" *) _0221_;
  assign _0350_ = we && (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:857" *) _0222_;
  assign _0351_ = we && (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:860" *) _0223_;
  assign _0352_ = we && (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:863" *) _0224_;
  assign _0353_ = we && (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:866" *) _0225_;
  assign _0354_ = we && (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:869" *) _0226_;
  assign _0355_ = we && (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:872" *) _0227_;
  assign _0356_ = we && (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:875" *) _0228_;
  assign _0357_ = we && (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:878" *) _0229_;
  assign _0358_ = we && (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:881" *) _0230_;
  assign _0359_ = we && (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:884" *) _0231_;
  assign _0360_ = we && (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:887" *) _0232_;
  assign _0361_ = we && (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:890" *) _0233_;
  assign _0362_ = we && (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:893" *) _0234_;
  assign _0363_ = we && (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:896" *) _0235_;
  assign _0364_ = we && (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:899" *) _0236_;
  assign _0365_ = we && (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:902" *) _0237_;
  assign _0366_ = we && (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:905" *) _0238_;
  assign _0367_ = we && (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:908" *) _0239_;
  assign _0368_ = we && (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:911" *) _0240_;
  assign _0369_ = we && (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:914" *) _0241_;
  assign _0370_ = we && (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:917" *) _0242_;
  assign _0371_ = we && (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:920" *) _0243_;
  assign _0372_ = we && (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:923" *) _0244_;
  assign _0373_ = we && (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:926" *) _0245_;
  assign _0374_ = we && (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:929" *) _0246_;
  assign _0375_ = we && (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:932" *) _0247_;
  assign _0376_ = we && (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:935" *) _0248_;
  assign _0377_ = we && (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:938" *) _0249_;
  assign _0378_ = we && (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:941" *) _0250_;
  assign _0379_ = we && (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:944" *) _0251_;
  assign _0380_ = we && (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:947" *) _0252_;
  assign _0381_ = we && (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:950" *) _0253_;
  assign _0382_ = we && (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:953" *) _0254_;
  assign _0383_ = we && (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:956" *) _0255_;
  assign _0384_ = we && (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:959" *) _0256_;
  always @(posedge clk_mgated)
      ram_ff0 <= _0001_;
  always @(posedge clk_mgated)
      ram_ff1 <= _0040_;
  always @(posedge clk_mgated)
      ram_ff2 <= _0051_;
  always @(posedge clk_mgated)
      ram_ff3 <= _0062_;
  always @(posedge clk_mgated)
      ram_ff4 <= _0073_;
  always @(posedge clk_mgated)
      ram_ff5 <= _0084_;
  always @(posedge clk_mgated)
      ram_ff6 <= _0095_;
  always @(posedge clk_mgated)
      ram_ff7 <= _0106_;
  always @(posedge clk_mgated)
      ram_ff8 <= _0117_;
  always @(posedge clk_mgated)
      ram_ff9 <= _0128_;
  always @(posedge clk_mgated)
      ram_ff10 <= _0012_;
  always @(posedge clk_mgated)
      ram_ff11 <= _0023_;
  always @(posedge clk_mgated)
      ram_ff12 <= _0032_;
  always @(posedge clk_mgated)
      ram_ff13 <= _0033_;
  always @(posedge clk_mgated)
      ram_ff14 <= _0034_;
  always @(posedge clk_mgated)
      ram_ff15 <= _0035_;
  always @(posedge clk_mgated)
      ram_ff16 <= _0036_;
  always @(posedge clk_mgated)
      ram_ff17 <= _0037_;
  always @(posedge clk_mgated)
      ram_ff18 <= _0038_;
  always @(posedge clk_mgated)
      ram_ff19 <= _0039_;
  always @(posedge clk_mgated)
      ram_ff20 <= _0041_;
  always @(posedge clk_mgated)
      ram_ff21 <= _0042_;
  always @(posedge clk_mgated)
      ram_ff22 <= _0043_;
  always @(posedge clk_mgated)
      ram_ff23 <= _0044_;
  always @(posedge clk_mgated)
      ram_ff24 <= _0045_;
  always @(posedge clk_mgated)
      ram_ff25 <= _0046_;
  always @(posedge clk_mgated)
      ram_ff26 <= _0047_;
  always @(posedge clk_mgated)
      ram_ff27 <= _0048_;
  always @(posedge clk_mgated)
      ram_ff28 <= _0049_;
  always @(posedge clk_mgated)
      ram_ff29 <= _0050_;
  always @(posedge clk_mgated)
      ram_ff30 <= _0052_;
  always @(posedge clk_mgated)
      ram_ff31 <= _0053_;
  always @(posedge clk_mgated)
      ram_ff32 <= _0054_;
  always @(posedge clk_mgated)
      ram_ff33 <= _0055_;
  always @(posedge clk_mgated)
      ram_ff34 <= _0056_;
  always @(posedge clk_mgated)
      ram_ff35 <= _0057_;
  always @(posedge clk_mgated)
      ram_ff36 <= _0058_;
  always @(posedge clk_mgated)
      ram_ff37 <= _0059_;
  always @(posedge clk_mgated)
      ram_ff38 <= _0060_;
  always @(posedge clk_mgated)
      ram_ff39 <= _0061_;
  always @(posedge clk_mgated)
      ram_ff40 <= _0063_;
  always @(posedge clk_mgated)
      ram_ff41 <= _0064_;
  always @(posedge clk_mgated)
      ram_ff42 <= _0065_;
  always @(posedge clk_mgated)
      ram_ff43 <= _0066_;
  always @(posedge clk_mgated)
      ram_ff44 <= _0067_;
  always @(posedge clk_mgated)
      ram_ff45 <= _0068_;
  always @(posedge clk_mgated)
      ram_ff46 <= _0069_;
  always @(posedge clk_mgated)
      ram_ff47 <= _0070_;
  always @(posedge clk_mgated)
      ram_ff48 <= _0071_;
  always @(posedge clk_mgated)
      ram_ff49 <= _0072_;
  always @(posedge clk_mgated)
      ram_ff50 <= _0074_;
  always @(posedge clk_mgated)
      ram_ff51 <= _0075_;
  always @(posedge clk_mgated)
      ram_ff52 <= _0076_;
  always @(posedge clk_mgated)
      ram_ff53 <= _0077_;
  always @(posedge clk_mgated)
      ram_ff54 <= _0078_;
  always @(posedge clk_mgated)
      ram_ff55 <= _0079_;
  always @(posedge clk_mgated)
      ram_ff56 <= _0080_;
  always @(posedge clk_mgated)
      ram_ff57 <= _0081_;
  always @(posedge clk_mgated)
      ram_ff58 <= _0082_;
  always @(posedge clk_mgated)
      ram_ff59 <= _0083_;
  always @(posedge clk_mgated)
      ram_ff60 <= _0085_;
  always @(posedge clk_mgated)
      ram_ff61 <= _0086_;
  always @(posedge clk_mgated)
      ram_ff62 <= _0087_;
  always @(posedge clk_mgated)
      ram_ff63 <= _0088_;
  always @(posedge clk_mgated)
      ram_ff64 <= _0089_;
  always @(posedge clk_mgated)
      ram_ff65 <= _0090_;
  always @(posedge clk_mgated)
      ram_ff66 <= _0091_;
  always @(posedge clk_mgated)
      ram_ff67 <= _0092_;
  always @(posedge clk_mgated)
      ram_ff68 <= _0093_;
  always @(posedge clk_mgated)
      ram_ff69 <= _0094_;
  always @(posedge clk_mgated)
      ram_ff70 <= _0096_;
  always @(posedge clk_mgated)
      ram_ff71 <= _0097_;
  always @(posedge clk_mgated)
      ram_ff72 <= _0098_;
  always @(posedge clk_mgated)
      ram_ff73 <= _0099_;
  always @(posedge clk_mgated)
      ram_ff74 <= _0100_;
  always @(posedge clk_mgated)
      ram_ff75 <= _0101_;
  always @(posedge clk_mgated)
      ram_ff76 <= _0102_;
  always @(posedge clk_mgated)
      ram_ff77 <= _0103_;
  always @(posedge clk_mgated)
      ram_ff78 <= _0104_;
  always @(posedge clk_mgated)
      ram_ff79 <= _0105_;
  always @(posedge clk_mgated)
      ram_ff80 <= _0107_;
  always @(posedge clk_mgated)
      ram_ff81 <= _0108_;
  always @(posedge clk_mgated)
      ram_ff82 <= _0109_;
  always @(posedge clk_mgated)
      ram_ff83 <= _0110_;
  always @(posedge clk_mgated)
      ram_ff84 <= _0111_;
  always @(posedge clk_mgated)
      ram_ff85 <= _0112_;
  always @(posedge clk_mgated)
      ram_ff86 <= _0113_;
  always @(posedge clk_mgated)
      ram_ff87 <= _0114_;
  always @(posedge clk_mgated)
      ram_ff88 <= _0115_;
  always @(posedge clk_mgated)
      ram_ff89 <= _0116_;
  always @(posedge clk_mgated)
      ram_ff90 <= _0118_;
  always @(posedge clk_mgated)
      ram_ff91 <= _0119_;
  always @(posedge clk_mgated)
      ram_ff92 <= _0120_;
  always @(posedge clk_mgated)
      ram_ff93 <= _0121_;
  always @(posedge clk_mgated)
      ram_ff94 <= _0122_;
  always @(posedge clk_mgated)
      ram_ff95 <= _0123_;
  always @(posedge clk_mgated)
      ram_ff96 <= _0124_;
  always @(posedge clk_mgated)
      ram_ff97 <= _0125_;
  always @(posedge clk_mgated)
      ram_ff98 <= _0126_;
  always @(posedge clk_mgated)
      ram_ff99 <= _0127_;
  always @(posedge clk_mgated)
      ram_ff100 <= _0002_;
  always @(posedge clk_mgated)
      ram_ff101 <= _0003_;
  always @(posedge clk_mgated)
      ram_ff102 <= _0004_;
  always @(posedge clk_mgated)
      ram_ff103 <= _0005_;
  always @(posedge clk_mgated)
      ram_ff104 <= _0006_;
  always @(posedge clk_mgated)
      ram_ff105 <= _0007_;
  always @(posedge clk_mgated)
      ram_ff106 <= _0008_;
  always @(posedge clk_mgated)
      ram_ff107 <= _0009_;
  always @(posedge clk_mgated)
      ram_ff108 <= _0010_;
  always @(posedge clk_mgated)
      ram_ff109 <= _0011_;
  always @(posedge clk_mgated)
      ram_ff110 <= _0013_;
  always @(posedge clk_mgated)
      ram_ff111 <= _0014_;
  always @(posedge clk_mgated)
      ram_ff112 <= _0015_;
  always @(posedge clk_mgated)
      ram_ff113 <= _0016_;
  always @(posedge clk_mgated)
      ram_ff114 <= _0017_;
  always @(posedge clk_mgated)
      ram_ff115 <= _0018_;
  always @(posedge clk_mgated)
      ram_ff116 <= _0019_;
  always @(posedge clk_mgated)
      ram_ff117 <= _0020_;
  always @(posedge clk_mgated)
      ram_ff118 <= _0021_;
  always @(posedge clk_mgated)
      ram_ff119 <= _0022_;
  always @(posedge clk_mgated)
      ram_ff120 <= _0024_;
  always @(posedge clk_mgated)
      ram_ff121 <= _0025_;
  always @(posedge clk_mgated)
      ram_ff122 <= _0026_;
  always @(posedge clk_mgated)
      ram_ff123 <= _0027_;
  always @(posedge clk_mgated)
      ram_ff124 <= _0028_;
  always @(posedge clk_mgated)
      ram_ff125 <= _0029_;
  always @(posedge clk_mgated)
      ram_ff126 <= _0030_;
  always @(posedge clk_mgated)
      ram_ff127 <= _0031_;
  always @(posedge clk)
      di_d <= _0000_;
  function [10:0] _0899_;
    input [10:0] a;
    input [1418:0] b;
    input [128:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:1094|./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:965" *)
    (* parallel_case *)
    casez (s)
      129'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1:
        _0899_ = b[10:0];
      129'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?:
        _0899_ = b[21:11];
      129'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??:
        _0899_ = b[32:22];
      129'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???:
        _0899_ = b[43:33];
      129'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????:
        _0899_ = b[54:44];
      129'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????:
        _0899_ = b[65:55];
      129'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????:
        _0899_ = b[76:66];
      129'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????:
        _0899_ = b[87:77];
      129'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????:
        _0899_ = b[98:88];
      129'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????:
        _0899_ = b[109:99];
      129'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????:
        _0899_ = b[120:110];
      129'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????:
        _0899_ = b[131:121];
      129'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????:
        _0899_ = b[142:132];
      129'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????:
        _0899_ = b[153:143];
      129'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????:
        _0899_ = b[164:154];
      129'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????:
        _0899_ = b[175:165];
      129'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????:
        _0899_ = b[186:176];
      129'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????:
        _0899_ = b[197:187];
      129'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????:
        _0899_ = b[208:198];
      129'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????:
        _0899_ = b[219:209];
      129'b????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????:
        _0899_ = b[230:220];
      129'b???????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????:
        _0899_ = b[241:231];
      129'b??????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????:
        _0899_ = b[252:242];
      129'b?????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????:
        _0899_ = b[263:253];
      129'b????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????:
        _0899_ = b[274:264];
      129'b???????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????:
        _0899_ = b[285:275];
      129'b??????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????:
        _0899_ = b[296:286];
      129'b?????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????:
        _0899_ = b[307:297];
      129'b????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????:
        _0899_ = b[318:308];
      129'b???????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????:
        _0899_ = b[329:319];
      129'b??????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????:
        _0899_ = b[340:330];
      129'b?????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????:
        _0899_ = b[351:341];
      129'b????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????:
        _0899_ = b[362:352];
      129'b???????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????:
        _0899_ = b[373:363];
      129'b??????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????:
        _0899_ = b[384:374];
      129'b?????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????:
        _0899_ = b[395:385];
      129'b????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????:
        _0899_ = b[406:396];
      129'b???????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????:
        _0899_ = b[417:407];
      129'b??????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????:
        _0899_ = b[428:418];
      129'b?????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????:
        _0899_ = b[439:429];
      129'b????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????:
        _0899_ = b[450:440];
      129'b???????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????:
        _0899_ = b[461:451];
      129'b??????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????:
        _0899_ = b[472:462];
      129'b?????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????:
        _0899_ = b[483:473];
      129'b????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????:
        _0899_ = b[494:484];
      129'b???????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????:
        _0899_ = b[505:495];
      129'b??????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????:
        _0899_ = b[516:506];
      129'b?????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????:
        _0899_ = b[527:517];
      129'b????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????:
        _0899_ = b[538:528];
      129'b???????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????:
        _0899_ = b[549:539];
      129'b??????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????:
        _0899_ = b[560:550];
      129'b?????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????:
        _0899_ = b[571:561];
      129'b????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????:
        _0899_ = b[582:572];
      129'b???????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????:
        _0899_ = b[593:583];
      129'b??????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????:
        _0899_ = b[604:594];
      129'b?????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????:
        _0899_ = b[615:605];
      129'b????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????:
        _0899_ = b[626:616];
      129'b???????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????:
        _0899_ = b[637:627];
      129'b??????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????:
        _0899_ = b[648:638];
      129'b?????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????:
        _0899_ = b[659:649];
      129'b????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????:
        _0899_ = b[670:660];
      129'b???????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????:
        _0899_ = b[681:671];
      129'b??????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????:
        _0899_ = b[692:682];
      129'b?????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????:
        _0899_ = b[703:693];
      129'b????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????:
        _0899_ = b[714:704];
      129'b???????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????:
        _0899_ = b[725:715];
      129'b??????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????:
        _0899_ = b[736:726];
      129'b?????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????:
        _0899_ = b[747:737];
      129'b????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????:
        _0899_ = b[758:748];
      129'b???????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????:
        _0899_ = b[769:759];
      129'b??????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????:
        _0899_ = b[780:770];
      129'b?????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????:
        _0899_ = b[791:781];
      129'b????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????:
        _0899_ = b[802:792];
      129'b???????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????:
        _0899_ = b[813:803];
      129'b??????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????:
        _0899_ = b[824:814];
      129'b?????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????:
        _0899_ = b[835:825];
      129'b????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????:
        _0899_ = b[846:836];
      129'b???????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????:
        _0899_ = b[857:847];
      129'b??????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????:
        _0899_ = b[868:858];
      129'b?????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????:
        _0899_ = b[879:869];
      129'b????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????:
        _0899_ = b[890:880];
      129'b???????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????:
        _0899_ = b[901:891];
      129'b??????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????:
        _0899_ = b[912:902];
      129'b?????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????:
        _0899_ = b[923:913];
      129'b????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????:
        _0899_ = b[934:924];
      129'b???????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????:
        _0899_ = b[945:935];
      129'b??????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????:
        _0899_ = b[956:946];
      129'b?????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????:
        _0899_ = b[967:957];
      129'b????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????:
        _0899_ = b[978:968];
      129'b???????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????:
        _0899_ = b[989:979];
      129'b??????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????:
        _0899_ = b[1000:990];
      129'b?????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????:
        _0899_ = b[1011:1001];
      129'b????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????:
        _0899_ = b[1022:1012];
      129'b???????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????:
        _0899_ = b[1033:1023];
      129'b??????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????:
        _0899_ = b[1044:1034];
      129'b?????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????:
        _0899_ = b[1055:1045];
      129'b????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????:
        _0899_ = b[1066:1056];
      129'b???????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????:
        _0899_ = b[1077:1067];
      129'b??????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????:
        _0899_ = b[1088:1078];
      129'b?????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????:
        _0899_ = b[1099:1089];
      129'b????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????:
        _0899_ = b[1110:1100];
      129'b???????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????:
        _0899_ = b[1121:1111];
      129'b??????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????:
        _0899_ = b[1132:1122];
      129'b?????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????:
        _0899_ = b[1143:1133];
      129'b????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _0899_ = b[1154:1144];
      129'b???????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _0899_ = b[1165:1155];
      129'b??????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _0899_ = b[1176:1166];
      129'b?????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _0899_ = b[1187:1177];
      129'b????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _0899_ = b[1198:1188];
      129'b???????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _0899_ = b[1209:1199];
      129'b??????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _0899_ = b[1220:1210];
      129'b?????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _0899_ = b[1231:1221];
      129'b????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _0899_ = b[1242:1232];
      129'b???????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _0899_ = b[1253:1243];
      129'b??????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _0899_ = b[1264:1254];
      129'b?????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _0899_ = b[1275:1265];
      129'b????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _0899_ = b[1286:1276];
      129'b???????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _0899_ = b[1297:1287];
      129'b??????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _0899_ = b[1308:1298];
      129'b?????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _0899_ = b[1319:1309];
      129'b????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _0899_ = b[1330:1320];
      129'b???????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _0899_ = b[1341:1331];
      129'b??????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _0899_ = b[1352:1342];
      129'b?????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _0899_ = b[1363:1353];
      129'b????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _0899_ = b[1374:1364];
      129'b???1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _0899_ = b[1385:1375];
      129'b??1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _0899_ = b[1396:1386];
      129'b?1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _0899_ = b[1407:1397];
      129'b1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _0899_ = b[1418:1408];
      default:
        _0899_ = a;
    endcase
  endfunction
  assign dout = _0899_(11'b00000000000, { ram_ff0, ram_ff1, ram_ff2, ram_ff3, ram_ff4, ram_ff5, ram_ff6, ram_ff7, ram_ff8, ram_ff9, ram_ff10, ram_ff11, ram_ff12, ram_ff13, ram_ff14, ram_ff15, ram_ff16, ram_ff17, ram_ff18, ram_ff19, ram_ff20, ram_ff21, ram_ff22, ram_ff23, ram_ff24, ram_ff25, ram_ff26, ram_ff27, ram_ff28, ram_ff29, ram_ff30, ram_ff31, ram_ff32, ram_ff33, ram_ff34, ram_ff35, ram_ff36, ram_ff37, ram_ff38, ram_ff39, ram_ff40, ram_ff41, ram_ff42, ram_ff43, ram_ff44, ram_ff45, ram_ff46, ram_ff47, ram_ff48, ram_ff49, ram_ff50, ram_ff51, ram_ff52, ram_ff53, ram_ff54, ram_ff55, ram_ff56, ram_ff57, ram_ff58, ram_ff59, ram_ff60, ram_ff61, ram_ff62, ram_ff63, ram_ff64, ram_ff65, ram_ff66, ram_ff67, ram_ff68, ram_ff69, ram_ff70, ram_ff71, ram_ff72, ram_ff73, ram_ff74, ram_ff75, ram_ff76, ram_ff77, ram_ff78, ram_ff79, ram_ff80, ram_ff81, ram_ff82, ram_ff83, ram_ff84, ram_ff85, ram_ff86, ram_ff87, ram_ff88, ram_ff89, ram_ff90, ram_ff91, ram_ff92, ram_ff93, ram_ff94, ram_ff95, ram_ff96, ram_ff97, ram_ff98, ram_ff99, ram_ff100, ram_ff101, ram_ff102, ram_ff103, ram_ff104, ram_ff105, ram_ff106, ram_ff107, ram_ff108, ram_ff109, ram_ff110, ram_ff111, ram_ff112, ram_ff113, ram_ff114, ram_ff115, ram_ff116, ram_ff117, ram_ff118, ram_ff119, ram_ff120, ram_ff121, ram_ff122, ram_ff123, ram_ff124, ram_ff125, ram_ff126, ram_ff127, di_d }, { _0513_, _0512_, _0511_, _0510_, _0509_, _0508_, _0507_, _0506_, _0505_, _0504_, _0503_, _0502_, _0501_, _0500_, _0499_, _0498_, _0497_, _0496_, _0495_, _0494_, _0493_, _0492_, _0491_, _0490_, _0489_, _0488_, _0487_, _0486_, _0485_, _0484_, _0483_, _0482_, _0481_, _0480_, _0479_, _0478_, _0477_, _0476_, _0475_, _0474_, _0473_, _0472_, _0471_, _0470_, _0469_, _0468_, _0467_, _0466_, _0465_, _0464_, _0463_, _0462_, _0461_, _0460_, _0459_, _0458_, _0457_, _0456_, _0455_, _0454_, _0453_, _0452_, _0451_, _0450_, _0449_, _0448_, _0447_, _0446_, _0445_, _0444_, _0443_, _0442_, _0441_, _0440_, _0439_, _0438_, _0437_, _0436_, _0435_, _0434_, _0433_, _0432_, _0431_, _0430_, _0429_, _0428_, _0427_, _0426_, _0425_, _0424_, _0423_, _0422_, _0421_, _0420_, _0419_, _0418_, _0417_, _0416_, _0415_, _0414_, _0413_, _0412_, _0411_, _0410_, _0409_, _0408_, _0407_, _0406_, _0405_, _0404_, _0403_, _0402_, _0401_, _0400_, _0399_, _0398_, _0397_, _0396_, _0395_, _0394_, _0393_, _0392_, _0391_, _0390_, _0389_, _0388_, _0387_, _0386_, _0385_ });
  assign _0385_ = ra == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:1094|./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:965" *) 8'b10000000;
  assign _0386_ = ra == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:1093|./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:965" *) 7'b1111111;
  assign _0387_ = ra == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:1092|./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:965" *) 7'b1111110;
  assign _0388_ = ra == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:1091|./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:965" *) 7'b1111101;
  assign _0389_ = ra == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:1090|./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:965" *) 7'b1111100;
  assign _0390_ = ra == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:1089|./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:965" *) 7'b1111011;
  assign _0391_ = ra == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:1088|./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:965" *) 7'b1111010;
  assign _0392_ = ra == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:1087|./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:965" *) 7'b1111001;
  assign _0393_ = ra == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:1086|./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:965" *) 7'b1111000;
  assign _0394_ = ra == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:1085|./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:965" *) 7'b1110111;
  assign _0395_ = ra == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:1084|./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:965" *) 7'b1110110;
  assign _0396_ = ra == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:1083|./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:965" *) 7'b1110101;
  assign _0397_ = ra == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:1082|./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:965" *) 7'b1110100;
  assign _0398_ = ra == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:1081|./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:965" *) 7'b1110011;
  assign _0399_ = ra == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:1080|./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:965" *) 7'b1110010;
  assign _0400_ = ra == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:1079|./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:965" *) 7'b1110001;
  assign _0401_ = ra == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:1078|./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:965" *) 7'b1110000;
  assign _0402_ = ra == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:1077|./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:965" *) 7'b1101111;
  assign _0403_ = ra == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:1076|./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:965" *) 7'b1101110;
  assign _0404_ = ra == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:1075|./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:965" *) 7'b1101101;
  assign _0405_ = ra == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:1074|./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:965" *) 7'b1101100;
  assign _0406_ = ra == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:1073|./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:965" *) 7'b1101011;
  assign _0407_ = ra == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:1072|./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:965" *) 7'b1101010;
  assign _0408_ = ra == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:1071|./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:965" *) 7'b1101001;
  assign _0409_ = ra == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:1070|./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:965" *) 7'b1101000;
  assign _0410_ = ra == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:1069|./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:965" *) 7'b1100111;
  assign _0411_ = ra == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:1068|./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:965" *) 7'b1100110;
  assign _0412_ = ra == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:1067|./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:965" *) 7'b1100101;
  assign _0413_ = ra == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:1066|./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:965" *) 7'b1100100;
  assign _0414_ = ra == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:1065|./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:965" *) 7'b1100011;
  assign _0415_ = ra == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:1064|./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:965" *) 7'b1100010;
  assign _0416_ = ra == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:1063|./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:965" *) 7'b1100001;
  assign _0417_ = ra == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:1062|./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:965" *) 7'b1100000;
  assign _0418_ = ra == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:1061|./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:965" *) 7'b1011111;
  assign _0419_ = ra == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:1060|./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:965" *) 7'b1011110;
  assign _0420_ = ra == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:1059|./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:965" *) 7'b1011101;
  assign _0421_ = ra == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:1058|./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:965" *) 7'b1011100;
  assign _0422_ = ra == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:1057|./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:965" *) 7'b1011011;
  assign _0423_ = ra == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:1056|./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:965" *) 7'b1011010;
  assign _0424_ = ra == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:1055|./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:965" *) 7'b1011001;
  assign _0425_ = ra == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:1054|./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:965" *) 7'b1011000;
  assign _0426_ = ra == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:1053|./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:965" *) 7'b1010111;
  assign _0427_ = ra == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:1052|./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:965" *) 7'b1010110;
  assign _0428_ = ra == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:1051|./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:965" *) 7'b1010101;
  assign _0429_ = ra == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:1050|./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:965" *) 7'b1010100;
  assign _0430_ = ra == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:1049|./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:965" *) 7'b1010011;
  assign _0431_ = ra == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:1048|./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:965" *) 7'b1010010;
  assign _0432_ = ra == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:1047|./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:965" *) 7'b1010001;
  assign _0433_ = ra == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:1046|./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:965" *) 7'b1010000;
  assign _0434_ = ra == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:1045|./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:965" *) 7'b1001111;
  assign _0435_ = ra == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:1044|./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:965" *) 7'b1001110;
  assign _0436_ = ra == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:1043|./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:965" *) 7'b1001101;
  assign _0437_ = ra == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:1042|./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:965" *) 7'b1001100;
  assign _0438_ = ra == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:1041|./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:965" *) 7'b1001011;
  assign _0439_ = ra == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:1040|./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:965" *) 7'b1001010;
  assign _0440_ = ra == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:1039|./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:965" *) 7'b1001001;
  assign _0441_ = ra == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:1038|./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:965" *) 7'b1001000;
  assign _0442_ = ra == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:1037|./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:965" *) 7'b1000111;
  assign _0443_ = ra == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:1036|./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:965" *) 7'b1000110;
  assign _0444_ = ra == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:1035|./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:965" *) 7'b1000101;
  assign _0445_ = ra == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:1034|./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:965" *) 7'b1000100;
  assign _0446_ = ra == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:1033|./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:965" *) 7'b1000011;
  assign _0447_ = ra == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:1032|./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:965" *) 7'b1000010;
  assign _0448_ = ra == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:1031|./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:965" *) 7'b1000001;
  assign _0449_ = ra == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:1030|./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:965" *) 7'b1000000;
  assign _0450_ = ra == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:1029|./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:965" *) 6'b111111;
  assign _0451_ = ra == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:1028|./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:965" *) 6'b111110;
  assign _0452_ = ra == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:1027|./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:965" *) 6'b111101;
  assign _0453_ = ra == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:1026|./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:965" *) 6'b111100;
  assign _0454_ = ra == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:1025|./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:965" *) 6'b111011;
  assign _0455_ = ra == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:1024|./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:965" *) 6'b111010;
  assign _0456_ = ra == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:1023|./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:965" *) 6'b111001;
  assign _0457_ = ra == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:1022|./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:965" *) 6'b111000;
  assign _0458_ = ra == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:1021|./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:965" *) 6'b110111;
  assign _0459_ = ra == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:1020|./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:965" *) 6'b110110;
  assign _0460_ = ra == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:1019|./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:965" *) 6'b110101;
  assign _0461_ = ra == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:1018|./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:965" *) 6'b110100;
  assign _0462_ = ra == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:1017|./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:965" *) 6'b110011;
  assign _0463_ = ra == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:1016|./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:965" *) 6'b110010;
  assign _0464_ = ra == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:1015|./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:965" *) 6'b110001;
  assign _0465_ = ra == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:1014|./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:965" *) 6'b110000;
  assign _0466_ = ra == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:1013|./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:965" *) 6'b101111;
  assign _0467_ = ra == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:1012|./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:965" *) 6'b101110;
  assign _0468_ = ra == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:1011|./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:965" *) 6'b101101;
  assign _0469_ = ra == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:1010|./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:965" *) 6'b101100;
  assign _0470_ = ra == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:1009|./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:965" *) 6'b101011;
  assign _0471_ = ra == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:1008|./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:965" *) 6'b101010;
  assign _0472_ = ra == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:1007|./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:965" *) 6'b101001;
  assign _0473_ = ra == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:1006|./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:965" *) 6'b101000;
  assign _0474_ = ra == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:1005|./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:965" *) 6'b100111;
  assign _0475_ = ra == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:1004|./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:965" *) 6'b100110;
  assign _0476_ = ra == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:1003|./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:965" *) 6'b100101;
  assign _0477_ = ra == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:1002|./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:965" *) 6'b100100;
  assign _0478_ = ra == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:1001|./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:965" *) 6'b100011;
  assign _0479_ = ra == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:1000|./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:965" *) 6'b100010;
  assign _0480_ = ra == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:999|./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:965" *) 6'b100001;
  assign _0481_ = ra == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:998|./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:965" *) 6'b100000;
  assign _0482_ = ra == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:997|./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:965" *) 5'b11111;
  assign _0483_ = ra == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:996|./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:965" *) 5'b11110;
  assign _0484_ = ra == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:995|./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:965" *) 5'b11101;
  assign _0485_ = ra == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:994|./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:965" *) 5'b11100;
  assign _0486_ = ra == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:993|./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:965" *) 5'b11011;
  assign _0487_ = ra == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:992|./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:965" *) 5'b11010;
  assign _0488_ = ra == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:991|./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:965" *) 5'b11001;
  assign _0489_ = ra == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:990|./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:965" *) 5'b11000;
  assign _0490_ = ra == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:989|./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:965" *) 5'b10111;
  assign _0491_ = ra == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:988|./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:965" *) 5'b10110;
  assign _0492_ = ra == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:987|./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:965" *) 5'b10101;
  assign _0493_ = ra == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:986|./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:965" *) 5'b10100;
  assign _0494_ = ra == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:985|./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:965" *) 5'b10011;
  assign _0495_ = ra == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:984|./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:965" *) 5'b10010;
  assign _0496_ = ra == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:983|./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:965" *) 5'b10001;
  assign _0497_ = ra == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:982|./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:965" *) 5'b10000;
  assign _0498_ = ra == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:981|./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:965" *) 4'b1111;
  assign _0499_ = ra == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:980|./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:965" *) 4'b1110;
  assign _0500_ = ra == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:979|./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:965" *) 4'b1101;
  assign _0501_ = ra == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:978|./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:965" *) 4'b1100;
  assign _0502_ = ra == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:977|./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:965" *) 4'b1011;
  assign _0503_ = ra == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:976|./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:965" *) 4'b1010;
  assign _0504_ = ra == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:975|./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:965" *) 4'b1001;
  assign _0505_ = ra == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:974|./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:965" *) 4'b1000;
  assign _0506_ = ra == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:973|./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:965" *) 3'b111;
  assign _0507_ = ra == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:972|./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:965" *) 3'b110;
  assign _0508_ = ra == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:971|./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:965" *) 3'b101;
  assign _0509_ = ra == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:970|./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:965" *) 3'b100;
  assign _0510_ = ra == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:969|./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:965" *) 2'b11;
  assign _0511_ = ra == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:968|./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:965" *) 2'b10;
  assign _0512_ = ra == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:967|./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:965" *) 1'b1;
  assign _0513_ = ! (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:966|./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:965" *) ra;
  assign _0031_ = _0384_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:959" *) di_d : ram_ff127;
  assign _0030_ = _0383_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:956" *) di_d : ram_ff126;
  assign _0029_ = _0382_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:953" *) di_d : ram_ff125;
  assign _0028_ = _0381_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:950" *) di_d : ram_ff124;
  assign _0027_ = _0380_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:947" *) di_d : ram_ff123;
  assign _0026_ = _0379_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:944" *) di_d : ram_ff122;
  assign _0025_ = _0378_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:941" *) di_d : ram_ff121;
  assign _0024_ = _0377_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:938" *) di_d : ram_ff120;
  assign _0022_ = _0376_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:935" *) di_d : ram_ff119;
  assign _0021_ = _0375_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:932" *) di_d : ram_ff118;
  assign _0020_ = _0374_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:929" *) di_d : ram_ff117;
  assign _0019_ = _0373_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:926" *) di_d : ram_ff116;
  assign _0018_ = _0372_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:923" *) di_d : ram_ff115;
  assign _0017_ = _0371_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:920" *) di_d : ram_ff114;
  assign _0016_ = _0370_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:917" *) di_d : ram_ff113;
  assign _0015_ = _0369_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:914" *) di_d : ram_ff112;
  assign _0014_ = _0368_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:911" *) di_d : ram_ff111;
  assign _0013_ = _0367_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:908" *) di_d : ram_ff110;
  assign _0011_ = _0366_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:905" *) di_d : ram_ff109;
  assign _0010_ = _0365_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:902" *) di_d : ram_ff108;
  assign _0009_ = _0364_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:899" *) di_d : ram_ff107;
  assign _0008_ = _0363_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:896" *) di_d : ram_ff106;
  assign _0007_ = _0362_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:893" *) di_d : ram_ff105;
  assign _0006_ = _0361_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:890" *) di_d : ram_ff104;
  assign _0005_ = _0360_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:887" *) di_d : ram_ff103;
  assign _0004_ = _0359_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:884" *) di_d : ram_ff102;
  assign _0003_ = _0358_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:881" *) di_d : ram_ff101;
  assign _0002_ = _0357_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:878" *) di_d : ram_ff100;
  assign _0127_ = _0356_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:875" *) di_d : ram_ff99;
  assign _0126_ = _0355_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:872" *) di_d : ram_ff98;
  assign _0125_ = _0354_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:869" *) di_d : ram_ff97;
  assign _0124_ = _0353_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:866" *) di_d : ram_ff96;
  assign _0123_ = _0352_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:863" *) di_d : ram_ff95;
  assign _0122_ = _0351_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:860" *) di_d : ram_ff94;
  assign _0121_ = _0350_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:857" *) di_d : ram_ff93;
  assign _0120_ = _0349_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:854" *) di_d : ram_ff92;
  assign _0119_ = _0348_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:851" *) di_d : ram_ff91;
  assign _0118_ = _0347_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:848" *) di_d : ram_ff90;
  assign _0116_ = _0346_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:845" *) di_d : ram_ff89;
  assign _0115_ = _0345_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:842" *) di_d : ram_ff88;
  assign _0114_ = _0344_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:839" *) di_d : ram_ff87;
  assign _0113_ = _0343_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:836" *) di_d : ram_ff86;
  assign _0112_ = _0342_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:833" *) di_d : ram_ff85;
  assign _0111_ = _0341_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:830" *) di_d : ram_ff84;
  assign _0110_ = _0340_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:827" *) di_d : ram_ff83;
  assign _0109_ = _0339_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:824" *) di_d : ram_ff82;
  assign _0108_ = _0338_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:821" *) di_d : ram_ff81;
  assign _0107_ = _0337_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:818" *) di_d : ram_ff80;
  assign _0105_ = _0336_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:815" *) di_d : ram_ff79;
  assign _0104_ = _0335_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:812" *) di_d : ram_ff78;
  assign _0103_ = _0334_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:809" *) di_d : ram_ff77;
  assign _0102_ = _0333_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:806" *) di_d : ram_ff76;
  assign _0101_ = _0332_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:803" *) di_d : ram_ff75;
  assign _0100_ = _0331_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:800" *) di_d : ram_ff74;
  assign _0099_ = _0330_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:797" *) di_d : ram_ff73;
  assign _0098_ = _0329_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:794" *) di_d : ram_ff72;
  assign _0097_ = _0328_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:791" *) di_d : ram_ff71;
  assign _0096_ = _0327_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:788" *) di_d : ram_ff70;
  assign _0094_ = _0326_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:785" *) di_d : ram_ff69;
  assign _0093_ = _0325_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:782" *) di_d : ram_ff68;
  assign _0092_ = _0324_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:779" *) di_d : ram_ff67;
  assign _0091_ = _0323_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:776" *) di_d : ram_ff66;
  assign _0090_ = _0322_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:773" *) di_d : ram_ff65;
  assign _0089_ = _0321_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:770" *) di_d : ram_ff64;
  assign _0088_ = _0320_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:767" *) di_d : ram_ff63;
  assign _0087_ = _0319_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:764" *) di_d : ram_ff62;
  assign _0086_ = _0318_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:761" *) di_d : ram_ff61;
  assign _0085_ = _0317_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:758" *) di_d : ram_ff60;
  assign _0083_ = _0316_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:755" *) di_d : ram_ff59;
  assign _0082_ = _0315_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:752" *) di_d : ram_ff58;
  assign _0081_ = _0314_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:749" *) di_d : ram_ff57;
  assign _0080_ = _0313_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:746" *) di_d : ram_ff56;
  assign _0079_ = _0312_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:743" *) di_d : ram_ff55;
  assign _0078_ = _0311_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:740" *) di_d : ram_ff54;
  assign _0077_ = _0310_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:737" *) di_d : ram_ff53;
  assign _0076_ = _0309_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:734" *) di_d : ram_ff52;
  assign _0075_ = _0308_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:731" *) di_d : ram_ff51;
  assign _0074_ = _0307_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:728" *) di_d : ram_ff50;
  assign _0072_ = _0306_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:725" *) di_d : ram_ff49;
  assign _0071_ = _0305_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:722" *) di_d : ram_ff48;
  assign _0070_ = _0304_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:719" *) di_d : ram_ff47;
  assign _0069_ = _0303_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:716" *) di_d : ram_ff46;
  assign _0068_ = _0302_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:713" *) di_d : ram_ff45;
  assign _0067_ = _0301_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:710" *) di_d : ram_ff44;
  assign _0066_ = _0300_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:707" *) di_d : ram_ff43;
  assign _0065_ = _0299_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:704" *) di_d : ram_ff42;
  assign _0064_ = _0298_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:701" *) di_d : ram_ff41;
  assign _0063_ = _0297_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:698" *) di_d : ram_ff40;
  assign _0061_ = _0296_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:695" *) di_d : ram_ff39;
  assign _0060_ = _0295_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:692" *) di_d : ram_ff38;
  assign _0059_ = _0294_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:689" *) di_d : ram_ff37;
  assign _0058_ = _0293_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:686" *) di_d : ram_ff36;
  assign _0057_ = _0292_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:683" *) di_d : ram_ff35;
  assign _0056_ = _0291_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:680" *) di_d : ram_ff34;
  assign _0055_ = _0290_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:677" *) di_d : ram_ff33;
  assign _0054_ = _0289_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:674" *) di_d : ram_ff32;
  assign _0053_ = _0288_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:671" *) di_d : ram_ff31;
  assign _0052_ = _0287_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:668" *) di_d : ram_ff30;
  assign _0050_ = _0286_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:665" *) di_d : ram_ff29;
  assign _0049_ = _0285_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:662" *) di_d : ram_ff28;
  assign _0048_ = _0284_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:659" *) di_d : ram_ff27;
  assign _0047_ = _0283_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:656" *) di_d : ram_ff26;
  assign _0046_ = _0282_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:653" *) di_d : ram_ff25;
  assign _0045_ = _0281_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:650" *) di_d : ram_ff24;
  assign _0044_ = _0280_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:647" *) di_d : ram_ff23;
  assign _0043_ = _0279_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:644" *) di_d : ram_ff22;
  assign _0042_ = _0278_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:641" *) di_d : ram_ff21;
  assign _0041_ = _0277_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:638" *) di_d : ram_ff20;
  assign _0039_ = _0276_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:635" *) di_d : ram_ff19;
  assign _0038_ = _0275_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:632" *) di_d : ram_ff18;
  assign _0037_ = _0274_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:629" *) di_d : ram_ff17;
  assign _0036_ = _0273_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:626" *) di_d : ram_ff16;
  assign _0035_ = _0272_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:623" *) di_d : ram_ff15;
  assign _0034_ = _0271_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:620" *) di_d : ram_ff14;
  assign _0033_ = _0270_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:617" *) di_d : ram_ff13;
  assign _0032_ = _0269_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:614" *) di_d : ram_ff12;
  assign _0023_ = _0268_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:611" *) di_d : ram_ff11;
  assign _0012_ = _0267_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:608" *) di_d : ram_ff10;
  assign _0128_ = _0266_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:605" *) di_d : ram_ff9;
  assign _0117_ = _0265_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:602" *) di_d : ram_ff8;
  assign _0106_ = _0264_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:599" *) di_d : ram_ff7;
  assign _0095_ = _0263_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:596" *) di_d : ram_ff6;
  assign _0084_ = _0262_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:593" *) di_d : ram_ff5;
  assign _0073_ = _0261_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:590" *) di_d : ram_ff4;
  assign _0062_ = _0260_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:587" *) di_d : ram_ff3;
  assign _0051_ = _0259_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:584" *) di_d : ram_ff2;
  assign _0040_ = _0258_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:581" *) di_d : ram_ff1;
  assign _0001_ = _0257_ ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:578" *) di_d : ram_ff0;
  assign _0000_ = iwe ? (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_IMG_sg2pack_fifo.v:423" *) di : di_d;
endmodule
