module SDP_X_chn_alu_out_rsci_unreg(in_0, outsig);
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:955" *)
  input in_0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:956" *)
  output outsig;
  assign outsig = in_0;
endmodule
