module one_round(clk, state_in, key, state_out);
  wire [7:0] _0000_;
  wire _0001_;
  wire _0002_;
  wire _0003_;
  wire _0004_;
  wire _0005_;
  wire _0006_;
  wire _0007_;
  wire _0008_;
  wire _0009_;
  wire _0010_;
  wire _0011_;
  wire _0012_;
  wire _0013_;
  wire _0014_;
  wire _0015_;
  wire _0016_;
  wire _0017_;
  wire _0018_;
  wire _0019_;
  wire _0020_;
  wire _0021_;
  wire _0022_;
  wire _0023_;
  wire _0024_;
  wire _0025_;
  wire _0026_;
  wire _0027_;
  wire _0028_;
  wire _0029_;
  wire _0030_;
  wire _0031_;
  wire _0032_;
  wire _0033_;
  wire _0034_;
  wire _0035_;
  wire _0036_;
  wire _0037_;
  wire _0038_;
  wire _0039_;
  wire _0040_;
  wire _0041_;
  wire _0042_;
  wire _0043_;
  wire _0044_;
  wire _0045_;
  wire _0046_;
  wire _0047_;
  wire _0048_;
  wire _0049_;
  wire _0050_;
  wire _0051_;
  wire _0052_;
  wire _0053_;
  wire _0054_;
  wire _0055_;
  wire _0056_;
  wire _0057_;
  wire _0058_;
  wire _0059_;
  wire _0060_;
  wire _0061_;
  wire _0062_;
  wire _0063_;
  wire _0064_;
  wire _0065_;
  wire _0066_;
  wire _0067_;
  wire _0068_;
  wire _0069_;
  wire _0070_;
  wire _0071_;
  wire _0072_;
  wire _0073_;
  wire _0074_;
  wire _0075_;
  wire _0076_;
  wire _0077_;
  wire _0078_;
  wire _0079_;
  wire _0080_;
  wire _0081_;
  wire _0082_;
  wire _0083_;
  wire _0084_;
  wire _0085_;
  wire _0086_;
  wire _0087_;
  wire _0088_;
  wire _0089_;
  wire _0090_;
  wire _0091_;
  wire _0092_;
  wire _0093_;
  wire _0094_;
  wire _0095_;
  wire _0096_;
  wire _0097_;
  wire _0098_;
  wire _0099_;
  wire _0100_;
  wire _0101_;
  wire _0102_;
  wire _0103_;
  wire _0104_;
  wire _0105_;
  wire _0106_;
  wire _0107_;
  wire _0108_;
  wire _0109_;
  wire _0110_;
  wire _0111_;
  wire _0112_;
  wire _0113_;
  wire _0114_;
  wire _0115_;
  wire _0116_;
  wire _0117_;
  wire _0118_;
  wire _0119_;
  wire _0120_;
  wire _0121_;
  wire _0122_;
  wire _0123_;
  wire _0124_;
  wire _0125_;
  wire _0126_;
  wire _0127_;
  wire _0128_;
  wire _0129_;
  wire _0130_;
  wire _0131_;
  wire _0132_;
  wire _0133_;
  wire _0134_;
  wire _0135_;
  wire _0136_;
  wire _0137_;
  wire _0138_;
  wire _0139_;
  wire _0140_;
  wire _0141_;
  wire _0142_;
  wire _0143_;
  wire _0144_;
  wire _0145_;
  wire _0146_;
  wire _0147_;
  wire _0148_;
  wire _0149_;
  wire _0150_;
  wire _0151_;
  wire _0152_;
  wire _0153_;
  wire _0154_;
  wire _0155_;
  wire _0156_;
  wire _0157_;
  wire _0158_;
  wire _0159_;
  wire _0160_;
  wire _0161_;
  wire _0162_;
  wire _0163_;
  wire _0164_;
  wire _0165_;
  wire _0166_;
  wire _0167_;
  wire _0168_;
  wire _0169_;
  wire _0170_;
  wire _0171_;
  wire _0172_;
  wire _0173_;
  wire _0174_;
  wire _0175_;
  wire _0176_;
  wire _0177_;
  wire _0178_;
  wire _0179_;
  wire _0180_;
  wire _0181_;
  wire _0182_;
  wire _0183_;
  wire _0184_;
  wire _0185_;
  wire _0186_;
  wire _0187_;
  wire _0188_;
  wire _0189_;
  wire _0190_;
  wire _0191_;
  wire _0192_;
  wire _0193_;
  wire _0194_;
  wire _0195_;
  wire _0196_;
  wire _0197_;
  wire _0198_;
  wire _0199_;
  wire _0200_;
  wire _0201_;
  wire _0202_;
  wire _0203_;
  wire _0204_;
  wire _0205_;
  wire _0206_;
  wire _0207_;
  wire _0208_;
  wire _0209_;
  wire _0210_;
  wire _0211_;
  wire _0212_;
  wire _0213_;
  wire _0214_;
  wire _0215_;
  wire _0216_;
  wire _0217_;
  wire _0218_;
  wire _0219_;
  wire _0220_;
  wire _0221_;
  wire _0222_;
  wire _0223_;
  wire _0224_;
  wire _0225_;
  wire _0226_;
  wire _0227_;
  wire _0228_;
  wire _0229_;
  wire _0230_;
  wire _0231_;
  wire _0232_;
  wire _0233_;
  wire _0234_;
  wire _0235_;
  wire _0236_;
  wire _0237_;
  wire _0238_;
  wire _0239_;
  wire _0240_;
  wire _0241_;
  wire _0242_;
  wire _0243_;
  wire _0244_;
  wire _0245_;
  wire _0246_;
  wire _0247_;
  wire _0248_;
  wire _0249_;
  wire _0250_;
  wire _0251_;
  wire _0252_;
  wire _0253_;
  wire _0254_;
  wire _0255_;
  wire _0256_;
  wire [7:0] _0257_;
  wire [7:0] _0258_;
  wire _0259_;
  wire _0260_;
  wire _0261_;
  wire _0262_;
  wire _0263_;
  wire _0264_;
  wire _0265_;
  wire _0266_;
  wire _0267_;
  wire _0268_;
  wire _0269_;
  wire _0270_;
  wire _0271_;
  wire _0272_;
  wire _0273_;
  wire _0274_;
  wire _0275_;
  wire _0276_;
  wire _0277_;
  wire _0278_;
  wire _0279_;
  wire _0280_;
  wire _0281_;
  wire _0282_;
  wire _0283_;
  wire _0284_;
  wire _0285_;
  wire _0286_;
  wire _0287_;
  wire _0288_;
  wire _0289_;
  wire _0290_;
  wire _0291_;
  wire _0292_;
  wire _0293_;
  wire _0294_;
  wire _0295_;
  wire _0296_;
  wire _0297_;
  wire _0298_;
  wire _0299_;
  wire _0300_;
  wire _0301_;
  wire _0302_;
  wire _0303_;
  wire _0304_;
  wire _0305_;
  wire _0306_;
  wire _0307_;
  wire _0308_;
  wire _0309_;
  wire _0310_;
  wire _0311_;
  wire _0312_;
  wire _0313_;
  wire _0314_;
  wire _0315_;
  wire _0316_;
  wire _0317_;
  wire _0318_;
  wire _0319_;
  wire _0320_;
  wire _0321_;
  wire _0322_;
  wire _0323_;
  wire _0324_;
  wire _0325_;
  wire _0326_;
  wire _0327_;
  wire _0328_;
  wire _0329_;
  wire _0330_;
  wire _0331_;
  wire _0332_;
  wire _0333_;
  wire _0334_;
  wire _0335_;
  wire _0336_;
  wire _0337_;
  wire _0338_;
  wire _0339_;
  wire _0340_;
  wire _0341_;
  wire _0342_;
  wire _0343_;
  wire _0344_;
  wire _0345_;
  wire _0346_;
  wire _0347_;
  wire _0348_;
  wire _0349_;
  wire _0350_;
  wire _0351_;
  wire _0352_;
  wire _0353_;
  wire _0354_;
  wire _0355_;
  wire _0356_;
  wire _0357_;
  wire _0358_;
  wire _0359_;
  wire _0360_;
  wire _0361_;
  wire _0362_;
  wire _0363_;
  wire _0364_;
  wire _0365_;
  wire _0366_;
  wire _0367_;
  wire _0368_;
  wire _0369_;
  wire _0370_;
  wire _0371_;
  wire _0372_;
  wire _0373_;
  wire _0374_;
  wire _0375_;
  wire _0376_;
  wire _0377_;
  wire _0378_;
  wire _0379_;
  wire _0380_;
  wire _0381_;
  wire _0382_;
  wire _0383_;
  wire _0384_;
  wire _0385_;
  wire _0386_;
  wire _0387_;
  wire _0388_;
  wire _0389_;
  wire _0390_;
  wire _0391_;
  wire _0392_;
  wire _0393_;
  wire _0394_;
  wire _0395_;
  wire _0396_;
  wire _0397_;
  wire _0398_;
  wire _0399_;
  wire _0400_;
  wire _0401_;
  wire _0402_;
  wire _0403_;
  wire _0404_;
  wire _0405_;
  wire _0406_;
  wire _0407_;
  wire _0408_;
  wire _0409_;
  wire _0410_;
  wire _0411_;
  wire _0412_;
  wire _0413_;
  wire _0414_;
  wire _0415_;
  wire _0416_;
  wire _0417_;
  wire _0418_;
  wire _0419_;
  wire _0420_;
  wire _0421_;
  wire _0422_;
  wire _0423_;
  wire _0424_;
  wire _0425_;
  wire _0426_;
  wire _0427_;
  wire _0428_;
  wire _0429_;
  wire _0430_;
  wire _0431_;
  wire _0432_;
  wire _0433_;
  wire _0434_;
  wire _0435_;
  wire _0436_;
  wire _0437_;
  wire _0438_;
  wire _0439_;
  wire _0440_;
  wire _0441_;
  wire _0442_;
  wire _0443_;
  wire _0444_;
  wire _0445_;
  wire _0446_;
  wire _0447_;
  wire _0448_;
  wire _0449_;
  wire _0450_;
  wire _0451_;
  wire _0452_;
  wire _0453_;
  wire _0454_;
  wire _0455_;
  wire _0456_;
  wire _0457_;
  wire _0458_;
  wire _0459_;
  wire _0460_;
  wire _0461_;
  wire _0462_;
  wire _0463_;
  wire _0464_;
  wire _0465_;
  wire _0466_;
  wire _0467_;
  wire _0468_;
  wire _0469_;
  wire _0470_;
  wire _0471_;
  wire _0472_;
  wire _0473_;
  wire _0474_;
  wire _0475_;
  wire _0476_;
  wire _0477_;
  wire _0478_;
  wire _0479_;
  wire _0480_;
  wire _0481_;
  wire _0482_;
  wire _0483_;
  wire _0484_;
  wire _0485_;
  wire _0486_;
  wire _0487_;
  wire _0488_;
  wire _0489_;
  wire _0490_;
  wire _0491_;
  wire _0492_;
  wire _0493_;
  wire _0494_;
  wire _0495_;
  wire _0496_;
  wire _0497_;
  wire _0498_;
  wire _0499_;
  wire _0500_;
  wire _0501_;
  wire _0502_;
  wire _0503_;
  wire _0504_;
  wire _0505_;
  wire _0506_;
  wire _0507_;
  wire _0508_;
  wire _0509_;
  wire _0510_;
  wire _0511_;
  wire _0512_;
  wire _0513_;
  wire _0514_;
  wire [7:0] _0515_;
  wire [7:0] _0516_;
  wire _0517_;
  wire _0518_;
  wire _0519_;
  wire _0520_;
  wire _0521_;
  wire _0522_;
  wire _0523_;
  wire _0524_;
  wire _0525_;
  wire _0526_;
  wire _0527_;
  wire _0528_;
  wire _0529_;
  wire _0530_;
  wire _0531_;
  wire _0532_;
  wire _0533_;
  wire _0534_;
  wire _0535_;
  wire _0536_;
  wire _0537_;
  wire _0538_;
  wire _0539_;
  wire _0540_;
  wire _0541_;
  wire _0542_;
  wire _0543_;
  wire _0544_;
  wire _0545_;
  wire _0546_;
  wire _0547_;
  wire _0548_;
  wire _0549_;
  wire _0550_;
  wire _0551_;
  wire _0552_;
  wire _0553_;
  wire _0554_;
  wire _0555_;
  wire _0556_;
  wire _0557_;
  wire _0558_;
  wire _0559_;
  wire _0560_;
  wire _0561_;
  wire _0562_;
  wire _0563_;
  wire _0564_;
  wire _0565_;
  wire _0566_;
  wire _0567_;
  wire _0568_;
  wire _0569_;
  wire _0570_;
  wire _0571_;
  wire _0572_;
  wire _0573_;
  wire _0574_;
  wire _0575_;
  wire _0576_;
  wire _0577_;
  wire _0578_;
  wire _0579_;
  wire _0580_;
  wire _0581_;
  wire _0582_;
  wire _0583_;
  wire _0584_;
  wire _0585_;
  wire _0586_;
  wire _0587_;
  wire _0588_;
  wire _0589_;
  wire _0590_;
  wire _0591_;
  wire _0592_;
  wire _0593_;
  wire _0594_;
  wire _0595_;
  wire _0596_;
  wire _0597_;
  wire _0598_;
  wire _0599_;
  wire _0600_;
  wire _0601_;
  wire _0602_;
  wire _0603_;
  wire _0604_;
  wire _0605_;
  wire _0606_;
  wire _0607_;
  wire _0608_;
  wire _0609_;
  wire _0610_;
  wire _0611_;
  wire _0612_;
  wire _0613_;
  wire _0614_;
  wire _0615_;
  wire _0616_;
  wire _0617_;
  wire _0618_;
  wire _0619_;
  wire _0620_;
  wire _0621_;
  wire _0622_;
  wire _0623_;
  wire _0624_;
  wire _0625_;
  wire _0626_;
  wire _0627_;
  wire _0628_;
  wire _0629_;
  wire _0630_;
  wire _0631_;
  wire _0632_;
  wire _0633_;
  wire _0634_;
  wire _0635_;
  wire _0636_;
  wire _0637_;
  wire _0638_;
  wire _0639_;
  wire _0640_;
  wire _0641_;
  wire _0642_;
  wire _0643_;
  wire _0644_;
  wire _0645_;
  wire _0646_;
  wire _0647_;
  wire _0648_;
  wire _0649_;
  wire _0650_;
  wire _0651_;
  wire _0652_;
  wire _0653_;
  wire _0654_;
  wire _0655_;
  wire _0656_;
  wire _0657_;
  wire _0658_;
  wire _0659_;
  wire _0660_;
  wire _0661_;
  wire _0662_;
  wire _0663_;
  wire _0664_;
  wire _0665_;
  wire _0666_;
  wire _0667_;
  wire _0668_;
  wire _0669_;
  wire _0670_;
  wire _0671_;
  wire _0672_;
  wire _0673_;
  wire _0674_;
  wire _0675_;
  wire _0676_;
  wire _0677_;
  wire _0678_;
  wire _0679_;
  wire _0680_;
  wire _0681_;
  wire _0682_;
  wire _0683_;
  wire _0684_;
  wire _0685_;
  wire _0686_;
  wire _0687_;
  wire _0688_;
  wire _0689_;
  wire _0690_;
  wire _0691_;
  wire _0692_;
  wire _0693_;
  wire _0694_;
  wire _0695_;
  wire _0696_;
  wire _0697_;
  wire _0698_;
  wire _0699_;
  wire _0700_;
  wire _0701_;
  wire _0702_;
  wire _0703_;
  wire _0704_;
  wire _0705_;
  wire _0706_;
  wire _0707_;
  wire _0708_;
  wire _0709_;
  wire _0710_;
  wire _0711_;
  wire _0712_;
  wire _0713_;
  wire _0714_;
  wire _0715_;
  wire _0716_;
  wire _0717_;
  wire _0718_;
  wire _0719_;
  wire _0720_;
  wire _0721_;
  wire _0722_;
  wire _0723_;
  wire _0724_;
  wire _0725_;
  wire _0726_;
  wire _0727_;
  wire _0728_;
  wire _0729_;
  wire _0730_;
  wire _0731_;
  wire _0732_;
  wire _0733_;
  wire _0734_;
  wire _0735_;
  wire _0736_;
  wire _0737_;
  wire _0738_;
  wire _0739_;
  wire _0740_;
  wire _0741_;
  wire _0742_;
  wire _0743_;
  wire _0744_;
  wire _0745_;
  wire _0746_;
  wire _0747_;
  wire _0748_;
  wire _0749_;
  wire _0750_;
  wire _0751_;
  wire _0752_;
  wire _0753_;
  wire _0754_;
  wire _0755_;
  wire _0756_;
  wire _0757_;
  wire _0758_;
  wire _0759_;
  wire _0760_;
  wire _0761_;
  wire _0762_;
  wire _0763_;
  wire _0764_;
  wire _0765_;
  wire _0766_;
  wire _0767_;
  wire _0768_;
  wire _0769_;
  wire _0770_;
  wire _0771_;
  wire _0772_;
  wire [7:0] _0773_;
  wire [7:0] _0774_;
  wire _0775_;
  wire _0776_;
  wire _0777_;
  wire _0778_;
  wire _0779_;
  wire _0780_;
  wire _0781_;
  wire _0782_;
  wire _0783_;
  wire _0784_;
  wire _0785_;
  wire _0786_;
  wire _0787_;
  wire _0788_;
  wire _0789_;
  wire _0790_;
  wire _0791_;
  wire _0792_;
  wire _0793_;
  wire _0794_;
  wire _0795_;
  wire _0796_;
  wire _0797_;
  wire _0798_;
  wire _0799_;
  wire _0800_;
  wire _0801_;
  wire _0802_;
  wire _0803_;
  wire _0804_;
  wire _0805_;
  wire _0806_;
  wire _0807_;
  wire _0808_;
  wire _0809_;
  wire _0810_;
  wire _0811_;
  wire _0812_;
  wire _0813_;
  wire _0814_;
  wire _0815_;
  wire _0816_;
  wire _0817_;
  wire _0818_;
  wire _0819_;
  wire _0820_;
  wire _0821_;
  wire _0822_;
  wire _0823_;
  wire _0824_;
  wire _0825_;
  wire _0826_;
  wire _0827_;
  wire _0828_;
  wire _0829_;
  wire _0830_;
  wire _0831_;
  wire _0832_;
  wire _0833_;
  wire _0834_;
  wire _0835_;
  wire _0836_;
  wire _0837_;
  wire _0838_;
  wire _0839_;
  wire _0840_;
  wire _0841_;
  wire _0842_;
  wire _0843_;
  wire _0844_;
  wire _0845_;
  wire _0846_;
  wire _0847_;
  wire _0848_;
  wire _0849_;
  wire _0850_;
  wire _0851_;
  wire _0852_;
  wire _0853_;
  wire _0854_;
  wire _0855_;
  wire _0856_;
  wire _0857_;
  wire _0858_;
  wire _0859_;
  wire _0860_;
  wire _0861_;
  wire _0862_;
  wire _0863_;
  wire _0864_;
  wire _0865_;
  wire _0866_;
  wire _0867_;
  wire _0868_;
  wire _0869_;
  wire _0870_;
  wire _0871_;
  wire _0872_;
  wire _0873_;
  wire _0874_;
  wire _0875_;
  wire _0876_;
  wire _0877_;
  wire _0878_;
  wire _0879_;
  wire _0880_;
  wire _0881_;
  wire _0882_;
  wire _0883_;
  wire _0884_;
  wire _0885_;
  wire _0886_;
  wire _0887_;
  wire _0888_;
  wire _0889_;
  wire _0890_;
  wire _0891_;
  wire _0892_;
  wire _0893_;
  wire _0894_;
  wire _0895_;
  wire _0896_;
  wire _0897_;
  wire _0898_;
  wire _0899_;
  wire _0900_;
  wire _0901_;
  wire _0902_;
  wire _0903_;
  wire _0904_;
  wire _0905_;
  wire _0906_;
  wire _0907_;
  wire _0908_;
  wire _0909_;
  wire _0910_;
  wire _0911_;
  wire _0912_;
  wire _0913_;
  wire _0914_;
  wire _0915_;
  wire _0916_;
  wire _0917_;
  wire _0918_;
  wire _0919_;
  wire _0920_;
  wire _0921_;
  wire _0922_;
  wire _0923_;
  wire _0924_;
  wire _0925_;
  wire _0926_;
  wire _0927_;
  wire _0928_;
  wire _0929_;
  wire _0930_;
  wire _0931_;
  wire _0932_;
  wire _0933_;
  wire _0934_;
  wire _0935_;
  wire _0936_;
  wire _0937_;
  wire _0938_;
  wire _0939_;
  wire _0940_;
  wire _0941_;
  wire _0942_;
  wire _0943_;
  wire _0944_;
  wire _0945_;
  wire _0946_;
  wire _0947_;
  wire _0948_;
  wire _0949_;
  wire _0950_;
  wire _0951_;
  wire _0952_;
  wire _0953_;
  wire _0954_;
  wire _0955_;
  wire _0956_;
  wire _0957_;
  wire _0958_;
  wire _0959_;
  wire _0960_;
  wire _0961_;
  wire _0962_;
  wire _0963_;
  wire _0964_;
  wire _0965_;
  wire _0966_;
  wire _0967_;
  wire _0968_;
  wire _0969_;
  wire _0970_;
  wire _0971_;
  wire _0972_;
  wire _0973_;
  wire _0974_;
  wire _0975_;
  wire _0976_;
  wire _0977_;
  wire _0978_;
  wire _0979_;
  wire _0980_;
  wire _0981_;
  wire _0982_;
  wire _0983_;
  wire _0984_;
  wire _0985_;
  wire _0986_;
  wire _0987_;
  wire _0988_;
  wire _0989_;
  wire _0990_;
  wire _0991_;
  wire _0992_;
  wire _0993_;
  wire _0994_;
  wire _0995_;
  wire _0996_;
  wire _0997_;
  wire _0998_;
  wire _0999_;
  wire _1000_;
  wire _1001_;
  wire _1002_;
  wire _1003_;
  wire _1004_;
  wire _1005_;
  wire _1006_;
  wire _1007_;
  wire _1008_;
  wire _1009_;
  wire _1010_;
  wire _1011_;
  wire _1012_;
  wire _1013_;
  wire _1014_;
  wire _1015_;
  wire _1016_;
  wire _1017_;
  wire _1018_;
  wire _1019_;
  wire _1020_;
  wire _1021_;
  wire _1022_;
  wire _1023_;
  wire _1024_;
  wire _1025_;
  wire _1026_;
  wire _1027_;
  wire _1028_;
  wire _1029_;
  wire _1030_;
  wire [7:0] _1031_;
  wire [7:0] _1032_;
  wire _1033_;
  wire _1034_;
  wire _1035_;
  wire _1036_;
  wire _1037_;
  wire _1038_;
  wire _1039_;
  wire _1040_;
  wire _1041_;
  wire _1042_;
  wire _1043_;
  wire _1044_;
  wire _1045_;
  wire _1046_;
  wire _1047_;
  wire _1048_;
  wire _1049_;
  wire _1050_;
  wire _1051_;
  wire _1052_;
  wire _1053_;
  wire _1054_;
  wire _1055_;
  wire _1056_;
  wire _1057_;
  wire _1058_;
  wire _1059_;
  wire _1060_;
  wire _1061_;
  wire _1062_;
  wire _1063_;
  wire _1064_;
  wire _1065_;
  wire _1066_;
  wire _1067_;
  wire _1068_;
  wire _1069_;
  wire _1070_;
  wire _1071_;
  wire _1072_;
  wire _1073_;
  wire _1074_;
  wire _1075_;
  wire _1076_;
  wire _1077_;
  wire _1078_;
  wire _1079_;
  wire _1080_;
  wire _1081_;
  wire _1082_;
  wire _1083_;
  wire _1084_;
  wire _1085_;
  wire _1086_;
  wire _1087_;
  wire _1088_;
  wire _1089_;
  wire _1090_;
  wire _1091_;
  wire _1092_;
  wire _1093_;
  wire _1094_;
  wire _1095_;
  wire _1096_;
  wire _1097_;
  wire _1098_;
  wire _1099_;
  wire _1100_;
  wire _1101_;
  wire _1102_;
  wire _1103_;
  wire _1104_;
  wire _1105_;
  wire _1106_;
  wire _1107_;
  wire _1108_;
  wire _1109_;
  wire _1110_;
  wire _1111_;
  wire _1112_;
  wire _1113_;
  wire _1114_;
  wire _1115_;
  wire _1116_;
  wire _1117_;
  wire _1118_;
  wire _1119_;
  wire _1120_;
  wire _1121_;
  wire _1122_;
  wire _1123_;
  wire _1124_;
  wire _1125_;
  wire _1126_;
  wire _1127_;
  wire _1128_;
  wire _1129_;
  wire _1130_;
  wire _1131_;
  wire _1132_;
  wire _1133_;
  wire _1134_;
  wire _1135_;
  wire _1136_;
  wire _1137_;
  wire _1138_;
  wire _1139_;
  wire _1140_;
  wire _1141_;
  wire _1142_;
  wire _1143_;
  wire _1144_;
  wire _1145_;
  wire _1146_;
  wire _1147_;
  wire _1148_;
  wire _1149_;
  wire _1150_;
  wire _1151_;
  wire _1152_;
  wire _1153_;
  wire _1154_;
  wire _1155_;
  wire _1156_;
  wire _1157_;
  wire _1158_;
  wire _1159_;
  wire _1160_;
  wire _1161_;
  wire _1162_;
  wire _1163_;
  wire _1164_;
  wire _1165_;
  wire _1166_;
  wire _1167_;
  wire _1168_;
  wire _1169_;
  wire _1170_;
  wire _1171_;
  wire _1172_;
  wire _1173_;
  wire _1174_;
  wire _1175_;
  wire _1176_;
  wire _1177_;
  wire _1178_;
  wire _1179_;
  wire _1180_;
  wire _1181_;
  wire _1182_;
  wire _1183_;
  wire _1184_;
  wire _1185_;
  wire _1186_;
  wire _1187_;
  wire _1188_;
  wire _1189_;
  wire _1190_;
  wire _1191_;
  wire _1192_;
  wire _1193_;
  wire _1194_;
  wire _1195_;
  wire _1196_;
  wire _1197_;
  wire _1198_;
  wire _1199_;
  wire _1200_;
  wire _1201_;
  wire _1202_;
  wire _1203_;
  wire _1204_;
  wire _1205_;
  wire _1206_;
  wire _1207_;
  wire _1208_;
  wire _1209_;
  wire _1210_;
  wire _1211_;
  wire _1212_;
  wire _1213_;
  wire _1214_;
  wire _1215_;
  wire _1216_;
  wire _1217_;
  wire _1218_;
  wire _1219_;
  wire _1220_;
  wire _1221_;
  wire _1222_;
  wire _1223_;
  wire _1224_;
  wire _1225_;
  wire _1226_;
  wire _1227_;
  wire _1228_;
  wire _1229_;
  wire _1230_;
  wire _1231_;
  wire _1232_;
  wire _1233_;
  wire _1234_;
  wire _1235_;
  wire _1236_;
  wire _1237_;
  wire _1238_;
  wire _1239_;
  wire _1240_;
  wire _1241_;
  wire _1242_;
  wire _1243_;
  wire _1244_;
  wire _1245_;
  wire _1246_;
  wire _1247_;
  wire _1248_;
  wire _1249_;
  wire _1250_;
  wire _1251_;
  wire _1252_;
  wire _1253_;
  wire _1254_;
  wire _1255_;
  wire _1256_;
  wire _1257_;
  wire _1258_;
  wire _1259_;
  wire _1260_;
  wire _1261_;
  wire _1262_;
  wire _1263_;
  wire _1264_;
  wire _1265_;
  wire _1266_;
  wire _1267_;
  wire _1268_;
  wire _1269_;
  wire _1270_;
  wire _1271_;
  wire _1272_;
  wire _1273_;
  wire _1274_;
  wire _1275_;
  wire _1276_;
  wire _1277_;
  wire _1278_;
  wire _1279_;
  wire _1280_;
  wire _1281_;
  wire _1282_;
  wire _1283_;
  wire _1284_;
  wire _1285_;
  wire _1286_;
  wire _1287_;
  wire _1288_;
  wire [7:0] _1289_;
  wire [7:0] _1290_;
  wire _1291_;
  wire _1292_;
  wire _1293_;
  wire _1294_;
  wire _1295_;
  wire _1296_;
  wire _1297_;
  wire _1298_;
  wire _1299_;
  wire _1300_;
  wire _1301_;
  wire _1302_;
  wire _1303_;
  wire _1304_;
  wire _1305_;
  wire _1306_;
  wire _1307_;
  wire _1308_;
  wire _1309_;
  wire _1310_;
  wire _1311_;
  wire _1312_;
  wire _1313_;
  wire _1314_;
  wire _1315_;
  wire _1316_;
  wire _1317_;
  wire _1318_;
  wire _1319_;
  wire _1320_;
  wire _1321_;
  wire _1322_;
  wire _1323_;
  wire _1324_;
  wire _1325_;
  wire _1326_;
  wire _1327_;
  wire _1328_;
  wire _1329_;
  wire _1330_;
  wire _1331_;
  wire _1332_;
  wire _1333_;
  wire _1334_;
  wire _1335_;
  wire _1336_;
  wire _1337_;
  wire _1338_;
  wire _1339_;
  wire _1340_;
  wire _1341_;
  wire _1342_;
  wire _1343_;
  wire _1344_;
  wire _1345_;
  wire _1346_;
  wire _1347_;
  wire _1348_;
  wire _1349_;
  wire _1350_;
  wire _1351_;
  wire _1352_;
  wire _1353_;
  wire _1354_;
  wire _1355_;
  wire _1356_;
  wire _1357_;
  wire _1358_;
  wire _1359_;
  wire _1360_;
  wire _1361_;
  wire _1362_;
  wire _1363_;
  wire _1364_;
  wire _1365_;
  wire _1366_;
  wire _1367_;
  wire _1368_;
  wire _1369_;
  wire _1370_;
  wire _1371_;
  wire _1372_;
  wire _1373_;
  wire _1374_;
  wire _1375_;
  wire _1376_;
  wire _1377_;
  wire _1378_;
  wire _1379_;
  wire _1380_;
  wire _1381_;
  wire _1382_;
  wire _1383_;
  wire _1384_;
  wire _1385_;
  wire _1386_;
  wire _1387_;
  wire _1388_;
  wire _1389_;
  wire _1390_;
  wire _1391_;
  wire _1392_;
  wire _1393_;
  wire _1394_;
  wire _1395_;
  wire _1396_;
  wire _1397_;
  wire _1398_;
  wire _1399_;
  wire _1400_;
  wire _1401_;
  wire _1402_;
  wire _1403_;
  wire _1404_;
  wire _1405_;
  wire _1406_;
  wire _1407_;
  wire _1408_;
  wire _1409_;
  wire _1410_;
  wire _1411_;
  wire _1412_;
  wire _1413_;
  wire _1414_;
  wire _1415_;
  wire _1416_;
  wire _1417_;
  wire _1418_;
  wire _1419_;
  wire _1420_;
  wire _1421_;
  wire _1422_;
  wire _1423_;
  wire _1424_;
  wire _1425_;
  wire _1426_;
  wire _1427_;
  wire _1428_;
  wire _1429_;
  wire _1430_;
  wire _1431_;
  wire _1432_;
  wire _1433_;
  wire _1434_;
  wire _1435_;
  wire _1436_;
  wire _1437_;
  wire _1438_;
  wire _1439_;
  wire _1440_;
  wire _1441_;
  wire _1442_;
  wire _1443_;
  wire _1444_;
  wire _1445_;
  wire _1446_;
  wire _1447_;
  wire _1448_;
  wire _1449_;
  wire _1450_;
  wire _1451_;
  wire _1452_;
  wire _1453_;
  wire _1454_;
  wire _1455_;
  wire _1456_;
  wire _1457_;
  wire _1458_;
  wire _1459_;
  wire _1460_;
  wire _1461_;
  wire _1462_;
  wire _1463_;
  wire _1464_;
  wire _1465_;
  wire _1466_;
  wire _1467_;
  wire _1468_;
  wire _1469_;
  wire _1470_;
  wire _1471_;
  wire _1472_;
  wire _1473_;
  wire _1474_;
  wire _1475_;
  wire _1476_;
  wire _1477_;
  wire _1478_;
  wire _1479_;
  wire _1480_;
  wire _1481_;
  wire _1482_;
  wire _1483_;
  wire _1484_;
  wire _1485_;
  wire _1486_;
  wire _1487_;
  wire _1488_;
  wire _1489_;
  wire _1490_;
  wire _1491_;
  wire _1492_;
  wire _1493_;
  wire _1494_;
  wire _1495_;
  wire _1496_;
  wire _1497_;
  wire _1498_;
  wire _1499_;
  wire _1500_;
  wire _1501_;
  wire _1502_;
  wire _1503_;
  wire _1504_;
  wire _1505_;
  wire _1506_;
  wire _1507_;
  wire _1508_;
  wire _1509_;
  wire _1510_;
  wire _1511_;
  wire _1512_;
  wire _1513_;
  wire _1514_;
  wire _1515_;
  wire _1516_;
  wire _1517_;
  wire _1518_;
  wire _1519_;
  wire _1520_;
  wire _1521_;
  wire _1522_;
  wire _1523_;
  wire _1524_;
  wire _1525_;
  wire _1526_;
  wire _1527_;
  wire _1528_;
  wire _1529_;
  wire _1530_;
  wire _1531_;
  wire _1532_;
  wire _1533_;
  wire _1534_;
  wire _1535_;
  wire _1536_;
  wire _1537_;
  wire _1538_;
  wire _1539_;
  wire _1540_;
  wire _1541_;
  wire _1542_;
  wire _1543_;
  wire _1544_;
  wire _1545_;
  wire _1546_;
  wire [7:0] _1547_;
  wire [7:0] _1548_;
  wire _1549_;
  wire _1550_;
  wire _1551_;
  wire _1552_;
  wire _1553_;
  wire _1554_;
  wire _1555_;
  wire _1556_;
  wire _1557_;
  wire _1558_;
  wire _1559_;
  wire _1560_;
  wire _1561_;
  wire _1562_;
  wire _1563_;
  wire _1564_;
  wire _1565_;
  wire _1566_;
  wire _1567_;
  wire _1568_;
  wire _1569_;
  wire _1570_;
  wire _1571_;
  wire _1572_;
  wire _1573_;
  wire _1574_;
  wire _1575_;
  wire _1576_;
  wire _1577_;
  wire _1578_;
  wire _1579_;
  wire _1580_;
  wire _1581_;
  wire _1582_;
  wire _1583_;
  wire _1584_;
  wire _1585_;
  wire _1586_;
  wire _1587_;
  wire _1588_;
  wire _1589_;
  wire _1590_;
  wire _1591_;
  wire _1592_;
  wire _1593_;
  wire _1594_;
  wire _1595_;
  wire _1596_;
  wire _1597_;
  wire _1598_;
  wire _1599_;
  wire _1600_;
  wire _1601_;
  wire _1602_;
  wire _1603_;
  wire _1604_;
  wire _1605_;
  wire _1606_;
  wire _1607_;
  wire _1608_;
  wire _1609_;
  wire _1610_;
  wire _1611_;
  wire _1612_;
  wire _1613_;
  wire _1614_;
  wire _1615_;
  wire _1616_;
  wire _1617_;
  wire _1618_;
  wire _1619_;
  wire _1620_;
  wire _1621_;
  wire _1622_;
  wire _1623_;
  wire _1624_;
  wire _1625_;
  wire _1626_;
  wire _1627_;
  wire _1628_;
  wire _1629_;
  wire _1630_;
  wire _1631_;
  wire _1632_;
  wire _1633_;
  wire _1634_;
  wire _1635_;
  wire _1636_;
  wire _1637_;
  wire _1638_;
  wire _1639_;
  wire _1640_;
  wire _1641_;
  wire _1642_;
  wire _1643_;
  wire _1644_;
  wire _1645_;
  wire _1646_;
  wire _1647_;
  wire _1648_;
  wire _1649_;
  wire _1650_;
  wire _1651_;
  wire _1652_;
  wire _1653_;
  wire _1654_;
  wire _1655_;
  wire _1656_;
  wire _1657_;
  wire _1658_;
  wire _1659_;
  wire _1660_;
  wire _1661_;
  wire _1662_;
  wire _1663_;
  wire _1664_;
  wire _1665_;
  wire _1666_;
  wire _1667_;
  wire _1668_;
  wire _1669_;
  wire _1670_;
  wire _1671_;
  wire _1672_;
  wire _1673_;
  wire _1674_;
  wire _1675_;
  wire _1676_;
  wire _1677_;
  wire _1678_;
  wire _1679_;
  wire _1680_;
  wire _1681_;
  wire _1682_;
  wire _1683_;
  wire _1684_;
  wire _1685_;
  wire _1686_;
  wire _1687_;
  wire _1688_;
  wire _1689_;
  wire _1690_;
  wire _1691_;
  wire _1692_;
  wire _1693_;
  wire _1694_;
  wire _1695_;
  wire _1696_;
  wire _1697_;
  wire _1698_;
  wire _1699_;
  wire _1700_;
  wire _1701_;
  wire _1702_;
  wire _1703_;
  wire _1704_;
  wire _1705_;
  wire _1706_;
  wire _1707_;
  wire _1708_;
  wire _1709_;
  wire _1710_;
  wire _1711_;
  wire _1712_;
  wire _1713_;
  wire _1714_;
  wire _1715_;
  wire _1716_;
  wire _1717_;
  wire _1718_;
  wire _1719_;
  wire _1720_;
  wire _1721_;
  wire _1722_;
  wire _1723_;
  wire _1724_;
  wire _1725_;
  wire _1726_;
  wire _1727_;
  wire _1728_;
  wire _1729_;
  wire _1730_;
  wire _1731_;
  wire _1732_;
  wire _1733_;
  wire _1734_;
  wire _1735_;
  wire _1736_;
  wire _1737_;
  wire _1738_;
  wire _1739_;
  wire _1740_;
  wire _1741_;
  wire _1742_;
  wire _1743_;
  wire _1744_;
  wire _1745_;
  wire _1746_;
  wire _1747_;
  wire _1748_;
  wire _1749_;
  wire _1750_;
  wire _1751_;
  wire _1752_;
  wire _1753_;
  wire _1754_;
  wire _1755_;
  wire _1756_;
  wire _1757_;
  wire _1758_;
  wire _1759_;
  wire _1760_;
  wire _1761_;
  wire _1762_;
  wire _1763_;
  wire _1764_;
  wire _1765_;
  wire _1766_;
  wire _1767_;
  wire _1768_;
  wire _1769_;
  wire _1770_;
  wire _1771_;
  wire _1772_;
  wire _1773_;
  wire _1774_;
  wire _1775_;
  wire _1776_;
  wire _1777_;
  wire _1778_;
  wire _1779_;
  wire _1780_;
  wire _1781_;
  wire _1782_;
  wire _1783_;
  wire _1784_;
  wire _1785_;
  wire _1786_;
  wire _1787_;
  wire _1788_;
  wire _1789_;
  wire _1790_;
  wire _1791_;
  wire _1792_;
  wire _1793_;
  wire _1794_;
  wire _1795_;
  wire _1796_;
  wire _1797_;
  wire _1798_;
  wire _1799_;
  wire _1800_;
  wire _1801_;
  wire _1802_;
  wire _1803_;
  wire _1804_;
  wire [7:0] _1805_;
  wire [7:0] _1806_;
  wire _1807_;
  wire _1808_;
  wire _1809_;
  wire _1810_;
  wire _1811_;
  wire _1812_;
  wire _1813_;
  wire _1814_;
  wire _1815_;
  wire _1816_;
  wire _1817_;
  wire _1818_;
  wire _1819_;
  wire _1820_;
  wire _1821_;
  wire _1822_;
  wire _1823_;
  wire _1824_;
  wire _1825_;
  wire _1826_;
  wire _1827_;
  wire _1828_;
  wire _1829_;
  wire _1830_;
  wire _1831_;
  wire _1832_;
  wire _1833_;
  wire _1834_;
  wire _1835_;
  wire _1836_;
  wire _1837_;
  wire _1838_;
  wire _1839_;
  wire _1840_;
  wire _1841_;
  wire _1842_;
  wire _1843_;
  wire _1844_;
  wire _1845_;
  wire _1846_;
  wire _1847_;
  wire _1848_;
  wire _1849_;
  wire _1850_;
  wire _1851_;
  wire _1852_;
  wire _1853_;
  wire _1854_;
  wire _1855_;
  wire _1856_;
  wire _1857_;
  wire _1858_;
  wire _1859_;
  wire _1860_;
  wire _1861_;
  wire _1862_;
  wire _1863_;
  wire _1864_;
  wire _1865_;
  wire _1866_;
  wire _1867_;
  wire _1868_;
  wire _1869_;
  wire _1870_;
  wire _1871_;
  wire _1872_;
  wire _1873_;
  wire _1874_;
  wire _1875_;
  wire _1876_;
  wire _1877_;
  wire _1878_;
  wire _1879_;
  wire _1880_;
  wire _1881_;
  wire _1882_;
  wire _1883_;
  wire _1884_;
  wire _1885_;
  wire _1886_;
  wire _1887_;
  wire _1888_;
  wire _1889_;
  wire _1890_;
  wire _1891_;
  wire _1892_;
  wire _1893_;
  wire _1894_;
  wire _1895_;
  wire _1896_;
  wire _1897_;
  wire _1898_;
  wire _1899_;
  wire _1900_;
  wire _1901_;
  wire _1902_;
  wire _1903_;
  wire _1904_;
  wire _1905_;
  wire _1906_;
  wire _1907_;
  wire _1908_;
  wire _1909_;
  wire _1910_;
  wire _1911_;
  wire _1912_;
  wire _1913_;
  wire _1914_;
  wire _1915_;
  wire _1916_;
  wire _1917_;
  wire _1918_;
  wire _1919_;
  wire _1920_;
  wire _1921_;
  wire _1922_;
  wire _1923_;
  wire _1924_;
  wire _1925_;
  wire _1926_;
  wire _1927_;
  wire _1928_;
  wire _1929_;
  wire _1930_;
  wire _1931_;
  wire _1932_;
  wire _1933_;
  wire _1934_;
  wire _1935_;
  wire _1936_;
  wire _1937_;
  wire _1938_;
  wire _1939_;
  wire _1940_;
  wire _1941_;
  wire _1942_;
  wire _1943_;
  wire _1944_;
  wire _1945_;
  wire _1946_;
  wire _1947_;
  wire _1948_;
  wire _1949_;
  wire _1950_;
  wire _1951_;
  wire _1952_;
  wire _1953_;
  wire _1954_;
  wire _1955_;
  wire _1956_;
  wire _1957_;
  wire _1958_;
  wire _1959_;
  wire _1960_;
  wire _1961_;
  wire _1962_;
  wire _1963_;
  wire _1964_;
  wire _1965_;
  wire _1966_;
  wire _1967_;
  wire _1968_;
  wire _1969_;
  wire _1970_;
  wire _1971_;
  wire _1972_;
  wire _1973_;
  wire _1974_;
  wire _1975_;
  wire _1976_;
  wire _1977_;
  wire _1978_;
  wire _1979_;
  wire _1980_;
  wire _1981_;
  wire _1982_;
  wire _1983_;
  wire _1984_;
  wire _1985_;
  wire _1986_;
  wire _1987_;
  wire _1988_;
  wire _1989_;
  wire _1990_;
  wire _1991_;
  wire _1992_;
  wire _1993_;
  wire _1994_;
  wire _1995_;
  wire _1996_;
  wire _1997_;
  wire _1998_;
  wire _1999_;
  wire _2000_;
  wire _2001_;
  wire _2002_;
  wire _2003_;
  wire _2004_;
  wire _2005_;
  wire _2006_;
  wire _2007_;
  wire _2008_;
  wire _2009_;
  wire _2010_;
  wire _2011_;
  wire _2012_;
  wire _2013_;
  wire _2014_;
  wire _2015_;
  wire _2016_;
  wire _2017_;
  wire _2018_;
  wire _2019_;
  wire _2020_;
  wire _2021_;
  wire _2022_;
  wire _2023_;
  wire _2024_;
  wire _2025_;
  wire _2026_;
  wire _2027_;
  wire _2028_;
  wire _2029_;
  wire _2030_;
  wire _2031_;
  wire _2032_;
  wire _2033_;
  wire _2034_;
  wire _2035_;
  wire _2036_;
  wire _2037_;
  wire _2038_;
  wire _2039_;
  wire _2040_;
  wire _2041_;
  wire _2042_;
  wire _2043_;
  wire _2044_;
  wire _2045_;
  wire _2046_;
  wire _2047_;
  wire _2048_;
  wire _2049_;
  wire _2050_;
  wire _2051_;
  wire _2052_;
  wire _2053_;
  wire _2054_;
  wire _2055_;
  wire _2056_;
  wire _2057_;
  wire _2058_;
  wire _2059_;
  wire _2060_;
  wire _2061_;
  wire _2062_;
  wire [7:0] _2063_;
  wire [7:0] _2064_;
  wire _2065_;
  wire _2066_;
  wire _2067_;
  wire _2068_;
  wire _2069_;
  wire _2070_;
  wire _2071_;
  wire _2072_;
  wire _2073_;
  wire _2074_;
  wire _2075_;
  wire _2076_;
  wire _2077_;
  wire _2078_;
  wire _2079_;
  wire _2080_;
  wire _2081_;
  wire _2082_;
  wire _2083_;
  wire _2084_;
  wire _2085_;
  wire _2086_;
  wire _2087_;
  wire _2088_;
  wire _2089_;
  wire _2090_;
  wire _2091_;
  wire _2092_;
  wire _2093_;
  wire _2094_;
  wire _2095_;
  wire _2096_;
  wire _2097_;
  wire _2098_;
  wire _2099_;
  wire _2100_;
  wire _2101_;
  wire _2102_;
  wire _2103_;
  wire _2104_;
  wire _2105_;
  wire _2106_;
  wire _2107_;
  wire _2108_;
  wire _2109_;
  wire _2110_;
  wire _2111_;
  wire _2112_;
  wire _2113_;
  wire _2114_;
  wire _2115_;
  wire _2116_;
  wire _2117_;
  wire _2118_;
  wire _2119_;
  wire _2120_;
  wire _2121_;
  wire _2122_;
  wire _2123_;
  wire _2124_;
  wire _2125_;
  wire _2126_;
  wire _2127_;
  wire _2128_;
  wire _2129_;
  wire _2130_;
  wire _2131_;
  wire _2132_;
  wire _2133_;
  wire _2134_;
  wire _2135_;
  wire _2136_;
  wire _2137_;
  wire _2138_;
  wire _2139_;
  wire _2140_;
  wire _2141_;
  wire _2142_;
  wire _2143_;
  wire _2144_;
  wire _2145_;
  wire _2146_;
  wire _2147_;
  wire _2148_;
  wire _2149_;
  wire _2150_;
  wire _2151_;
  wire _2152_;
  wire _2153_;
  wire _2154_;
  wire _2155_;
  wire _2156_;
  wire _2157_;
  wire _2158_;
  wire _2159_;
  wire _2160_;
  wire _2161_;
  wire _2162_;
  wire _2163_;
  wire _2164_;
  wire _2165_;
  wire _2166_;
  wire _2167_;
  wire _2168_;
  wire _2169_;
  wire _2170_;
  wire _2171_;
  wire _2172_;
  wire _2173_;
  wire _2174_;
  wire _2175_;
  wire _2176_;
  wire _2177_;
  wire _2178_;
  wire _2179_;
  wire _2180_;
  wire _2181_;
  wire _2182_;
  wire _2183_;
  wire _2184_;
  wire _2185_;
  wire _2186_;
  wire _2187_;
  wire _2188_;
  wire _2189_;
  wire _2190_;
  wire _2191_;
  wire _2192_;
  wire _2193_;
  wire _2194_;
  wire _2195_;
  wire _2196_;
  wire _2197_;
  wire _2198_;
  wire _2199_;
  wire _2200_;
  wire _2201_;
  wire _2202_;
  wire _2203_;
  wire _2204_;
  wire _2205_;
  wire _2206_;
  wire _2207_;
  wire _2208_;
  wire _2209_;
  wire _2210_;
  wire _2211_;
  wire _2212_;
  wire _2213_;
  wire _2214_;
  wire _2215_;
  wire _2216_;
  wire _2217_;
  wire _2218_;
  wire _2219_;
  wire _2220_;
  wire _2221_;
  wire _2222_;
  wire _2223_;
  wire _2224_;
  wire _2225_;
  wire _2226_;
  wire _2227_;
  wire _2228_;
  wire _2229_;
  wire _2230_;
  wire _2231_;
  wire _2232_;
  wire _2233_;
  wire _2234_;
  wire _2235_;
  wire _2236_;
  wire _2237_;
  wire _2238_;
  wire _2239_;
  wire _2240_;
  wire _2241_;
  wire _2242_;
  wire _2243_;
  wire _2244_;
  wire _2245_;
  wire _2246_;
  wire _2247_;
  wire _2248_;
  wire _2249_;
  wire _2250_;
  wire _2251_;
  wire _2252_;
  wire _2253_;
  wire _2254_;
  wire _2255_;
  wire _2256_;
  wire _2257_;
  wire _2258_;
  wire _2259_;
  wire _2260_;
  wire _2261_;
  wire _2262_;
  wire _2263_;
  wire _2264_;
  wire _2265_;
  wire _2266_;
  wire _2267_;
  wire _2268_;
  wire _2269_;
  wire _2270_;
  wire _2271_;
  wire _2272_;
  wire _2273_;
  wire _2274_;
  wire _2275_;
  wire _2276_;
  wire _2277_;
  wire _2278_;
  wire _2279_;
  wire _2280_;
  wire _2281_;
  wire _2282_;
  wire _2283_;
  wire _2284_;
  wire _2285_;
  wire _2286_;
  wire _2287_;
  wire _2288_;
  wire _2289_;
  wire _2290_;
  wire _2291_;
  wire _2292_;
  wire _2293_;
  wire _2294_;
  wire _2295_;
  wire _2296_;
  wire _2297_;
  wire _2298_;
  wire _2299_;
  wire _2300_;
  wire _2301_;
  wire _2302_;
  wire _2303_;
  wire _2304_;
  wire _2305_;
  wire _2306_;
  wire _2307_;
  wire _2308_;
  wire _2309_;
  wire _2310_;
  wire _2311_;
  wire _2312_;
  wire _2313_;
  wire _2314_;
  wire _2315_;
  wire _2316_;
  wire _2317_;
  wire _2318_;
  wire _2319_;
  wire _2320_;
  wire [7:0] _2321_;
  wire [7:0] _2322_;
  wire _2323_;
  wire _2324_;
  wire _2325_;
  wire _2326_;
  wire _2327_;
  wire _2328_;
  wire _2329_;
  wire _2330_;
  wire _2331_;
  wire _2332_;
  wire _2333_;
  wire _2334_;
  wire _2335_;
  wire _2336_;
  wire _2337_;
  wire _2338_;
  wire _2339_;
  wire _2340_;
  wire _2341_;
  wire _2342_;
  wire _2343_;
  wire _2344_;
  wire _2345_;
  wire _2346_;
  wire _2347_;
  wire _2348_;
  wire _2349_;
  wire _2350_;
  wire _2351_;
  wire _2352_;
  wire _2353_;
  wire _2354_;
  wire _2355_;
  wire _2356_;
  wire _2357_;
  wire _2358_;
  wire _2359_;
  wire _2360_;
  wire _2361_;
  wire _2362_;
  wire _2363_;
  wire _2364_;
  wire _2365_;
  wire _2366_;
  wire _2367_;
  wire _2368_;
  wire _2369_;
  wire _2370_;
  wire _2371_;
  wire _2372_;
  wire _2373_;
  wire _2374_;
  wire _2375_;
  wire _2376_;
  wire _2377_;
  wire _2378_;
  wire _2379_;
  wire _2380_;
  wire _2381_;
  wire _2382_;
  wire _2383_;
  wire _2384_;
  wire _2385_;
  wire _2386_;
  wire _2387_;
  wire _2388_;
  wire _2389_;
  wire _2390_;
  wire _2391_;
  wire _2392_;
  wire _2393_;
  wire _2394_;
  wire _2395_;
  wire _2396_;
  wire _2397_;
  wire _2398_;
  wire _2399_;
  wire _2400_;
  wire _2401_;
  wire _2402_;
  wire _2403_;
  wire _2404_;
  wire _2405_;
  wire _2406_;
  wire _2407_;
  wire _2408_;
  wire _2409_;
  wire _2410_;
  wire _2411_;
  wire _2412_;
  wire _2413_;
  wire _2414_;
  wire _2415_;
  wire _2416_;
  wire _2417_;
  wire _2418_;
  wire _2419_;
  wire _2420_;
  wire _2421_;
  wire _2422_;
  wire _2423_;
  wire _2424_;
  wire _2425_;
  wire _2426_;
  wire _2427_;
  wire _2428_;
  wire _2429_;
  wire _2430_;
  wire _2431_;
  wire _2432_;
  wire _2433_;
  wire _2434_;
  wire _2435_;
  wire _2436_;
  wire _2437_;
  wire _2438_;
  wire _2439_;
  wire _2440_;
  wire _2441_;
  wire _2442_;
  wire _2443_;
  wire _2444_;
  wire _2445_;
  wire _2446_;
  wire _2447_;
  wire _2448_;
  wire _2449_;
  wire _2450_;
  wire _2451_;
  wire _2452_;
  wire _2453_;
  wire _2454_;
  wire _2455_;
  wire _2456_;
  wire _2457_;
  wire _2458_;
  wire _2459_;
  wire _2460_;
  wire _2461_;
  wire _2462_;
  wire _2463_;
  wire _2464_;
  wire _2465_;
  wire _2466_;
  wire _2467_;
  wire _2468_;
  wire _2469_;
  wire _2470_;
  wire _2471_;
  wire _2472_;
  wire _2473_;
  wire _2474_;
  wire _2475_;
  wire _2476_;
  wire _2477_;
  wire _2478_;
  wire _2479_;
  wire _2480_;
  wire _2481_;
  wire _2482_;
  wire _2483_;
  wire _2484_;
  wire _2485_;
  wire _2486_;
  wire _2487_;
  wire _2488_;
  wire _2489_;
  wire _2490_;
  wire _2491_;
  wire _2492_;
  wire _2493_;
  wire _2494_;
  wire _2495_;
  wire _2496_;
  wire _2497_;
  wire _2498_;
  wire _2499_;
  wire _2500_;
  wire _2501_;
  wire _2502_;
  wire _2503_;
  wire _2504_;
  wire _2505_;
  wire _2506_;
  wire _2507_;
  wire _2508_;
  wire _2509_;
  wire _2510_;
  wire _2511_;
  wire _2512_;
  wire _2513_;
  wire _2514_;
  wire _2515_;
  wire _2516_;
  wire _2517_;
  wire _2518_;
  wire _2519_;
  wire _2520_;
  wire _2521_;
  wire _2522_;
  wire _2523_;
  wire _2524_;
  wire _2525_;
  wire _2526_;
  wire _2527_;
  wire _2528_;
  wire _2529_;
  wire _2530_;
  wire _2531_;
  wire _2532_;
  wire _2533_;
  wire _2534_;
  wire _2535_;
  wire _2536_;
  wire _2537_;
  wire _2538_;
  wire _2539_;
  wire _2540_;
  wire _2541_;
  wire _2542_;
  wire _2543_;
  wire _2544_;
  wire _2545_;
  wire _2546_;
  wire _2547_;
  wire _2548_;
  wire _2549_;
  wire _2550_;
  wire _2551_;
  wire _2552_;
  wire _2553_;
  wire _2554_;
  wire _2555_;
  wire _2556_;
  wire _2557_;
  wire _2558_;
  wire _2559_;
  wire _2560_;
  wire _2561_;
  wire _2562_;
  wire _2563_;
  wire _2564_;
  wire _2565_;
  wire _2566_;
  wire _2567_;
  wire _2568_;
  wire _2569_;
  wire _2570_;
  wire _2571_;
  wire _2572_;
  wire _2573_;
  wire _2574_;
  wire _2575_;
  wire _2576_;
  wire _2577_;
  wire _2578_;
  wire [7:0] _2579_;
  wire [7:0] _2580_;
  wire _2581_;
  wire _2582_;
  wire _2583_;
  wire _2584_;
  wire _2585_;
  wire _2586_;
  wire _2587_;
  wire _2588_;
  wire _2589_;
  wire _2590_;
  wire _2591_;
  wire _2592_;
  wire _2593_;
  wire _2594_;
  wire _2595_;
  wire _2596_;
  wire _2597_;
  wire _2598_;
  wire _2599_;
  wire _2600_;
  wire _2601_;
  wire _2602_;
  wire _2603_;
  wire _2604_;
  wire _2605_;
  wire _2606_;
  wire _2607_;
  wire _2608_;
  wire _2609_;
  wire _2610_;
  wire _2611_;
  wire _2612_;
  wire _2613_;
  wire _2614_;
  wire _2615_;
  wire _2616_;
  wire _2617_;
  wire _2618_;
  wire _2619_;
  wire _2620_;
  wire _2621_;
  wire _2622_;
  wire _2623_;
  wire _2624_;
  wire _2625_;
  wire _2626_;
  wire _2627_;
  wire _2628_;
  wire _2629_;
  wire _2630_;
  wire _2631_;
  wire _2632_;
  wire _2633_;
  wire _2634_;
  wire _2635_;
  wire _2636_;
  wire _2637_;
  wire _2638_;
  wire _2639_;
  wire _2640_;
  wire _2641_;
  wire _2642_;
  wire _2643_;
  wire _2644_;
  wire _2645_;
  wire _2646_;
  wire _2647_;
  wire _2648_;
  wire _2649_;
  wire _2650_;
  wire _2651_;
  wire _2652_;
  wire _2653_;
  wire _2654_;
  wire _2655_;
  wire _2656_;
  wire _2657_;
  wire _2658_;
  wire _2659_;
  wire _2660_;
  wire _2661_;
  wire _2662_;
  wire _2663_;
  wire _2664_;
  wire _2665_;
  wire _2666_;
  wire _2667_;
  wire _2668_;
  wire _2669_;
  wire _2670_;
  wire _2671_;
  wire _2672_;
  wire _2673_;
  wire _2674_;
  wire _2675_;
  wire _2676_;
  wire _2677_;
  wire _2678_;
  wire _2679_;
  wire _2680_;
  wire _2681_;
  wire _2682_;
  wire _2683_;
  wire _2684_;
  wire _2685_;
  wire _2686_;
  wire _2687_;
  wire _2688_;
  wire _2689_;
  wire _2690_;
  wire _2691_;
  wire _2692_;
  wire _2693_;
  wire _2694_;
  wire _2695_;
  wire _2696_;
  wire _2697_;
  wire _2698_;
  wire _2699_;
  wire _2700_;
  wire _2701_;
  wire _2702_;
  wire _2703_;
  wire _2704_;
  wire _2705_;
  wire _2706_;
  wire _2707_;
  wire _2708_;
  wire _2709_;
  wire _2710_;
  wire _2711_;
  wire _2712_;
  wire _2713_;
  wire _2714_;
  wire _2715_;
  wire _2716_;
  wire _2717_;
  wire _2718_;
  wire _2719_;
  wire _2720_;
  wire _2721_;
  wire _2722_;
  wire _2723_;
  wire _2724_;
  wire _2725_;
  wire _2726_;
  wire _2727_;
  wire _2728_;
  wire _2729_;
  wire _2730_;
  wire _2731_;
  wire _2732_;
  wire _2733_;
  wire _2734_;
  wire _2735_;
  wire _2736_;
  wire _2737_;
  wire _2738_;
  wire _2739_;
  wire _2740_;
  wire _2741_;
  wire _2742_;
  wire _2743_;
  wire _2744_;
  wire _2745_;
  wire _2746_;
  wire _2747_;
  wire _2748_;
  wire _2749_;
  wire _2750_;
  wire _2751_;
  wire _2752_;
  wire _2753_;
  wire _2754_;
  wire _2755_;
  wire _2756_;
  wire _2757_;
  wire _2758_;
  wire _2759_;
  wire _2760_;
  wire _2761_;
  wire _2762_;
  wire _2763_;
  wire _2764_;
  wire _2765_;
  wire _2766_;
  wire _2767_;
  wire _2768_;
  wire _2769_;
  wire _2770_;
  wire _2771_;
  wire _2772_;
  wire _2773_;
  wire _2774_;
  wire _2775_;
  wire _2776_;
  wire _2777_;
  wire _2778_;
  wire _2779_;
  wire _2780_;
  wire _2781_;
  wire _2782_;
  wire _2783_;
  wire _2784_;
  wire _2785_;
  wire _2786_;
  wire _2787_;
  wire _2788_;
  wire _2789_;
  wire _2790_;
  wire _2791_;
  wire _2792_;
  wire _2793_;
  wire _2794_;
  wire _2795_;
  wire _2796_;
  wire _2797_;
  wire _2798_;
  wire _2799_;
  wire _2800_;
  wire _2801_;
  wire _2802_;
  wire _2803_;
  wire _2804_;
  wire _2805_;
  wire _2806_;
  wire _2807_;
  wire _2808_;
  wire _2809_;
  wire _2810_;
  wire _2811_;
  wire _2812_;
  wire _2813_;
  wire _2814_;
  wire _2815_;
  wire _2816_;
  wire _2817_;
  wire _2818_;
  wire _2819_;
  wire _2820_;
  wire _2821_;
  wire _2822_;
  wire _2823_;
  wire _2824_;
  wire _2825_;
  wire _2826_;
  wire _2827_;
  wire _2828_;
  wire _2829_;
  wire _2830_;
  wire _2831_;
  wire _2832_;
  wire _2833_;
  wire _2834_;
  wire _2835_;
  wire _2836_;
  wire [7:0] _2837_;
  wire [7:0] _2838_;
  wire _2839_;
  wire _2840_;
  wire _2841_;
  wire _2842_;
  wire _2843_;
  wire _2844_;
  wire _2845_;
  wire _2846_;
  wire _2847_;
  wire _2848_;
  wire _2849_;
  wire _2850_;
  wire _2851_;
  wire _2852_;
  wire _2853_;
  wire _2854_;
  wire _2855_;
  wire _2856_;
  wire _2857_;
  wire _2858_;
  wire _2859_;
  wire _2860_;
  wire _2861_;
  wire _2862_;
  wire _2863_;
  wire _2864_;
  wire _2865_;
  wire _2866_;
  wire _2867_;
  wire _2868_;
  wire _2869_;
  wire _2870_;
  wire _2871_;
  wire _2872_;
  wire _2873_;
  wire _2874_;
  wire _2875_;
  wire _2876_;
  wire _2877_;
  wire _2878_;
  wire _2879_;
  wire _2880_;
  wire _2881_;
  wire _2882_;
  wire _2883_;
  wire _2884_;
  wire _2885_;
  wire _2886_;
  wire _2887_;
  wire _2888_;
  wire _2889_;
  wire _2890_;
  wire _2891_;
  wire _2892_;
  wire _2893_;
  wire _2894_;
  wire _2895_;
  wire _2896_;
  wire _2897_;
  wire _2898_;
  wire _2899_;
  wire _2900_;
  wire _2901_;
  wire _2902_;
  wire _2903_;
  wire _2904_;
  wire _2905_;
  wire _2906_;
  wire _2907_;
  wire _2908_;
  wire _2909_;
  wire _2910_;
  wire _2911_;
  wire _2912_;
  wire _2913_;
  wire _2914_;
  wire _2915_;
  wire _2916_;
  wire _2917_;
  wire _2918_;
  wire _2919_;
  wire _2920_;
  wire _2921_;
  wire _2922_;
  wire _2923_;
  wire _2924_;
  wire _2925_;
  wire _2926_;
  wire _2927_;
  wire _2928_;
  wire _2929_;
  wire _2930_;
  wire _2931_;
  wire _2932_;
  wire _2933_;
  wire _2934_;
  wire _2935_;
  wire _2936_;
  wire _2937_;
  wire _2938_;
  wire _2939_;
  wire _2940_;
  wire _2941_;
  wire _2942_;
  wire _2943_;
  wire _2944_;
  wire _2945_;
  wire _2946_;
  wire _2947_;
  wire _2948_;
  wire _2949_;
  wire _2950_;
  wire _2951_;
  wire _2952_;
  wire _2953_;
  wire _2954_;
  wire _2955_;
  wire _2956_;
  wire _2957_;
  wire _2958_;
  wire _2959_;
  wire _2960_;
  wire _2961_;
  wire _2962_;
  wire _2963_;
  wire _2964_;
  wire _2965_;
  wire _2966_;
  wire _2967_;
  wire _2968_;
  wire _2969_;
  wire _2970_;
  wire _2971_;
  wire _2972_;
  wire _2973_;
  wire _2974_;
  wire _2975_;
  wire _2976_;
  wire _2977_;
  wire _2978_;
  wire _2979_;
  wire _2980_;
  wire _2981_;
  wire _2982_;
  wire _2983_;
  wire _2984_;
  wire _2985_;
  wire _2986_;
  wire _2987_;
  wire _2988_;
  wire _2989_;
  wire _2990_;
  wire _2991_;
  wire _2992_;
  wire _2993_;
  wire _2994_;
  wire _2995_;
  wire _2996_;
  wire _2997_;
  wire _2998_;
  wire _2999_;
  wire _3000_;
  wire _3001_;
  wire _3002_;
  wire _3003_;
  wire _3004_;
  wire _3005_;
  wire _3006_;
  wire _3007_;
  wire _3008_;
  wire _3009_;
  wire _3010_;
  wire _3011_;
  wire _3012_;
  wire _3013_;
  wire _3014_;
  wire _3015_;
  wire _3016_;
  wire _3017_;
  wire _3018_;
  wire _3019_;
  wire _3020_;
  wire _3021_;
  wire _3022_;
  wire _3023_;
  wire _3024_;
  wire _3025_;
  wire _3026_;
  wire _3027_;
  wire _3028_;
  wire _3029_;
  wire _3030_;
  wire _3031_;
  wire _3032_;
  wire _3033_;
  wire _3034_;
  wire _3035_;
  wire _3036_;
  wire _3037_;
  wire _3038_;
  wire _3039_;
  wire _3040_;
  wire _3041_;
  wire _3042_;
  wire _3043_;
  wire _3044_;
  wire _3045_;
  wire _3046_;
  wire _3047_;
  wire _3048_;
  wire _3049_;
  wire _3050_;
  wire _3051_;
  wire _3052_;
  wire _3053_;
  wire _3054_;
  wire _3055_;
  wire _3056_;
  wire _3057_;
  wire _3058_;
  wire _3059_;
  wire _3060_;
  wire _3061_;
  wire _3062_;
  wire _3063_;
  wire _3064_;
  wire _3065_;
  wire _3066_;
  wire _3067_;
  wire _3068_;
  wire _3069_;
  wire _3070_;
  wire _3071_;
  wire _3072_;
  wire _3073_;
  wire _3074_;
  wire _3075_;
  wire _3076_;
  wire _3077_;
  wire _3078_;
  wire _3079_;
  wire _3080_;
  wire _3081_;
  wire _3082_;
  wire _3083_;
  wire _3084_;
  wire _3085_;
  wire _3086_;
  wire _3087_;
  wire _3088_;
  wire _3089_;
  wire _3090_;
  wire _3091_;
  wire _3092_;
  wire _3093_;
  wire _3094_;
  wire [7:0] _3095_;
  wire [7:0] _3096_;
  wire _3097_;
  wire _3098_;
  wire _3099_;
  wire _3100_;
  wire _3101_;
  wire _3102_;
  wire _3103_;
  wire _3104_;
  wire _3105_;
  wire _3106_;
  wire _3107_;
  wire _3108_;
  wire _3109_;
  wire _3110_;
  wire _3111_;
  wire _3112_;
  wire _3113_;
  wire _3114_;
  wire _3115_;
  wire _3116_;
  wire _3117_;
  wire _3118_;
  wire _3119_;
  wire _3120_;
  wire _3121_;
  wire _3122_;
  wire _3123_;
  wire _3124_;
  wire _3125_;
  wire _3126_;
  wire _3127_;
  wire _3128_;
  wire _3129_;
  wire _3130_;
  wire _3131_;
  wire _3132_;
  wire _3133_;
  wire _3134_;
  wire _3135_;
  wire _3136_;
  wire _3137_;
  wire _3138_;
  wire _3139_;
  wire _3140_;
  wire _3141_;
  wire _3142_;
  wire _3143_;
  wire _3144_;
  wire _3145_;
  wire _3146_;
  wire _3147_;
  wire _3148_;
  wire _3149_;
  wire _3150_;
  wire _3151_;
  wire _3152_;
  wire _3153_;
  wire _3154_;
  wire _3155_;
  wire _3156_;
  wire _3157_;
  wire _3158_;
  wire _3159_;
  wire _3160_;
  wire _3161_;
  wire _3162_;
  wire _3163_;
  wire _3164_;
  wire _3165_;
  wire _3166_;
  wire _3167_;
  wire _3168_;
  wire _3169_;
  wire _3170_;
  wire _3171_;
  wire _3172_;
  wire _3173_;
  wire _3174_;
  wire _3175_;
  wire _3176_;
  wire _3177_;
  wire _3178_;
  wire _3179_;
  wire _3180_;
  wire _3181_;
  wire _3182_;
  wire _3183_;
  wire _3184_;
  wire _3185_;
  wire _3186_;
  wire _3187_;
  wire _3188_;
  wire _3189_;
  wire _3190_;
  wire _3191_;
  wire _3192_;
  wire _3193_;
  wire _3194_;
  wire _3195_;
  wire _3196_;
  wire _3197_;
  wire _3198_;
  wire _3199_;
  wire _3200_;
  wire _3201_;
  wire _3202_;
  wire _3203_;
  wire _3204_;
  wire _3205_;
  wire _3206_;
  wire _3207_;
  wire _3208_;
  wire _3209_;
  wire _3210_;
  wire _3211_;
  wire _3212_;
  wire _3213_;
  wire _3214_;
  wire _3215_;
  wire _3216_;
  wire _3217_;
  wire _3218_;
  wire _3219_;
  wire _3220_;
  wire _3221_;
  wire _3222_;
  wire _3223_;
  wire _3224_;
  wire _3225_;
  wire _3226_;
  wire _3227_;
  wire _3228_;
  wire _3229_;
  wire _3230_;
  wire _3231_;
  wire _3232_;
  wire _3233_;
  wire _3234_;
  wire _3235_;
  wire _3236_;
  wire _3237_;
  wire _3238_;
  wire _3239_;
  wire _3240_;
  wire _3241_;
  wire _3242_;
  wire _3243_;
  wire _3244_;
  wire _3245_;
  wire _3246_;
  wire _3247_;
  wire _3248_;
  wire _3249_;
  wire _3250_;
  wire _3251_;
  wire _3252_;
  wire _3253_;
  wire _3254_;
  wire _3255_;
  wire _3256_;
  wire _3257_;
  wire _3258_;
  wire _3259_;
  wire _3260_;
  wire _3261_;
  wire _3262_;
  wire _3263_;
  wire _3264_;
  wire _3265_;
  wire _3266_;
  wire _3267_;
  wire _3268_;
  wire _3269_;
  wire _3270_;
  wire _3271_;
  wire _3272_;
  wire _3273_;
  wire _3274_;
  wire _3275_;
  wire _3276_;
  wire _3277_;
  wire _3278_;
  wire _3279_;
  wire _3280_;
  wire _3281_;
  wire _3282_;
  wire _3283_;
  wire _3284_;
  wire _3285_;
  wire _3286_;
  wire _3287_;
  wire _3288_;
  wire _3289_;
  wire _3290_;
  wire _3291_;
  wire _3292_;
  wire _3293_;
  wire _3294_;
  wire _3295_;
  wire _3296_;
  wire _3297_;
  wire _3298_;
  wire _3299_;
  wire _3300_;
  wire _3301_;
  wire _3302_;
  wire _3303_;
  wire _3304_;
  wire _3305_;
  wire _3306_;
  wire _3307_;
  wire _3308_;
  wire _3309_;
  wire _3310_;
  wire _3311_;
  wire _3312_;
  wire _3313_;
  wire _3314_;
  wire _3315_;
  wire _3316_;
  wire _3317_;
  wire _3318_;
  wire _3319_;
  wire _3320_;
  wire _3321_;
  wire _3322_;
  wire _3323_;
  wire _3324_;
  wire _3325_;
  wire _3326_;
  wire _3327_;
  wire _3328_;
  wire _3329_;
  wire _3330_;
  wire _3331_;
  wire _3332_;
  wire _3333_;
  wire _3334_;
  wire _3335_;
  wire _3336_;
  wire _3337_;
  wire _3338_;
  wire _3339_;
  wire _3340_;
  wire _3341_;
  wire _3342_;
  wire _3343_;
  wire _3344_;
  wire _3345_;
  wire _3346_;
  wire _3347_;
  wire _3348_;
  wire _3349_;
  wire _3350_;
  wire _3351_;
  wire _3352_;
  wire [7:0] _3353_;
  wire [7:0] _3354_;
  wire _3355_;
  wire _3356_;
  wire _3357_;
  wire _3358_;
  wire _3359_;
  wire _3360_;
  wire _3361_;
  wire _3362_;
  wire _3363_;
  wire _3364_;
  wire _3365_;
  wire _3366_;
  wire _3367_;
  wire _3368_;
  wire _3369_;
  wire _3370_;
  wire _3371_;
  wire _3372_;
  wire _3373_;
  wire _3374_;
  wire _3375_;
  wire _3376_;
  wire _3377_;
  wire _3378_;
  wire _3379_;
  wire _3380_;
  wire _3381_;
  wire _3382_;
  wire _3383_;
  wire _3384_;
  wire _3385_;
  wire _3386_;
  wire _3387_;
  wire _3388_;
  wire _3389_;
  wire _3390_;
  wire _3391_;
  wire _3392_;
  wire _3393_;
  wire _3394_;
  wire _3395_;
  wire _3396_;
  wire _3397_;
  wire _3398_;
  wire _3399_;
  wire _3400_;
  wire _3401_;
  wire _3402_;
  wire _3403_;
  wire _3404_;
  wire _3405_;
  wire _3406_;
  wire _3407_;
  wire _3408_;
  wire _3409_;
  wire _3410_;
  wire _3411_;
  wire _3412_;
  wire _3413_;
  wire _3414_;
  wire _3415_;
  wire _3416_;
  wire _3417_;
  wire _3418_;
  wire _3419_;
  wire _3420_;
  wire _3421_;
  wire _3422_;
  wire _3423_;
  wire _3424_;
  wire _3425_;
  wire _3426_;
  wire _3427_;
  wire _3428_;
  wire _3429_;
  wire _3430_;
  wire _3431_;
  wire _3432_;
  wire _3433_;
  wire _3434_;
  wire _3435_;
  wire _3436_;
  wire _3437_;
  wire _3438_;
  wire _3439_;
  wire _3440_;
  wire _3441_;
  wire _3442_;
  wire _3443_;
  wire _3444_;
  wire _3445_;
  wire _3446_;
  wire _3447_;
  wire _3448_;
  wire _3449_;
  wire _3450_;
  wire _3451_;
  wire _3452_;
  wire _3453_;
  wire _3454_;
  wire _3455_;
  wire _3456_;
  wire _3457_;
  wire _3458_;
  wire _3459_;
  wire _3460_;
  wire _3461_;
  wire _3462_;
  wire _3463_;
  wire _3464_;
  wire _3465_;
  wire _3466_;
  wire _3467_;
  wire _3468_;
  wire _3469_;
  wire _3470_;
  wire _3471_;
  wire _3472_;
  wire _3473_;
  wire _3474_;
  wire _3475_;
  wire _3476_;
  wire _3477_;
  wire _3478_;
  wire _3479_;
  wire _3480_;
  wire _3481_;
  wire _3482_;
  wire _3483_;
  wire _3484_;
  wire _3485_;
  wire _3486_;
  wire _3487_;
  wire _3488_;
  wire _3489_;
  wire _3490_;
  wire _3491_;
  wire _3492_;
  wire _3493_;
  wire _3494_;
  wire _3495_;
  wire _3496_;
  wire _3497_;
  wire _3498_;
  wire _3499_;
  wire _3500_;
  wire _3501_;
  wire _3502_;
  wire _3503_;
  wire _3504_;
  wire _3505_;
  wire _3506_;
  wire _3507_;
  wire _3508_;
  wire _3509_;
  wire _3510_;
  wire _3511_;
  wire _3512_;
  wire _3513_;
  wire _3514_;
  wire _3515_;
  wire _3516_;
  wire _3517_;
  wire _3518_;
  wire _3519_;
  wire _3520_;
  wire _3521_;
  wire _3522_;
  wire _3523_;
  wire _3524_;
  wire _3525_;
  wire _3526_;
  wire _3527_;
  wire _3528_;
  wire _3529_;
  wire _3530_;
  wire _3531_;
  wire _3532_;
  wire _3533_;
  wire _3534_;
  wire _3535_;
  wire _3536_;
  wire _3537_;
  wire _3538_;
  wire _3539_;
  wire _3540_;
  wire _3541_;
  wire _3542_;
  wire _3543_;
  wire _3544_;
  wire _3545_;
  wire _3546_;
  wire _3547_;
  wire _3548_;
  wire _3549_;
  wire _3550_;
  wire _3551_;
  wire _3552_;
  wire _3553_;
  wire _3554_;
  wire _3555_;
  wire _3556_;
  wire _3557_;
  wire _3558_;
  wire _3559_;
  wire _3560_;
  wire _3561_;
  wire _3562_;
  wire _3563_;
  wire _3564_;
  wire _3565_;
  wire _3566_;
  wire _3567_;
  wire _3568_;
  wire _3569_;
  wire _3570_;
  wire _3571_;
  wire _3572_;
  wire _3573_;
  wire _3574_;
  wire _3575_;
  wire _3576_;
  wire _3577_;
  wire _3578_;
  wire _3579_;
  wire _3580_;
  wire _3581_;
  wire _3582_;
  wire _3583_;
  wire _3584_;
  wire _3585_;
  wire _3586_;
  wire _3587_;
  wire _3588_;
  wire _3589_;
  wire _3590_;
  wire _3591_;
  wire _3592_;
  wire _3593_;
  wire _3594_;
  wire _3595_;
  wire _3596_;
  wire _3597_;
  wire _3598_;
  wire _3599_;
  wire _3600_;
  wire _3601_;
  wire _3602_;
  wire _3603_;
  wire _3604_;
  wire _3605_;
  wire _3606_;
  wire _3607_;
  wire _3608_;
  wire _3609_;
  wire _3610_;
  wire [7:0] _3611_;
  wire [7:0] _3612_;
  wire _3613_;
  wire _3614_;
  wire _3615_;
  wire _3616_;
  wire _3617_;
  wire _3618_;
  wire _3619_;
  wire _3620_;
  wire _3621_;
  wire _3622_;
  wire _3623_;
  wire _3624_;
  wire _3625_;
  wire _3626_;
  wire _3627_;
  wire _3628_;
  wire _3629_;
  wire _3630_;
  wire _3631_;
  wire _3632_;
  wire _3633_;
  wire _3634_;
  wire _3635_;
  wire _3636_;
  wire _3637_;
  wire _3638_;
  wire _3639_;
  wire _3640_;
  wire _3641_;
  wire _3642_;
  wire _3643_;
  wire _3644_;
  wire _3645_;
  wire _3646_;
  wire _3647_;
  wire _3648_;
  wire _3649_;
  wire _3650_;
  wire _3651_;
  wire _3652_;
  wire _3653_;
  wire _3654_;
  wire _3655_;
  wire _3656_;
  wire _3657_;
  wire _3658_;
  wire _3659_;
  wire _3660_;
  wire _3661_;
  wire _3662_;
  wire _3663_;
  wire _3664_;
  wire _3665_;
  wire _3666_;
  wire _3667_;
  wire _3668_;
  wire _3669_;
  wire _3670_;
  wire _3671_;
  wire _3672_;
  wire _3673_;
  wire _3674_;
  wire _3675_;
  wire _3676_;
  wire _3677_;
  wire _3678_;
  wire _3679_;
  wire _3680_;
  wire _3681_;
  wire _3682_;
  wire _3683_;
  wire _3684_;
  wire _3685_;
  wire _3686_;
  wire _3687_;
  wire _3688_;
  wire _3689_;
  wire _3690_;
  wire _3691_;
  wire _3692_;
  wire _3693_;
  wire _3694_;
  wire _3695_;
  wire _3696_;
  wire _3697_;
  wire _3698_;
  wire _3699_;
  wire _3700_;
  wire _3701_;
  wire _3702_;
  wire _3703_;
  wire _3704_;
  wire _3705_;
  wire _3706_;
  wire _3707_;
  wire _3708_;
  wire _3709_;
  wire _3710_;
  wire _3711_;
  wire _3712_;
  wire _3713_;
  wire _3714_;
  wire _3715_;
  wire _3716_;
  wire _3717_;
  wire _3718_;
  wire _3719_;
  wire _3720_;
  wire _3721_;
  wire _3722_;
  wire _3723_;
  wire _3724_;
  wire _3725_;
  wire _3726_;
  wire _3727_;
  wire _3728_;
  wire _3729_;
  wire _3730_;
  wire _3731_;
  wire _3732_;
  wire _3733_;
  wire _3734_;
  wire _3735_;
  wire _3736_;
  wire _3737_;
  wire _3738_;
  wire _3739_;
  wire _3740_;
  wire _3741_;
  wire _3742_;
  wire _3743_;
  wire _3744_;
  wire _3745_;
  wire _3746_;
  wire _3747_;
  wire _3748_;
  wire _3749_;
  wire _3750_;
  wire _3751_;
  wire _3752_;
  wire _3753_;
  wire _3754_;
  wire _3755_;
  wire _3756_;
  wire _3757_;
  wire _3758_;
  wire _3759_;
  wire _3760_;
  wire _3761_;
  wire _3762_;
  wire _3763_;
  wire _3764_;
  wire _3765_;
  wire _3766_;
  wire _3767_;
  wire _3768_;
  wire _3769_;
  wire _3770_;
  wire _3771_;
  wire _3772_;
  wire _3773_;
  wire _3774_;
  wire _3775_;
  wire _3776_;
  wire _3777_;
  wire _3778_;
  wire _3779_;
  wire _3780_;
  wire _3781_;
  wire _3782_;
  wire _3783_;
  wire _3784_;
  wire _3785_;
  wire _3786_;
  wire _3787_;
  wire _3788_;
  wire _3789_;
  wire _3790_;
  wire _3791_;
  wire _3792_;
  wire _3793_;
  wire _3794_;
  wire _3795_;
  wire _3796_;
  wire _3797_;
  wire _3798_;
  wire _3799_;
  wire _3800_;
  wire _3801_;
  wire _3802_;
  wire _3803_;
  wire _3804_;
  wire _3805_;
  wire _3806_;
  wire _3807_;
  wire _3808_;
  wire _3809_;
  wire _3810_;
  wire _3811_;
  wire _3812_;
  wire _3813_;
  wire _3814_;
  wire _3815_;
  wire _3816_;
  wire _3817_;
  wire _3818_;
  wire _3819_;
  wire _3820_;
  wire _3821_;
  wire _3822_;
  wire _3823_;
  wire _3824_;
  wire _3825_;
  wire _3826_;
  wire _3827_;
  wire _3828_;
  wire _3829_;
  wire _3830_;
  wire _3831_;
  wire _3832_;
  wire _3833_;
  wire _3834_;
  wire _3835_;
  wire _3836_;
  wire _3837_;
  wire _3838_;
  wire _3839_;
  wire _3840_;
  wire _3841_;
  wire _3842_;
  wire _3843_;
  wire _3844_;
  wire _3845_;
  wire _3846_;
  wire _3847_;
  wire _3848_;
  wire _3849_;
  wire _3850_;
  wire _3851_;
  wire _3852_;
  wire _3853_;
  wire _3854_;
  wire _3855_;
  wire _3856_;
  wire _3857_;
  wire _3858_;
  wire _3859_;
  wire _3860_;
  wire _3861_;
  wire _3862_;
  wire _3863_;
  wire _3864_;
  wire _3865_;
  wire _3866_;
  wire _3867_;
  wire _3868_;
  wire [7:0] _3869_;
  wire [7:0] _3870_;
  wire _3871_;
  wire _3872_;
  wire _3873_;
  wire _3874_;
  wire _3875_;
  wire _3876_;
  wire _3877_;
  wire _3878_;
  wire _3879_;
  wire _3880_;
  wire _3881_;
  wire _3882_;
  wire _3883_;
  wire _3884_;
  wire _3885_;
  wire _3886_;
  wire _3887_;
  wire _3888_;
  wire _3889_;
  wire _3890_;
  wire _3891_;
  wire _3892_;
  wire _3893_;
  wire _3894_;
  wire _3895_;
  wire _3896_;
  wire _3897_;
  wire _3898_;
  wire _3899_;
  wire _3900_;
  wire _3901_;
  wire _3902_;
  wire _3903_;
  wire _3904_;
  wire _3905_;
  wire _3906_;
  wire _3907_;
  wire _3908_;
  wire _3909_;
  wire _3910_;
  wire _3911_;
  wire _3912_;
  wire _3913_;
  wire _3914_;
  wire _3915_;
  wire _3916_;
  wire _3917_;
  wire _3918_;
  wire _3919_;
  wire _3920_;
  wire _3921_;
  wire _3922_;
  wire _3923_;
  wire _3924_;
  wire _3925_;
  wire _3926_;
  wire _3927_;
  wire _3928_;
  wire _3929_;
  wire _3930_;
  wire _3931_;
  wire _3932_;
  wire _3933_;
  wire _3934_;
  wire _3935_;
  wire _3936_;
  wire _3937_;
  wire _3938_;
  wire _3939_;
  wire _3940_;
  wire _3941_;
  wire _3942_;
  wire _3943_;
  wire _3944_;
  wire _3945_;
  wire _3946_;
  wire _3947_;
  wire _3948_;
  wire _3949_;
  wire _3950_;
  wire _3951_;
  wire _3952_;
  wire _3953_;
  wire _3954_;
  wire _3955_;
  wire _3956_;
  wire _3957_;
  wire _3958_;
  wire _3959_;
  wire _3960_;
  wire _3961_;
  wire _3962_;
  wire _3963_;
  wire _3964_;
  wire _3965_;
  wire _3966_;
  wire _3967_;
  wire _3968_;
  wire _3969_;
  wire _3970_;
  wire _3971_;
  wire _3972_;
  wire _3973_;
  wire _3974_;
  wire _3975_;
  wire _3976_;
  wire _3977_;
  wire _3978_;
  wire _3979_;
  wire _3980_;
  wire _3981_;
  wire _3982_;
  wire _3983_;
  wire _3984_;
  wire _3985_;
  wire _3986_;
  wire _3987_;
  wire _3988_;
  wire _3989_;
  wire _3990_;
  wire _3991_;
  wire _3992_;
  wire _3993_;
  wire _3994_;
  wire _3995_;
  wire _3996_;
  wire _3997_;
  wire _3998_;
  wire _3999_;
  wire _4000_;
  wire _4001_;
  wire _4002_;
  wire _4003_;
  wire _4004_;
  wire _4005_;
  wire _4006_;
  wire _4007_;
  wire _4008_;
  wire _4009_;
  wire _4010_;
  wire _4011_;
  wire _4012_;
  wire _4013_;
  wire _4014_;
  wire _4015_;
  wire _4016_;
  wire _4017_;
  wire _4018_;
  wire _4019_;
  wire _4020_;
  wire _4021_;
  wire _4022_;
  wire _4023_;
  wire _4024_;
  wire _4025_;
  wire _4026_;
  wire _4027_;
  wire _4028_;
  wire _4029_;
  wire _4030_;
  wire _4031_;
  wire _4032_;
  wire _4033_;
  wire _4034_;
  wire _4035_;
  wire _4036_;
  wire _4037_;
  wire _4038_;
  wire _4039_;
  wire _4040_;
  wire _4041_;
  wire _4042_;
  wire _4043_;
  wire _4044_;
  wire _4045_;
  wire _4046_;
  wire _4047_;
  wire _4048_;
  wire _4049_;
  wire _4050_;
  wire _4051_;
  wire _4052_;
  wire _4053_;
  wire _4054_;
  wire _4055_;
  wire _4056_;
  wire _4057_;
  wire _4058_;
  wire _4059_;
  wire _4060_;
  wire _4061_;
  wire _4062_;
  wire _4063_;
  wire _4064_;
  wire _4065_;
  wire _4066_;
  wire _4067_;
  wire _4068_;
  wire _4069_;
  wire _4070_;
  wire _4071_;
  wire _4072_;
  wire _4073_;
  wire _4074_;
  wire _4075_;
  wire _4076_;
  wire _4077_;
  wire _4078_;
  wire _4079_;
  wire _4080_;
  wire _4081_;
  wire _4082_;
  wire _4083_;
  wire _4084_;
  wire _4085_;
  wire _4086_;
  wire _4087_;
  wire _4088_;
  wire _4089_;
  wire _4090_;
  wire _4091_;
  wire _4092_;
  wire _4093_;
  wire _4094_;
  wire _4095_;
  wire _4096_;
  wire _4097_;
  wire _4098_;
  wire _4099_;
  wire _4100_;
  wire _4101_;
  wire _4102_;
  wire _4103_;
  wire _4104_;
  wire _4105_;
  wire _4106_;
  wire _4107_;
  wire _4108_;
  wire _4109_;
  wire _4110_;
  wire _4111_;
  wire _4112_;
  wire _4113_;
  wire _4114_;
  wire _4115_;
  wire _4116_;
  wire _4117_;
  wire _4118_;
  wire _4119_;
  wire _4120_;
  wire _4121_;
  wire _4122_;
  wire _4123_;
  wire _4124_;
  wire _4125_;
  wire _4126_;
  wire [7:0] _4127_;
  wire [31:0] _4128_;
  wire [31:0] _4129_;
  wire [31:0] _4130_;
  wire [31:0] _4131_;
  wire [31:0] _4132_;
  wire [31:0] _4133_;
  wire [31:0] _4134_;
  wire [31:0] _4135_;
  wire [31:0] _4136_;
  wire [31:0] _4137_;
  wire [31:0] _4138_;
  wire [31:0] _4139_;
  input clk;
  wire [31:0] k0;
  wire [31:0] k1;
  wire [31:0] k2;
  wire [31:0] k3;
  input [127:0] key;
  wire [31:0] p00;
  wire [31:0] p01;
  wire [31:0] p02;
  wire [31:0] p03;
  wire [31:0] p10;
  wire [31:0] p11;
  wire [31:0] p12;
  wire [31:0] p13;
  wire [31:0] p20;
  wire [31:0] p21;
  wire [31:0] p22;
  wire [31:0] p23;
  wire [31:0] p30;
  wire [31:0] p31;
  wire [31:0] p32;
  wire [31:0] p33;
  wire [31:0] s0;
  wire [31:0] s1;
  wire [31:0] s2;
  wire [31:0] s3;
  input [127:0] state_in;
  output [127:0] state_out;
  reg [127:0] state_out;
  wire [7:0] \t0.b0 ;
  wire [7:0] \t0.b1 ;
  wire [7:0] \t0.b2 ;
  wire [7:0] \t0.b3 ;
  wire \t0.clk ;
  wire [31:0] \t0.p0 ;
  wire [31:0] \t0.p1 ;
  wire [31:0] \t0.p2 ;
  wire [31:0] \t0.p3 ;
  wire [31:0] \t0.state ;
  wire \t0.t0.clk ;
  wire [7:0] \t0.t0.in ;
  wire [31:0] \t0.t0.out ;
  wire \t0.t0.s0.clk ;
  wire [7:0] \t0.t0.s0.in ;
  reg [7:0] \t0.t0.s0.out ;
  wire \t0.t0.s4.clk ;
  wire [7:0] \t0.t0.s4.in ;
  reg [7:0] \t0.t0.s4.out ;
  wire \t0.t1.clk ;
  wire [7:0] \t0.t1.in ;
  wire [31:0] \t0.t1.out ;
  wire \t0.t1.s0.clk ;
  wire [7:0] \t0.t1.s0.in ;
  reg [7:0] \t0.t1.s0.out ;
  wire \t0.t1.s4.clk ;
  wire [7:0] \t0.t1.s4.in ;
  reg [7:0] \t0.t1.s4.out ;
  wire \t0.t2.clk ;
  wire [7:0] \t0.t2.in ;
  wire [31:0] \t0.t2.out ;
  wire \t0.t2.s0.clk ;
  wire [7:0] \t0.t2.s0.in ;
  reg [7:0] \t0.t2.s0.out ;
  wire \t0.t2.s4.clk ;
  wire [7:0] \t0.t2.s4.in ;
  reg [7:0] \t0.t2.s4.out ;
  wire \t0.t3.clk ;
  wire [7:0] \t0.t3.in ;
  wire [31:0] \t0.t3.out ;
  wire \t0.t3.s0.clk ;
  wire [7:0] \t0.t3.s0.in ;
  reg [7:0] \t0.t3.s0.out ;
  wire \t0.t3.s4.clk ;
  wire [7:0] \t0.t3.s4.in ;
  reg [7:0] \t0.t3.s4.out ;
  wire [7:0] \t1.b0 ;
  wire [7:0] \t1.b1 ;
  wire [7:0] \t1.b2 ;
  wire [7:0] \t1.b3 ;
  wire \t1.clk ;
  wire [31:0] \t1.p0 ;
  wire [31:0] \t1.p1 ;
  wire [31:0] \t1.p2 ;
  wire [31:0] \t1.p3 ;
  wire [31:0] \t1.state ;
  wire \t1.t0.clk ;
  wire [7:0] \t1.t0.in ;
  wire [31:0] \t1.t0.out ;
  wire \t1.t0.s0.clk ;
  wire [7:0] \t1.t0.s0.in ;
  reg [7:0] \t1.t0.s0.out ;
  wire \t1.t0.s4.clk ;
  wire [7:0] \t1.t0.s4.in ;
  reg [7:0] \t1.t0.s4.out ;
  wire \t1.t1.clk ;
  wire [7:0] \t1.t1.in ;
  wire [31:0] \t1.t1.out ;
  wire \t1.t1.s0.clk ;
  wire [7:0] \t1.t1.s0.in ;
  reg [7:0] \t1.t1.s0.out ;
  wire \t1.t1.s4.clk ;
  wire [7:0] \t1.t1.s4.in ;
  reg [7:0] \t1.t1.s4.out ;
  wire \t1.t2.clk ;
  wire [7:0] \t1.t2.in ;
  wire [31:0] \t1.t2.out ;
  wire \t1.t2.s0.clk ;
  wire [7:0] \t1.t2.s0.in ;
  reg [7:0] \t1.t2.s0.out ;
  wire \t1.t2.s4.clk ;
  wire [7:0] \t1.t2.s4.in ;
  reg [7:0] \t1.t2.s4.out ;
  wire \t1.t3.clk ;
  wire [7:0] \t1.t3.in ;
  wire [31:0] \t1.t3.out ;
  wire \t1.t3.s0.clk ;
  wire [7:0] \t1.t3.s0.in ;
  reg [7:0] \t1.t3.s0.out ;
  wire \t1.t3.s4.clk ;
  wire [7:0] \t1.t3.s4.in ;
  reg [7:0] \t1.t3.s4.out ;
  wire [7:0] \t2.b0 ;
  wire [7:0] \t2.b1 ;
  wire [7:0] \t2.b2 ;
  wire [7:0] \t2.b3 ;
  wire \t2.clk ;
  wire [31:0] \t2.p0 ;
  wire [31:0] \t2.p1 ;
  wire [31:0] \t2.p2 ;
  wire [31:0] \t2.p3 ;
  wire [31:0] \t2.state ;
  wire \t2.t0.clk ;
  wire [7:0] \t2.t0.in ;
  wire [31:0] \t2.t0.out ;
  wire \t2.t0.s0.clk ;
  wire [7:0] \t2.t0.s0.in ;
  reg [7:0] \t2.t0.s0.out ;
  wire \t2.t0.s4.clk ;
  wire [7:0] \t2.t0.s4.in ;
  reg [7:0] \t2.t0.s4.out ;
  wire \t2.t1.clk ;
  wire [7:0] \t2.t1.in ;
  wire [31:0] \t2.t1.out ;
  wire \t2.t1.s0.clk ;
  wire [7:0] \t2.t1.s0.in ;
  reg [7:0] \t2.t1.s0.out ;
  wire \t2.t1.s4.clk ;
  wire [7:0] \t2.t1.s4.in ;
  reg [7:0] \t2.t1.s4.out ;
  wire \t2.t2.clk ;
  wire [7:0] \t2.t2.in ;
  wire [31:0] \t2.t2.out ;
  wire \t2.t2.s0.clk ;
  wire [7:0] \t2.t2.s0.in ;
  reg [7:0] \t2.t2.s0.out ;
  wire \t2.t2.s4.clk ;
  wire [7:0] \t2.t2.s4.in ;
  reg [7:0] \t2.t2.s4.out ;
  wire \t2.t3.clk ;
  wire [7:0] \t2.t3.in ;
  wire [31:0] \t2.t3.out ;
  wire \t2.t3.s0.clk ;
  wire [7:0] \t2.t3.s0.in ;
  reg [7:0] \t2.t3.s0.out ;
  wire \t2.t3.s4.clk ;
  wire [7:0] \t2.t3.s4.in ;
  reg [7:0] \t2.t3.s4.out ;
  wire [7:0] \t3.b0 ;
  wire [7:0] \t3.b1 ;
  wire [7:0] \t3.b2 ;
  wire [7:0] \t3.b3 ;
  wire \t3.clk ;
  wire [31:0] \t3.p0 ;
  wire [31:0] \t3.p1 ;
  wire [31:0] \t3.p2 ;
  wire [31:0] \t3.p3 ;
  wire [31:0] \t3.state ;
  wire \t3.t0.clk ;
  wire [7:0] \t3.t0.in ;
  wire [31:0] \t3.t0.out ;
  wire \t3.t0.s0.clk ;
  wire [7:0] \t3.t0.s0.in ;
  reg [7:0] \t3.t0.s0.out ;
  wire \t3.t0.s4.clk ;
  wire [7:0] \t3.t0.s4.in ;
  reg [7:0] \t3.t0.s4.out ;
  wire \t3.t1.clk ;
  wire [7:0] \t3.t1.in ;
  wire [31:0] \t3.t1.out ;
  wire \t3.t1.s0.clk ;
  wire [7:0] \t3.t1.s0.in ;
  reg [7:0] \t3.t1.s0.out ;
  wire \t3.t1.s4.clk ;
  wire [7:0] \t3.t1.s4.in ;
  reg [7:0] \t3.t1.s4.out ;
  wire \t3.t2.clk ;
  wire [7:0] \t3.t2.in ;
  wire [31:0] \t3.t2.out ;
  wire \t3.t2.s0.clk ;
  wire [7:0] \t3.t2.s0.in ;
  reg [7:0] \t3.t2.s0.out ;
  wire \t3.t2.s4.clk ;
  wire [7:0] \t3.t2.s4.in ;
  reg [7:0] \t3.t2.s4.out ;
  wire \t3.t3.clk ;
  wire [7:0] \t3.t3.in ;
  wire [31:0] \t3.t3.out ;
  wire \t3.t3.s0.clk ;
  wire [7:0] \t3.t3.s0.in ;
  reg [7:0] \t3.t3.s0.out ;
  wire \t3.t3.s4.clk ;
  wire [7:0] \t3.t3.s4.in ;
  reg [7:0] \t3.t3.s4.out ;
  wire [31:0] z0;
  wire [31:0] z1;
  wire [31:0] z2;
  wire [31:0] z3;

  wire [127:0] fangyuan0;
  assign fangyuan0 = { z0, z1, z2, z3 };
  always @(posedge clk)
      state_out <= fangyuan0;
  assign p00[7:0] = \t0.t0.s0.out ^ \t0.t0.s4.out ;
  always @(posedge clk)
      \t0.t0.s0.out <= _0000_;
  wire [255:0] fangyuan1;
  assign fangyuan1 = { _0256_, _0255_, _0254_, _0253_, _0252_, _0251_, _0250_, _0249_, _0248_, _0247_, _0246_, _0245_, _0244_, _0243_, _0242_, _0241_, _0240_, _0239_, _0238_, _0237_, _0236_, _0235_, _0234_, _0233_, _0232_, _0231_, _0230_, _0229_, _0228_, _0227_, _0226_, _0225_, _0224_, _0223_, _0222_, _0221_, _0220_, _0219_, _0218_, _0217_, _0216_, _0215_, _0214_, _0213_, _0212_, _0211_, _0210_, _0209_, _0208_, _0207_, _0206_, _0205_, _0204_, _0203_, _0202_, _0201_, _0200_, _0199_, _0198_, _0197_, _0196_, _0195_, _0194_, _0193_, _0192_, _0191_, _0190_, _0189_, _0188_, _0187_, _0186_, _0185_, _0184_, _0183_, _0182_, _0181_, _0180_, _0179_, _0178_, _0177_, _0176_, _0175_, _0174_, _0173_, _0172_, _0171_, _0170_, _0169_, _0168_, _0167_, _0166_, _0165_, _0164_, _0163_, _0162_, _0161_, _0160_, _0159_, _0158_, _0157_, _0156_, _0155_, _0154_, _0153_, _0152_, _0151_, _0150_, _0149_, _0148_, _0147_, _0146_, _0145_, _0144_, _0143_, _0142_, _0141_, _0140_, _0139_, _0138_, _0137_, _0136_, _0135_, _0134_, _0133_, _0132_, _0131_, _0130_, _0129_, _0128_, _0127_, _0126_, _0125_, _0124_, _0123_, _0122_, _0121_, _0120_, _0119_, _0118_, _0117_, _0116_, _0115_, _0114_, _0113_, _0112_, _0111_, _0110_, _0109_, _0108_, _0107_, _0106_, _0105_, _0104_, _0103_, _0102_, _0101_, _0100_, _0099_, _0098_, _0097_, _0096_, _0095_, _0094_, _0093_, _0092_, _0091_, _0090_, _0089_, _0088_, _0087_, _0086_, _0085_, _0084_, _0083_, _0082_, _0081_, _0080_, _0079_, _0078_, _0077_, _0076_, _0075_, _0074_, _0073_, _0072_, _0071_, _0070_, _0069_, _0068_, _0067_, _0066_, _0065_, _0064_, _0063_, _0062_, _0061_, _0060_, _0059_, _0058_, _0057_, _0056_, _0055_, _0054_, _0053_, _0052_, _0051_, _0050_, _0049_, _0048_, _0047_, _0046_, _0045_, _0044_, _0043_, _0042_, _0041_, _0040_, _0039_, _0038_, _0037_, _0036_, _0035_, _0034_, _0033_, _0032_, _0031_, _0030_, _0029_, _0028_, _0027_, _0026_, _0025_, _0024_, _0023_, _0022_, _0021_, _0020_, _0019_, _0018_, _0017_, _0016_, _0015_, _0014_, _0013_, _0012_, _0011_, _0010_, _0009_, _0008_, _0007_, _0006_, _0005_, _0004_, _0003_, _0002_, _0001_ };

  always @(\t0.t0.s0.out or fangyuan1) begin
    casez (fangyuan1)
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1 :
        _0000_ = 8'b00010110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1? :
        _0000_ = 8'b10111011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?? :
        _0000_ = 8'b01010100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??? :
        _0000_ = 8'b10110000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???? :
        _0000_ = 8'b00001111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????? :
        _0000_ = 8'b00101101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????? :
        _0000_ = 8'b10011001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????? :
        _0000_ = 8'b01000001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????? :
        _0000_ = 8'b01101000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????? :
        _0000_ = 8'b01000010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????? :
        _0000_ = 8'b11100110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????? :
        _0000_ = 8'b10111111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????? :
        _0000_ = 8'b00001101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????? :
        _0000_ = 8'b10001001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????? :
        _0000_ = 8'b10100001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????? :
        _0000_ = 8'b10001100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????? :
        _0000_ = 8'b11011111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????? :
        _0000_ = 8'b00101000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????? :
        _0000_ = 8'b01010101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????? :
        _0000_ = 8'b11001110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????? :
        _0000_ = 8'b11101001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????? :
        _0000_ = 8'b10000111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????? :
        _0000_ = 8'b00011110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????? :
        _0000_ = 8'b10011011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????? :
        _0000_ = 8'b10010100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????? :
        _0000_ = 8'b10001110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????? :
        _0000_ = 8'b11011001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????? :
        _0000_ = 8'b01101001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????? :
        _0000_ = 8'b00010001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????? :
        _0000_ = 8'b10011000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????? :
        _0000_ = 8'b11111000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????? :
        _0000_ = 8'b11100001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????? :
        _0000_ = 8'b10011110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????? :
        _0000_ = 8'b00011101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????? :
        _0000_ = 8'b11000001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????? :
        _0000_ = 8'b10000110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????? :
        _0000_ = 8'b10111001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????? :
        _0000_ = 8'b01010111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????? :
        _0000_ = 8'b00110101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????? :
        _0000_ = 8'b01100001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????? :
        _0000_ = 8'b00001110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????? :
        _0000_ = 8'b11110110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????? :
        _0000_ = 8'b00000011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????? :
        _0000_ = 8'b01001000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????? :
        _0000_ = 8'b01100110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????? :
        _0000_ = 8'b10110101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????? :
        _0000_ = 8'b00111110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????? :
        _0000_ = 8'b01110000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????? :
        _0000_ = 8'b10001010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????? :
        _0000_ = 8'b10001011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????? :
        _0000_ = 8'b10111101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????? :
        _0000_ = 8'b01001011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????? :
        _0000_ = 8'b00011111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????? :
        _0000_ = 8'b01110100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????? :
        _0000_ = 8'b11011101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????? :
        _0000_ = 8'b11101000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????? :
        _0000_ = 8'b11000110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????? :
        _0000_ = 8'b10110100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????? :
        _0000_ = 8'b10100110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????? :
        _0000_ = 8'b00011100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????? :
        _0000_ = 8'b00101110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????? :
        _0000_ = 8'b00100101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????? :
        _0000_ = 8'b01111000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????? :
        _0000_ = 8'b10111010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????? :
        _0000_ = 8'b00001000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b10101110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b01111010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b01100101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b11101010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b11110100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b01010110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b01101100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b10101001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b01001110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b11010101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b10001101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b01101101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b00110111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b11001000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b11100111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b01111001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b11100100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b10010101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b10010001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b01100010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b10101100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b11010011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b11000010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b01011100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b00100100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b00000110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b01001001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b00001010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b00111010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b00110010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b11100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b11011011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b00001011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b01011110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b11011110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b00010100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b10111000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b11101110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b01000110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b10001000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b10010000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b00101010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b00100010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b11011100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b01001111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b10000001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b01100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b01110011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b00011001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b01011101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b01100100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b00111101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b01111110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b10100111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b11000100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b00010111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b01000100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b10010111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b01011111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b11101100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b00010011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b00001100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b11001101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b11010010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b11110011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b11111111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b00010000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b00100001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b11011010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b10110110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b10111100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b11110101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b00111000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b10011101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b10010010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b10001111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b01000000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b10100011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b01010001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b10101000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b10011111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b00111100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b01010000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b01111111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b00000010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b11111001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b01000101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b10000101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b00110011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b01001101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b01000011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b11111011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b10101010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b11101111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b11010000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b11001111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b01011000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b01001100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b01001010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b00111001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b10111110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b11001011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b01101010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b01011011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b10110001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b11111100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b00100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b11101101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b00000000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b11010001 ;
      256'b????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b01010011 ;
      256'b???????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b10000100 ;
      256'b??????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b00101111 ;
      256'b?????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b11100011 ;
      256'b????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b00101001 ;
      256'b???????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b10110011 ;
      256'b??????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b11010110 ;
      256'b?????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b00111011 ;
      256'b????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b01010010 ;
      256'b???????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b10100000 ;
      256'b??????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b01011010 ;
      256'b?????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b01101110 ;
      256'b????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b00011011 ;
      256'b???????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b00011010 ;
      256'b??????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b00101100 ;
      256'b?????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b10000011 ;
      256'b????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b00001001 ;
      256'b???????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b01110101 ;
      256'b??????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b10110010 ;
      256'b?????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b00100111 ;
      256'b????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b11101011 ;
      256'b???????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b11100010 ;
      256'b??????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b10000000 ;
      256'b?????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b00010010 ;
      256'b????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b00000111 ;
      256'b???????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b10011010 ;
      256'b??????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b00000101 ;
      256'b?????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b10010110 ;
      256'b????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b00011000 ;
      256'b???????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b11000011 ;
      256'b??????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b00100011 ;
      256'b?????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b11000111 ;
      256'b????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b00000100 ;
      256'b???????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b00010101 ;
      256'b??????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b00110001 ;
      256'b?????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b11011000 ;
      256'b????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b01110001 ;
      256'b???????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b11110001 ;
      256'b??????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b11100101 ;
      256'b?????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b10100101 ;
      256'b????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b00110100 ;
      256'b???????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b11001100 ;
      256'b??????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b11110111 ;
      256'b?????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b00111111 ;
      256'b????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b00110110 ;
      256'b???????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b00100110 ;
      256'b??????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b10010011 ;
      256'b?????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b11111101 ;
      256'b????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b10110111 ;
      256'b???????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b11000000 ;
      256'b??????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b01110010 ;
      256'b?????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b10100100 ;
      256'b????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b10011100 ;
      256'b???????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b10101111 ;
      256'b??????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b10100010 ;
      256'b?????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b11010100 ;
      256'b????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b10101101 ;
      256'b???????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b11110000 ;
      256'b??????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b01000111 ;
      256'b?????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b01011001 ;
      256'b????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b11111010 ;
      256'b???????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b01111101 ;
      256'b??????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b11001001 ;
      256'b?????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b10000010 ;
      256'b????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b11001010 ;
      256'b???????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b01110110 ;
      256'b??????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b10101011 ;
      256'b?????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b11010111 ;
      256'b????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b11111110 ;
      256'b???????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b00101011 ;
      256'b??????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b01100111 ;
      256'b?????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b00000001 ;
      256'b????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b00110000 ;
      256'b???????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b11000101 ;
      256'b??????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b01101111 ;
      256'b?????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b01101011 ;
      256'b????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b11110010 ;
      256'b???1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b01111011 ;
      256'b??1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b01110111 ;
      256'b?1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b01111100 ;
      256'b1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b01100011 ;
      default:
        _0000_ = \t0.t0.s0.out ;
    endcase
  end
  assign _0001_ = state_in[127:120] == 8'b11111111;
  assign _0002_ = state_in[127:120] == 8'b11111110;
  assign _0003_ = state_in[127:120] == 8'b11111101;
  assign _0004_ = state_in[127:120] == 8'b11111100;
  assign _0005_ = state_in[127:120] == 8'b11111011;
  assign _0006_ = state_in[127:120] == 8'b11111010;
  assign _0007_ = state_in[127:120] == 8'b11111001;
  assign _0008_ = state_in[127:120] == 8'b11111000;
  assign _0009_ = state_in[127:120] == 8'b11110111;
  assign _0010_ = state_in[127:120] == 8'b11110110;
  assign _0011_ = state_in[127:120] == 8'b11110101;
  assign _0012_ = state_in[127:120] == 8'b11110100;
  assign _0013_ = state_in[127:120] == 8'b11110011;
  assign _0014_ = state_in[127:120] == 8'b11110010;
  assign _0015_ = state_in[127:120] == 8'b11110001;
  assign _0016_ = state_in[127:120] == 8'b11110000;
  assign _0017_ = state_in[127:120] == 8'b11101111;
  assign _0018_ = state_in[127:120] == 8'b11101110;
  assign _0019_ = state_in[127:120] == 8'b11101101;
  assign _0020_ = state_in[127:120] == 8'b11101100;
  assign _0021_ = state_in[127:120] == 8'b11101011;
  assign _0022_ = state_in[127:120] == 8'b11101010;
  assign _0023_ = state_in[127:120] == 8'b11101001;
  assign _0024_ = state_in[127:120] == 8'b11101000;
  assign _0025_ = state_in[127:120] == 8'b11100111;
  assign _0026_ = state_in[127:120] == 8'b11100110;
  assign _0027_ = state_in[127:120] == 8'b11100101;
  assign _0028_ = state_in[127:120] == 8'b11100100;
  assign _0029_ = state_in[127:120] == 8'b11100011;
  assign _0030_ = state_in[127:120] == 8'b11100010;
  assign _0031_ = state_in[127:120] == 8'b11100001;
  assign _0032_ = state_in[127:120] == 8'b11100000;
  assign _0033_ = state_in[127:120] == 8'b11011111;
  assign _0034_ = state_in[127:120] == 8'b11011110;
  assign _0035_ = state_in[127:120] == 8'b11011101;
  assign _0036_ = state_in[127:120] == 8'b11011100;
  assign _0037_ = state_in[127:120] == 8'b11011011;
  assign _0038_ = state_in[127:120] == 8'b11011010;
  assign _0039_ = state_in[127:120] == 8'b11011001;
  assign _0040_ = state_in[127:120] == 8'b11011000;
  assign _0041_ = state_in[127:120] == 8'b11010111;
  assign _0042_ = state_in[127:120] == 8'b11010110;
  assign _0043_ = state_in[127:120] == 8'b11010101;
  assign _0044_ = state_in[127:120] == 8'b11010100;
  assign _0045_ = state_in[127:120] == 8'b11010011;
  assign _0046_ = state_in[127:120] == 8'b11010010;
  assign _0047_ = state_in[127:120] == 8'b11010001;
  assign _0048_ = state_in[127:120] == 8'b11010000;
  assign _0049_ = state_in[127:120] == 8'b11001111;
  assign _0050_ = state_in[127:120] == 8'b11001110;
  assign _0051_ = state_in[127:120] == 8'b11001101;
  assign _0052_ = state_in[127:120] == 8'b11001100;
  assign _0053_ = state_in[127:120] == 8'b11001011;
  assign _0054_ = state_in[127:120] == 8'b11001010;
  assign _0055_ = state_in[127:120] == 8'b11001001;
  assign _0056_ = state_in[127:120] == 8'b11001000;
  assign _0057_ = state_in[127:120] == 8'b11000111;
  assign _0058_ = state_in[127:120] == 8'b11000110;
  assign _0059_ = state_in[127:120] == 8'b11000101;
  assign _0060_ = state_in[127:120] == 8'b11000100;
  assign _0061_ = state_in[127:120] == 8'b11000011;
  assign _0062_ = state_in[127:120] == 8'b11000010;
  assign _0063_ = state_in[127:120] == 8'b11000001;
  assign _0064_ = state_in[127:120] == 8'b11000000;
  assign _0065_ = state_in[127:120] == 8'b10111111;
  assign _0066_ = state_in[127:120] == 8'b10111110;
  assign _0067_ = state_in[127:120] == 8'b10111101;
  assign _0068_ = state_in[127:120] == 8'b10111100;
  assign _0069_ = state_in[127:120] == 8'b10111011;
  assign _0070_ = state_in[127:120] == 8'b10111010;
  assign _0071_ = state_in[127:120] == 8'b10111001;
  assign _0072_ = state_in[127:120] == 8'b10111000;
  assign _0073_ = state_in[127:120] == 8'b10110111;
  assign _0074_ = state_in[127:120] == 8'b10110110;
  assign _0075_ = state_in[127:120] == 8'b10110101;
  assign _0076_ = state_in[127:120] == 8'b10110100;
  assign _0077_ = state_in[127:120] == 8'b10110011;
  assign _0078_ = state_in[127:120] == 8'b10110010;
  assign _0079_ = state_in[127:120] == 8'b10110001;
  assign _0080_ = state_in[127:120] == 8'b10110000;
  assign _0081_ = state_in[127:120] == 8'b10101111;
  assign _0082_ = state_in[127:120] == 8'b10101110;
  assign _0083_ = state_in[127:120] == 8'b10101101;
  assign _0084_ = state_in[127:120] == 8'b10101100;
  assign _0085_ = state_in[127:120] == 8'b10101011;
  assign _0086_ = state_in[127:120] == 8'b10101010;
  assign _0087_ = state_in[127:120] == 8'b10101001;
  assign _0088_ = state_in[127:120] == 8'b10101000;
  assign _0089_ = state_in[127:120] == 8'b10100111;
  assign _0090_ = state_in[127:120] == 8'b10100110;
  assign _0091_ = state_in[127:120] == 8'b10100101;
  assign _0092_ = state_in[127:120] == 8'b10100100;
  assign _0093_ = state_in[127:120] == 8'b10100011;
  assign _0094_ = state_in[127:120] == 8'b10100010;
  assign _0095_ = state_in[127:120] == 8'b10100001;
  assign _0096_ = state_in[127:120] == 8'b10100000;
  assign _0097_ = state_in[127:120] == 8'b10011111;
  assign _0098_ = state_in[127:120] == 8'b10011110;
  assign _0099_ = state_in[127:120] == 8'b10011101;
  assign _0100_ = state_in[127:120] == 8'b10011100;
  assign _0101_ = state_in[127:120] == 8'b10011011;
  assign _0102_ = state_in[127:120] == 8'b10011010;
  assign _0103_ = state_in[127:120] == 8'b10011001;
  assign _0104_ = state_in[127:120] == 8'b10011000;
  assign _0105_ = state_in[127:120] == 8'b10010111;
  assign _0106_ = state_in[127:120] == 8'b10010110;
  assign _0107_ = state_in[127:120] == 8'b10010101;
  assign _0108_ = state_in[127:120] == 8'b10010100;
  assign _0109_ = state_in[127:120] == 8'b10010011;
  assign _0110_ = state_in[127:120] == 8'b10010010;
  assign _0111_ = state_in[127:120] == 8'b10010001;
  assign _0112_ = state_in[127:120] == 8'b10010000;
  assign _0113_ = state_in[127:120] == 8'b10001111;
  assign _0114_ = state_in[127:120] == 8'b10001110;
  assign _0115_ = state_in[127:120] == 8'b10001101;
  assign _0116_ = state_in[127:120] == 8'b10001100;
  assign _0117_ = state_in[127:120] == 8'b10001011;
  assign _0118_ = state_in[127:120] == 8'b10001010;
  assign _0119_ = state_in[127:120] == 8'b10001001;
  assign _0120_ = state_in[127:120] == 8'b10001000;
  assign _0121_ = state_in[127:120] == 8'b10000111;
  assign _0122_ = state_in[127:120] == 8'b10000110;
  assign _0123_ = state_in[127:120] == 8'b10000101;
  assign _0124_ = state_in[127:120] == 8'b10000100;
  assign _0125_ = state_in[127:120] == 8'b10000011;
  assign _0126_ = state_in[127:120] == 8'b10000010;
  assign _0127_ = state_in[127:120] == 8'b10000001;
  assign _0128_ = state_in[127:120] == 8'b10000000;
  assign _0129_ = state_in[127:120] == 7'b1111111;
  assign _0130_ = state_in[127:120] == 7'b1111110;
  assign _0131_ = state_in[127:120] == 7'b1111101;
  assign _0132_ = state_in[127:120] == 7'b1111100;
  assign _0133_ = state_in[127:120] == 7'b1111011;
  assign _0134_ = state_in[127:120] == 7'b1111010;
  assign _0135_ = state_in[127:120] == 7'b1111001;
  assign _0136_ = state_in[127:120] == 7'b1111000;
  assign _0137_ = state_in[127:120] == 7'b1110111;
  assign _0138_ = state_in[127:120] == 7'b1110110;
  assign _0139_ = state_in[127:120] == 7'b1110101;
  assign _0140_ = state_in[127:120] == 7'b1110100;
  assign _0141_ = state_in[127:120] == 7'b1110011;
  assign _0142_ = state_in[127:120] == 7'b1110010;
  assign _0143_ = state_in[127:120] == 7'b1110001;
  assign _0144_ = state_in[127:120] == 7'b1110000;
  assign _0145_ = state_in[127:120] == 7'b1101111;
  assign _0146_ = state_in[127:120] == 7'b1101110;
  assign _0147_ = state_in[127:120] == 7'b1101101;
  assign _0148_ = state_in[127:120] == 7'b1101100;
  assign _0149_ = state_in[127:120] == 7'b1101011;
  assign _0150_ = state_in[127:120] == 7'b1101010;
  assign _0151_ = state_in[127:120] == 7'b1101001;
  assign _0152_ = state_in[127:120] == 7'b1101000;
  assign _0153_ = state_in[127:120] == 7'b1100111;
  assign _0154_ = state_in[127:120] == 7'b1100110;
  assign _0155_ = state_in[127:120] == 7'b1100101;
  assign _0156_ = state_in[127:120] == 7'b1100100;
  assign _0157_ = state_in[127:120] == 7'b1100011;
  assign _0158_ = state_in[127:120] == 7'b1100010;
  assign _0159_ = state_in[127:120] == 7'b1100001;
  assign _0160_ = state_in[127:120] == 7'b1100000;
  assign _0161_ = state_in[127:120] == 7'b1011111;
  assign _0162_ = state_in[127:120] == 7'b1011110;
  assign _0163_ = state_in[127:120] == 7'b1011101;
  assign _0164_ = state_in[127:120] == 7'b1011100;
  assign _0165_ = state_in[127:120] == 7'b1011011;
  assign _0166_ = state_in[127:120] == 7'b1011010;
  assign _0167_ = state_in[127:120] == 7'b1011001;
  assign _0168_ = state_in[127:120] == 7'b1011000;
  assign _0169_ = state_in[127:120] == 7'b1010111;
  assign _0170_ = state_in[127:120] == 7'b1010110;
  assign _0171_ = state_in[127:120] == 7'b1010101;
  assign _0172_ = state_in[127:120] == 7'b1010100;
  assign _0173_ = state_in[127:120] == 7'b1010011;
  assign _0174_ = state_in[127:120] == 7'b1010010;
  assign _0175_ = state_in[127:120] == 7'b1010001;
  assign _0176_ = state_in[127:120] == 7'b1010000;
  assign _0177_ = state_in[127:120] == 7'b1001111;
  assign _0178_ = state_in[127:120] == 7'b1001110;
  assign _0179_ = state_in[127:120] == 7'b1001101;
  assign _0180_ = state_in[127:120] == 7'b1001100;
  assign _0181_ = state_in[127:120] == 7'b1001011;
  assign _0182_ = state_in[127:120] == 7'b1001010;
  assign _0183_ = state_in[127:120] == 7'b1001001;
  assign _0184_ = state_in[127:120] == 7'b1001000;
  assign _0185_ = state_in[127:120] == 7'b1000111;
  assign _0186_ = state_in[127:120] == 7'b1000110;
  assign _0187_ = state_in[127:120] == 7'b1000101;
  assign _0188_ = state_in[127:120] == 7'b1000100;
  assign _0189_ = state_in[127:120] == 7'b1000011;
  assign _0190_ = state_in[127:120] == 7'b1000010;
  assign _0191_ = state_in[127:120] == 7'b1000001;
  assign _0192_ = state_in[127:120] == 7'b1000000;
  assign _0193_ = state_in[127:120] == 6'b111111;
  assign _0194_ = state_in[127:120] == 6'b111110;
  assign _0195_ = state_in[127:120] == 6'b111101;
  assign _0196_ = state_in[127:120] == 6'b111100;
  assign _0197_ = state_in[127:120] == 6'b111011;
  assign _0198_ = state_in[127:120] == 6'b111010;
  assign _0199_ = state_in[127:120] == 6'b111001;
  assign _0200_ = state_in[127:120] == 6'b111000;
  assign _0201_ = state_in[127:120] == 6'b110111;
  assign _0202_ = state_in[127:120] == 6'b110110;
  assign _0203_ = state_in[127:120] == 6'b110101;
  assign _0204_ = state_in[127:120] == 6'b110100;
  assign _0205_ = state_in[127:120] == 6'b110011;
  assign _0206_ = state_in[127:120] == 6'b110010;
  assign _0207_ = state_in[127:120] == 6'b110001;
  assign _0208_ = state_in[127:120] == 6'b110000;
  assign _0209_ = state_in[127:120] == 6'b101111;
  assign _0210_ = state_in[127:120] == 6'b101110;
  assign _0211_ = state_in[127:120] == 6'b101101;
  assign _0212_ = state_in[127:120] == 6'b101100;
  assign _0213_ = state_in[127:120] == 6'b101011;
  assign _0214_ = state_in[127:120] == 6'b101010;
  assign _0215_ = state_in[127:120] == 6'b101001;
  assign _0216_ = state_in[127:120] == 6'b101000;
  assign _0217_ = state_in[127:120] == 6'b100111;
  assign _0218_ = state_in[127:120] == 6'b100110;
  assign _0219_ = state_in[127:120] == 6'b100101;
  assign _0220_ = state_in[127:120] == 6'b100100;
  assign _0221_ = state_in[127:120] == 6'b100011;
  assign _0222_ = state_in[127:120] == 6'b100010;
  assign _0223_ = state_in[127:120] == 6'b100001;
  assign _0224_ = state_in[127:120] == 6'b100000;
  assign _0225_ = state_in[127:120] == 5'b11111;
  assign _0226_ = state_in[127:120] == 5'b11110;
  assign _0227_ = state_in[127:120] == 5'b11101;
  assign _0228_ = state_in[127:120] == 5'b11100;
  assign _0229_ = state_in[127:120] == 5'b11011;
  assign _0230_ = state_in[127:120] == 5'b11010;
  assign _0231_ = state_in[127:120] == 5'b11001;
  assign _0232_ = state_in[127:120] == 5'b11000;
  assign _0233_ = state_in[127:120] == 5'b10111;
  assign _0234_ = state_in[127:120] == 5'b10110;
  assign _0235_ = state_in[127:120] == 5'b10101;
  assign _0236_ = state_in[127:120] == 5'b10100;
  assign _0237_ = state_in[127:120] == 5'b10011;
  assign _0238_ = state_in[127:120] == 5'b10010;
  assign _0239_ = state_in[127:120] == 5'b10001;
  assign _0240_ = state_in[127:120] == 5'b10000;
  assign _0241_ = state_in[127:120] == 4'b1111;
  assign _0242_ = state_in[127:120] == 4'b1110;
  assign _0243_ = state_in[127:120] == 4'b1101;
  assign _0244_ = state_in[127:120] == 4'b1100;
  assign _0245_ = state_in[127:120] == 4'b1011;
  assign _0246_ = state_in[127:120] == 4'b1010;
  assign _0247_ = state_in[127:120] == 4'b1001;
  assign _0248_ = state_in[127:120] == 4'b1000;
  assign _0249_ = state_in[127:120] == 3'b111;
  assign _0250_ = state_in[127:120] == 3'b110;
  assign _0251_ = state_in[127:120] == 3'b101;
  assign _0252_ = state_in[127:120] == 3'b100;
  assign _0253_ = state_in[127:120] == 2'b11;
  assign _0254_ = state_in[127:120] == 2'b10;
  assign _0255_ = state_in[127:120] == 1'b1;
  assign _0256_ = ! state_in[127:120];
  always @(posedge clk)
      \t0.t0.s4.out <= _0257_;
  wire [255:0] fangyuan2;
  assign fangyuan2 = { _0256_, _0255_, _0254_, _0253_, _0252_, _0251_, _0250_, _0249_, _0248_, _0247_, _0246_, _0245_, _0244_, _0243_, _0242_, _0241_, _0240_, _0239_, _0238_, _0237_, _0236_, _0235_, _0234_, _0233_, _0232_, _0231_, _0230_, _0229_, _0228_, _0227_, _0226_, _0225_, _0224_, _0223_, _0222_, _0221_, _0220_, _0219_, _0218_, _0217_, _0216_, _0215_, _0214_, _0213_, _0212_, _0211_, _0210_, _0209_, _0208_, _0207_, _0206_, _0205_, _0204_, _0203_, _0202_, _0201_, _0200_, _0199_, _0198_, _0197_, _0196_, _0195_, _0194_, _0193_, _0192_, _0191_, _0190_, _0189_, _0188_, _0187_, _0186_, _0185_, _0184_, _0183_, _0182_, _0181_, _0180_, _0179_, _0178_, _0177_, _0176_, _0175_, _0174_, _0173_, _0172_, _0171_, _0170_, _0169_, _0168_, _0167_, _0166_, _0165_, _0164_, _0163_, _0162_, _0161_, _0160_, _0159_, _0158_, _0157_, _0156_, _0155_, _0154_, _0153_, _0152_, _0151_, _0150_, _0149_, _0148_, _0147_, _0146_, _0145_, _0144_, _0143_, _0142_, _0141_, _0140_, _0139_, _0138_, _0137_, _0136_, _0135_, _0134_, _0133_, _0132_, _0131_, _0130_, _0129_, _0128_, _0127_, _0126_, _0125_, _0124_, _0123_, _0122_, _0121_, _0120_, _0119_, _0118_, _0117_, _0116_, _0115_, _0114_, _0113_, _0112_, _0111_, _0110_, _0109_, _0108_, _0107_, _0106_, _0105_, _0104_, _0103_, _0102_, _0101_, _0100_, _0099_, _0098_, _0097_, _0096_, _0095_, _0094_, _0093_, _0092_, _0091_, _0090_, _0089_, _0088_, _0087_, _0086_, _0085_, _0084_, _0083_, _0082_, _0081_, _0080_, _0079_, _0078_, _0077_, _0076_, _0075_, _0074_, _0073_, _0072_, _0071_, _0070_, _0069_, _0068_, _0067_, _0066_, _0065_, _0064_, _0063_, _0062_, _0061_, _0060_, _0059_, _0058_, _0057_, _0056_, _0055_, _0054_, _0053_, _0052_, _0051_, _0050_, _0049_, _0048_, _0047_, _0046_, _0045_, _0044_, _0043_, _0042_, _0041_, _0040_, _0039_, _0038_, _0037_, _0036_, _0035_, _0034_, _0033_, _0032_, _0031_, _0030_, _0029_, _0028_, _0027_, _0026_, _0025_, _0024_, _0023_, _0022_, _0021_, _0020_, _0019_, _0018_, _0017_, _0016_, _0015_, _0014_, _0013_, _0012_, _0011_, _0010_, _0009_, _0008_, _0007_, _0006_, _0005_, _0004_, _0003_, _0002_, _0001_ };

  always @(\t0.t0.s4.out or fangyuan2) begin
    casez (fangyuan2)
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1 :
        _0257_ = 8'b00101100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1? :
        _0257_ = 8'b01101101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?? :
        _0257_ = 8'b10101000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??? :
        _0257_ = 8'b01111011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???? :
        _0257_ = 8'b00011110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????? :
        _0257_ = 8'b01011010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????? :
        _0257_ = 8'b00101001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????? :
        _0257_ = 8'b10000010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????? :
        _0257_ = 8'b11010000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????? :
        _0257_ = 8'b10000100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????? :
        _0257_ = 8'b11010111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????? :
        _0257_ = 8'b01100101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????? :
        _0257_ = 8'b00011010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????? :
        _0257_ = 8'b00001001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????? :
        _0257_ = 8'b01011001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????? :
        _0257_ = 8'b00000011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????? :
        _0257_ = 8'b10100101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????? :
        _0257_ = 8'b01010000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????? :
        _0257_ = 8'b10101010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????? :
        _0257_ = 8'b10000111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????? :
        _0257_ = 8'b11001001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????? :
        _0257_ = 8'b00010101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????? :
        _0257_ = 8'b00111100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????? :
        _0257_ = 8'b00101101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????? :
        _0257_ = 8'b00110011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????? :
        _0257_ = 8'b00000111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????? :
        _0257_ = 8'b10101001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????? :
        _0257_ = 8'b11010010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????? :
        _0257_ = 8'b00100010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????? :
        _0257_ = 8'b00101011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????? :
        _0257_ = 8'b11101011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????? :
        _0257_ = 8'b11011001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????? :
        _0257_ = 8'b00100111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????? :
        _0257_ = 8'b00111010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????? :
        _0257_ = 8'b10011001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????? :
        _0257_ = 8'b00010111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????? :
        _0257_ = 8'b01101001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????? :
        _0257_ = 8'b10101110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????? :
        _0257_ = 8'b01101010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????? :
        _0257_ = 8'b11000010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????? :
        _0257_ = 8'b00011100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????? :
        _0257_ = 8'b11110111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????? :
        _0257_ = 8'b00000110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????? :
        _0257_ = 8'b10010000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????? :
        _0257_ = 8'b11001100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????? :
        _0257_ = 8'b01110001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????? :
        _0257_ = 8'b01111100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????? :
        _0257_ = 8'b11100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????? :
        _0257_ = 8'b00001111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????? :
        _0257_ = 8'b00001101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????? :
        _0257_ = 8'b01100001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????? :
        _0257_ = 8'b10010110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????? :
        _0257_ = 8'b00111110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????? :
        _0257_ = 8'b11101000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????? :
        _0257_ = 8'b10100001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????? :
        _0257_ = 8'b11001011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????? :
        _0257_ = 8'b10010111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????? :
        _0257_ = 8'b01110011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????? :
        _0257_ = 8'b01010111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????? :
        _0257_ = 8'b00111000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????? :
        _0257_ = 8'b01011100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????? :
        _0257_ = 8'b01001010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????? :
        _0257_ = 8'b11110000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????? :
        _0257_ = 8'b01101111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????? :
        _0257_ = 8'b00010000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b01000111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b11110100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b11001010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b11001111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b11110011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b10101100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b11011000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b01001001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b10011100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b10110001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b00000001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b11011010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b01101110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b10001011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b11010101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b11110010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b11010011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b00110001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b00111001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b11000100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b01000011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b10111101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b10011111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b10111000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b01001000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b00001100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b10010010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b00010100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b01110100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b01100100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b11011011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b10101101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b00010110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b10111100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b10100111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b00101000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b01101011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b11000111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b10001100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b00001011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b00111011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b01010100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b01000100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b10100011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b10011110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b00011001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b11000000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b11100110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b00110010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b10111010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b11001000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b01111010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b11111100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b01010101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b10010011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b00101110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b10001000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b00110101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b10111110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b11000011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b00100110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b00011000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b10000001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b10111111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b11111101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b11100101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b00100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b01000010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b10101111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b01110111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b01100011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b11110001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b01110000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b00100001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b00111111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b00000101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b10000000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b01011101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b10100010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b01001011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b00100101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b01111000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b10100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b11111110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b00000100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b11101001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b10001010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b00010001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b01100110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b10011010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b10000110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b11101101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b01001111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b11000101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b10111011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b10000101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b10110000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b10011000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b10010100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b01110010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b01100111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b10001101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b11010100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b10110110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b01111001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b11100011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b01000000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b11000001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b00000000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b10111001 ;
      256'b????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b10100110 ;
      256'b???????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b00010011 ;
      256'b??????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b01011110 ;
      256'b?????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b11011101 ;
      256'b????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b01010010 ;
      256'b???????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b01111101 ;
      256'b??????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b10110111 ;
      256'b?????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b01110110 ;
      256'b????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b10100100 ;
      256'b???????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b01011011 ;
      256'b??????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b10110100 ;
      256'b?????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b11011100 ;
      256'b????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b00110110 ;
      256'b???????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b00110100 ;
      256'b??????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b01011000 ;
      256'b?????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b00011101 ;
      256'b????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b00010010 ;
      256'b???????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b11101010 ;
      256'b??????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b01111111 ;
      256'b?????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b01001110 ;
      256'b????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b11001101 ;
      256'b???????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b11011111 ;
      256'b??????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b00011011 ;
      256'b?????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b00100100 ;
      256'b????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b00001110 ;
      256'b???????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b00101111 ;
      256'b??????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b00001010 ;
      256'b?????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b00110111 ;
      256'b????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b00110000 ;
      256'b???????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b10011101 ;
      256'b??????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b01000110 ;
      256'b?????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b10010101 ;
      256'b????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b00001000 ;
      256'b???????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b00101010 ;
      256'b??????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b01100010 ;
      256'b?????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b10101011 ;
      256'b????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b11100010 ;
      256'b???????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b11111001 ;
      256'b??????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b11010001 ;
      256'b?????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b01010001 ;
      256'b????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b01101000 ;
      256'b???????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b10000011 ;
      256'b??????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b11110101 ;
      256'b?????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b01111110 ;
      256'b????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b01101100 ;
      256'b???????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b01001100 ;
      256'b??????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b00111101 ;
      256'b?????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b11100001 ;
      256'b????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b01110101 ;
      256'b???????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b10011011 ;
      256'b??????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b11100100 ;
      256'b?????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b01010011 ;
      256'b????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b00100011 ;
      256'b???????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b01000101 ;
      256'b??????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b01011111 ;
      256'b?????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b10110011 ;
      256'b????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b01000001 ;
      256'b???????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b11111011 ;
      256'b??????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b10001110 ;
      256'b?????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b10110010 ;
      256'b????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b11101111 ;
      256'b???????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b11111010 ;
      256'b??????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b10001001 ;
      256'b?????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b00011111 ;
      256'b????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b10001111 ;
      256'b???????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b11101100 ;
      256'b??????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b01001101 ;
      256'b?????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b10110101 ;
      256'b????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b11100111 ;
      256'b???????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b01010110 ;
      256'b??????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b11001110 ;
      256'b?????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b00000010 ;
      256'b????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b01100000 ;
      256'b???????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b10010001 ;
      256'b??????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b11011110 ;
      256'b?????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b11010110 ;
      256'b????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b11111111 ;
      256'b???1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b11110110 ;
      256'b??1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b11101110 ;
      256'b?1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b11111000 ;
      256'b1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b11000110 ;
      default:
        _0257_ = \t0.t0.s4.out ;
    endcase
  end
  assign p01[31:24] = \t0.t1.s0.out ^ \t0.t1.s4.out ;
  always @(posedge clk)
      \t0.t1.s0.out <= _0258_;
  wire [255:0] fangyuan3;
  assign fangyuan3 = { _0514_, _0513_, _0512_, _0511_, _0510_, _0509_, _0508_, _0507_, _0506_, _0505_, _0504_, _0503_, _0502_, _0501_, _0500_, _0499_, _0498_, _0497_, _0496_, _0495_, _0494_, _0493_, _0492_, _0491_, _0490_, _0489_, _0488_, _0487_, _0486_, _0485_, _0484_, _0483_, _0482_, _0481_, _0480_, _0479_, _0478_, _0477_, _0476_, _0475_, _0474_, _0473_, _0472_, _0471_, _0470_, _0469_, _0468_, _0467_, _0466_, _0465_, _0464_, _0463_, _0462_, _0461_, _0460_, _0459_, _0458_, _0457_, _0456_, _0455_, _0454_, _0453_, _0452_, _0451_, _0450_, _0449_, _0448_, _0447_, _0446_, _0445_, _0444_, _0443_, _0442_, _0441_, _0440_, _0439_, _0438_, _0437_, _0436_, _0435_, _0434_, _0433_, _0432_, _0431_, _0430_, _0429_, _0428_, _0427_, _0426_, _0425_, _0424_, _0423_, _0422_, _0421_, _0420_, _0419_, _0418_, _0417_, _0416_, _0415_, _0414_, _0413_, _0412_, _0411_, _0410_, _0409_, _0408_, _0407_, _0406_, _0405_, _0404_, _0403_, _0402_, _0401_, _0400_, _0399_, _0398_, _0397_, _0396_, _0395_, _0394_, _0393_, _0392_, _0391_, _0390_, _0389_, _0388_, _0387_, _0386_, _0385_, _0384_, _0383_, _0382_, _0381_, _0380_, _0379_, _0378_, _0377_, _0376_, _0375_, _0374_, _0373_, _0372_, _0371_, _0370_, _0369_, _0368_, _0367_, _0366_, _0365_, _0364_, _0363_, _0362_, _0361_, _0360_, _0359_, _0358_, _0357_, _0356_, _0355_, _0354_, _0353_, _0352_, _0351_, _0350_, _0349_, _0348_, _0347_, _0346_, _0345_, _0344_, _0343_, _0342_, _0341_, _0340_, _0339_, _0338_, _0337_, _0336_, _0335_, _0334_, _0333_, _0332_, _0331_, _0330_, _0329_, _0328_, _0327_, _0326_, _0325_, _0324_, _0323_, _0322_, _0321_, _0320_, _0319_, _0318_, _0317_, _0316_, _0315_, _0314_, _0313_, _0312_, _0311_, _0310_, _0309_, _0308_, _0307_, _0306_, _0305_, _0304_, _0303_, _0302_, _0301_, _0300_, _0299_, _0298_, _0297_, _0296_, _0295_, _0294_, _0293_, _0292_, _0291_, _0290_, _0289_, _0288_, _0287_, _0286_, _0285_, _0284_, _0283_, _0282_, _0281_, _0280_, _0279_, _0278_, _0277_, _0276_, _0275_, _0274_, _0273_, _0272_, _0271_, _0270_, _0269_, _0268_, _0267_, _0266_, _0265_, _0264_, _0263_, _0262_, _0261_, _0260_, _0259_ };

  always @(\t0.t1.s0.out or fangyuan3) begin
    casez (fangyuan3)
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1 :
        _0258_ = 8'b00010110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1? :
        _0258_ = 8'b10111011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?? :
        _0258_ = 8'b01010100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??? :
        _0258_ = 8'b10110000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???? :
        _0258_ = 8'b00001111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????? :
        _0258_ = 8'b00101101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????? :
        _0258_ = 8'b10011001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????? :
        _0258_ = 8'b01000001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????? :
        _0258_ = 8'b01101000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????? :
        _0258_ = 8'b01000010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????? :
        _0258_ = 8'b11100110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????? :
        _0258_ = 8'b10111111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????? :
        _0258_ = 8'b00001101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????? :
        _0258_ = 8'b10001001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????? :
        _0258_ = 8'b10100001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????? :
        _0258_ = 8'b10001100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????? :
        _0258_ = 8'b11011111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????? :
        _0258_ = 8'b00101000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????? :
        _0258_ = 8'b01010101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????? :
        _0258_ = 8'b11001110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????? :
        _0258_ = 8'b11101001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????? :
        _0258_ = 8'b10000111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????? :
        _0258_ = 8'b00011110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????? :
        _0258_ = 8'b10011011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????? :
        _0258_ = 8'b10010100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????? :
        _0258_ = 8'b10001110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????? :
        _0258_ = 8'b11011001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????? :
        _0258_ = 8'b01101001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????? :
        _0258_ = 8'b00010001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????? :
        _0258_ = 8'b10011000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????? :
        _0258_ = 8'b11111000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????? :
        _0258_ = 8'b11100001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????? :
        _0258_ = 8'b10011110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????? :
        _0258_ = 8'b00011101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????? :
        _0258_ = 8'b11000001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????? :
        _0258_ = 8'b10000110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????? :
        _0258_ = 8'b10111001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????? :
        _0258_ = 8'b01010111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????? :
        _0258_ = 8'b00110101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????? :
        _0258_ = 8'b01100001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????? :
        _0258_ = 8'b00001110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????? :
        _0258_ = 8'b11110110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????? :
        _0258_ = 8'b00000011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????? :
        _0258_ = 8'b01001000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????? :
        _0258_ = 8'b01100110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????? :
        _0258_ = 8'b10110101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????? :
        _0258_ = 8'b00111110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????? :
        _0258_ = 8'b01110000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????? :
        _0258_ = 8'b10001010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????? :
        _0258_ = 8'b10001011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????? :
        _0258_ = 8'b10111101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????? :
        _0258_ = 8'b01001011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????? :
        _0258_ = 8'b00011111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????? :
        _0258_ = 8'b01110100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????? :
        _0258_ = 8'b11011101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????? :
        _0258_ = 8'b11101000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????? :
        _0258_ = 8'b11000110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????? :
        _0258_ = 8'b10110100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????? :
        _0258_ = 8'b10100110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????? :
        _0258_ = 8'b00011100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????? :
        _0258_ = 8'b00101110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????? :
        _0258_ = 8'b00100101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????? :
        _0258_ = 8'b01111000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????? :
        _0258_ = 8'b10111010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????? :
        _0258_ = 8'b00001000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b10101110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b01111010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b01100101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b11101010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b11110100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b01010110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b01101100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b10101001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b01001110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b11010101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b10001101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b01101101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b00110111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b11001000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b11100111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b01111001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b11100100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b10010101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b10010001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b01100010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b10101100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b11010011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b11000010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b01011100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b00100100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b00000110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b01001001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b00001010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b00111010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b00110010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b11100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b11011011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b00001011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b01011110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b11011110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b00010100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b10111000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b11101110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b01000110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b10001000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b10010000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b00101010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b00100010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b11011100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b01001111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b10000001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b01100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b01110011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b00011001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b01011101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b01100100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b00111101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b01111110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b10100111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b11000100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b00010111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b01000100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b10010111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b01011111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b11101100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b00010011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b00001100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b11001101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b11010010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b11110011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b11111111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b00010000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b00100001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b11011010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b10110110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b10111100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b11110101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b00111000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b10011101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b10010010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b10001111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b01000000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b10100011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b01010001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b10101000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b10011111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b00111100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b01010000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b01111111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b00000010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b11111001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b01000101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b10000101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b00110011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b01001101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b01000011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b11111011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b10101010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b11101111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b11010000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b11001111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b01011000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b01001100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b01001010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b00111001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b10111110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b11001011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b01101010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b01011011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b10110001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b11111100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b00100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b11101101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b00000000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b11010001 ;
      256'b????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b01010011 ;
      256'b???????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b10000100 ;
      256'b??????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b00101111 ;
      256'b?????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b11100011 ;
      256'b????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b00101001 ;
      256'b???????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b10110011 ;
      256'b??????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b11010110 ;
      256'b?????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b00111011 ;
      256'b????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b01010010 ;
      256'b???????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b10100000 ;
      256'b??????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b01011010 ;
      256'b?????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b01101110 ;
      256'b????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b00011011 ;
      256'b???????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b00011010 ;
      256'b??????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b00101100 ;
      256'b?????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b10000011 ;
      256'b????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b00001001 ;
      256'b???????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b01110101 ;
      256'b??????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b10110010 ;
      256'b?????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b00100111 ;
      256'b????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b11101011 ;
      256'b???????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b11100010 ;
      256'b??????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b10000000 ;
      256'b?????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b00010010 ;
      256'b????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b00000111 ;
      256'b???????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b10011010 ;
      256'b??????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b00000101 ;
      256'b?????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b10010110 ;
      256'b????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b00011000 ;
      256'b???????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b11000011 ;
      256'b??????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b00100011 ;
      256'b?????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b11000111 ;
      256'b????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b00000100 ;
      256'b???????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b00010101 ;
      256'b??????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b00110001 ;
      256'b?????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b11011000 ;
      256'b????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b01110001 ;
      256'b???????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b11110001 ;
      256'b??????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b11100101 ;
      256'b?????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b10100101 ;
      256'b????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b00110100 ;
      256'b???????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b11001100 ;
      256'b??????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b11110111 ;
      256'b?????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b00111111 ;
      256'b????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b00110110 ;
      256'b???????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b00100110 ;
      256'b??????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b10010011 ;
      256'b?????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b11111101 ;
      256'b????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b10110111 ;
      256'b???????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b11000000 ;
      256'b??????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b01110010 ;
      256'b?????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b10100100 ;
      256'b????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b10011100 ;
      256'b???????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b10101111 ;
      256'b??????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b10100010 ;
      256'b?????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b11010100 ;
      256'b????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b10101101 ;
      256'b???????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b11110000 ;
      256'b??????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b01000111 ;
      256'b?????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b01011001 ;
      256'b????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b11111010 ;
      256'b???????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b01111101 ;
      256'b??????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b11001001 ;
      256'b?????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b10000010 ;
      256'b????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b11001010 ;
      256'b???????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b01110110 ;
      256'b??????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b10101011 ;
      256'b?????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b11010111 ;
      256'b????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b11111110 ;
      256'b???????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b00101011 ;
      256'b??????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b01100111 ;
      256'b?????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b00000001 ;
      256'b????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b00110000 ;
      256'b???????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b11000101 ;
      256'b??????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b01101111 ;
      256'b?????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b01101011 ;
      256'b????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b11110010 ;
      256'b???1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b01111011 ;
      256'b??1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b01110111 ;
      256'b?1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b01111100 ;
      256'b1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b01100011 ;
      default:
        _0258_ = \t0.t1.s0.out ;
    endcase
  end
  assign _0259_ = state_in[119:112] == 8'b11111111;
  assign _0260_ = state_in[119:112] == 8'b11111110;
  assign _0261_ = state_in[119:112] == 8'b11111101;
  assign _0262_ = state_in[119:112] == 8'b11111100;
  assign _0263_ = state_in[119:112] == 8'b11111011;
  assign _0264_ = state_in[119:112] == 8'b11111010;
  assign _0265_ = state_in[119:112] == 8'b11111001;
  assign _0266_ = state_in[119:112] == 8'b11111000;
  assign _0267_ = state_in[119:112] == 8'b11110111;
  assign _0268_ = state_in[119:112] == 8'b11110110;
  assign _0269_ = state_in[119:112] == 8'b11110101;
  assign _0270_ = state_in[119:112] == 8'b11110100;
  assign _0271_ = state_in[119:112] == 8'b11110011;
  assign _0272_ = state_in[119:112] == 8'b11110010;
  assign _0273_ = state_in[119:112] == 8'b11110001;
  assign _0274_ = state_in[119:112] == 8'b11110000;
  assign _0275_ = state_in[119:112] == 8'b11101111;
  assign _0276_ = state_in[119:112] == 8'b11101110;
  assign _0277_ = state_in[119:112] == 8'b11101101;
  assign _0278_ = state_in[119:112] == 8'b11101100;
  assign _0279_ = state_in[119:112] == 8'b11101011;
  assign _0280_ = state_in[119:112] == 8'b11101010;
  assign _0281_ = state_in[119:112] == 8'b11101001;
  assign _0282_ = state_in[119:112] == 8'b11101000;
  assign _0283_ = state_in[119:112] == 8'b11100111;
  assign _0284_ = state_in[119:112] == 8'b11100110;
  assign _0285_ = state_in[119:112] == 8'b11100101;
  assign _0286_ = state_in[119:112] == 8'b11100100;
  assign _0287_ = state_in[119:112] == 8'b11100011;
  assign _0288_ = state_in[119:112] == 8'b11100010;
  assign _0289_ = state_in[119:112] == 8'b11100001;
  assign _0290_ = state_in[119:112] == 8'b11100000;
  assign _0291_ = state_in[119:112] == 8'b11011111;
  assign _0292_ = state_in[119:112] == 8'b11011110;
  assign _0293_ = state_in[119:112] == 8'b11011101;
  assign _0294_ = state_in[119:112] == 8'b11011100;
  assign _0295_ = state_in[119:112] == 8'b11011011;
  assign _0296_ = state_in[119:112] == 8'b11011010;
  assign _0297_ = state_in[119:112] == 8'b11011001;
  assign _0298_ = state_in[119:112] == 8'b11011000;
  assign _0299_ = state_in[119:112] == 8'b11010111;
  assign _0300_ = state_in[119:112] == 8'b11010110;
  assign _0301_ = state_in[119:112] == 8'b11010101;
  assign _0302_ = state_in[119:112] == 8'b11010100;
  assign _0303_ = state_in[119:112] == 8'b11010011;
  assign _0304_ = state_in[119:112] == 8'b11010010;
  assign _0305_ = state_in[119:112] == 8'b11010001;
  assign _0306_ = state_in[119:112] == 8'b11010000;
  assign _0307_ = state_in[119:112] == 8'b11001111;
  assign _0308_ = state_in[119:112] == 8'b11001110;
  assign _0309_ = state_in[119:112] == 8'b11001101;
  assign _0310_ = state_in[119:112] == 8'b11001100;
  assign _0311_ = state_in[119:112] == 8'b11001011;
  assign _0312_ = state_in[119:112] == 8'b11001010;
  assign _0313_ = state_in[119:112] == 8'b11001001;
  assign _0314_ = state_in[119:112] == 8'b11001000;
  assign _0315_ = state_in[119:112] == 8'b11000111;
  assign _0316_ = state_in[119:112] == 8'b11000110;
  assign _0317_ = state_in[119:112] == 8'b11000101;
  assign _0318_ = state_in[119:112] == 8'b11000100;
  assign _0319_ = state_in[119:112] == 8'b11000011;
  assign _0320_ = state_in[119:112] == 8'b11000010;
  assign _0321_ = state_in[119:112] == 8'b11000001;
  assign _0322_ = state_in[119:112] == 8'b11000000;
  assign _0323_ = state_in[119:112] == 8'b10111111;
  assign _0324_ = state_in[119:112] == 8'b10111110;
  assign _0325_ = state_in[119:112] == 8'b10111101;
  assign _0326_ = state_in[119:112] == 8'b10111100;
  assign _0327_ = state_in[119:112] == 8'b10111011;
  assign _0328_ = state_in[119:112] == 8'b10111010;
  assign _0329_ = state_in[119:112] == 8'b10111001;
  assign _0330_ = state_in[119:112] == 8'b10111000;
  assign _0331_ = state_in[119:112] == 8'b10110111;
  assign _0332_ = state_in[119:112] == 8'b10110110;
  assign _0333_ = state_in[119:112] == 8'b10110101;
  assign _0334_ = state_in[119:112] == 8'b10110100;
  assign _0335_ = state_in[119:112] == 8'b10110011;
  assign _0336_ = state_in[119:112] == 8'b10110010;
  assign _0337_ = state_in[119:112] == 8'b10110001;
  assign _0338_ = state_in[119:112] == 8'b10110000;
  assign _0339_ = state_in[119:112] == 8'b10101111;
  assign _0340_ = state_in[119:112] == 8'b10101110;
  assign _0341_ = state_in[119:112] == 8'b10101101;
  assign _0342_ = state_in[119:112] == 8'b10101100;
  assign _0343_ = state_in[119:112] == 8'b10101011;
  assign _0344_ = state_in[119:112] == 8'b10101010;
  assign _0345_ = state_in[119:112] == 8'b10101001;
  assign _0346_ = state_in[119:112] == 8'b10101000;
  assign _0347_ = state_in[119:112] == 8'b10100111;
  assign _0348_ = state_in[119:112] == 8'b10100110;
  assign _0349_ = state_in[119:112] == 8'b10100101;
  assign _0350_ = state_in[119:112] == 8'b10100100;
  assign _0351_ = state_in[119:112] == 8'b10100011;
  assign _0352_ = state_in[119:112] == 8'b10100010;
  assign _0353_ = state_in[119:112] == 8'b10100001;
  assign _0354_ = state_in[119:112] == 8'b10100000;
  assign _0355_ = state_in[119:112] == 8'b10011111;
  assign _0356_ = state_in[119:112] == 8'b10011110;
  assign _0357_ = state_in[119:112] == 8'b10011101;
  assign _0358_ = state_in[119:112] == 8'b10011100;
  assign _0359_ = state_in[119:112] == 8'b10011011;
  assign _0360_ = state_in[119:112] == 8'b10011010;
  assign _0361_ = state_in[119:112] == 8'b10011001;
  assign _0362_ = state_in[119:112] == 8'b10011000;
  assign _0363_ = state_in[119:112] == 8'b10010111;
  assign _0364_ = state_in[119:112] == 8'b10010110;
  assign _0365_ = state_in[119:112] == 8'b10010101;
  assign _0366_ = state_in[119:112] == 8'b10010100;
  assign _0367_ = state_in[119:112] == 8'b10010011;
  assign _0368_ = state_in[119:112] == 8'b10010010;
  assign _0369_ = state_in[119:112] == 8'b10010001;
  assign _0370_ = state_in[119:112] == 8'b10010000;
  assign _0371_ = state_in[119:112] == 8'b10001111;
  assign _0372_ = state_in[119:112] == 8'b10001110;
  assign _0373_ = state_in[119:112] == 8'b10001101;
  assign _0374_ = state_in[119:112] == 8'b10001100;
  assign _0375_ = state_in[119:112] == 8'b10001011;
  assign _0376_ = state_in[119:112] == 8'b10001010;
  assign _0377_ = state_in[119:112] == 8'b10001001;
  assign _0378_ = state_in[119:112] == 8'b10001000;
  assign _0379_ = state_in[119:112] == 8'b10000111;
  assign _0380_ = state_in[119:112] == 8'b10000110;
  assign _0381_ = state_in[119:112] == 8'b10000101;
  assign _0382_ = state_in[119:112] == 8'b10000100;
  assign _0383_ = state_in[119:112] == 8'b10000011;
  assign _0384_ = state_in[119:112] == 8'b10000010;
  assign _0385_ = state_in[119:112] == 8'b10000001;
  assign _0386_ = state_in[119:112] == 8'b10000000;
  assign _0387_ = state_in[119:112] == 7'b1111111;
  assign _0388_ = state_in[119:112] == 7'b1111110;
  assign _0389_ = state_in[119:112] == 7'b1111101;
  assign _0390_ = state_in[119:112] == 7'b1111100;
  assign _0391_ = state_in[119:112] == 7'b1111011;
  assign _0392_ = state_in[119:112] == 7'b1111010;
  assign _0393_ = state_in[119:112] == 7'b1111001;
  assign _0394_ = state_in[119:112] == 7'b1111000;
  assign _0395_ = state_in[119:112] == 7'b1110111;
  assign _0396_ = state_in[119:112] == 7'b1110110;
  assign _0397_ = state_in[119:112] == 7'b1110101;
  assign _0398_ = state_in[119:112] == 7'b1110100;
  assign _0399_ = state_in[119:112] == 7'b1110011;
  assign _0400_ = state_in[119:112] == 7'b1110010;
  assign _0401_ = state_in[119:112] == 7'b1110001;
  assign _0402_ = state_in[119:112] == 7'b1110000;
  assign _0403_ = state_in[119:112] == 7'b1101111;
  assign _0404_ = state_in[119:112] == 7'b1101110;
  assign _0405_ = state_in[119:112] == 7'b1101101;
  assign _0406_ = state_in[119:112] == 7'b1101100;
  assign _0407_ = state_in[119:112] == 7'b1101011;
  assign _0408_ = state_in[119:112] == 7'b1101010;
  assign _0409_ = state_in[119:112] == 7'b1101001;
  assign _0410_ = state_in[119:112] == 7'b1101000;
  assign _0411_ = state_in[119:112] == 7'b1100111;
  assign _0412_ = state_in[119:112] == 7'b1100110;
  assign _0413_ = state_in[119:112] == 7'b1100101;
  assign _0414_ = state_in[119:112] == 7'b1100100;
  assign _0415_ = state_in[119:112] == 7'b1100011;
  assign _0416_ = state_in[119:112] == 7'b1100010;
  assign _0417_ = state_in[119:112] == 7'b1100001;
  assign _0418_ = state_in[119:112] == 7'b1100000;
  assign _0419_ = state_in[119:112] == 7'b1011111;
  assign _0420_ = state_in[119:112] == 7'b1011110;
  assign _0421_ = state_in[119:112] == 7'b1011101;
  assign _0422_ = state_in[119:112] == 7'b1011100;
  assign _0423_ = state_in[119:112] == 7'b1011011;
  assign _0424_ = state_in[119:112] == 7'b1011010;
  assign _0425_ = state_in[119:112] == 7'b1011001;
  assign _0426_ = state_in[119:112] == 7'b1011000;
  assign _0427_ = state_in[119:112] == 7'b1010111;
  assign _0428_ = state_in[119:112] == 7'b1010110;
  assign _0429_ = state_in[119:112] == 7'b1010101;
  assign _0430_ = state_in[119:112] == 7'b1010100;
  assign _0431_ = state_in[119:112] == 7'b1010011;
  assign _0432_ = state_in[119:112] == 7'b1010010;
  assign _0433_ = state_in[119:112] == 7'b1010001;
  assign _0434_ = state_in[119:112] == 7'b1010000;
  assign _0435_ = state_in[119:112] == 7'b1001111;
  assign _0436_ = state_in[119:112] == 7'b1001110;
  assign _0437_ = state_in[119:112] == 7'b1001101;
  assign _0438_ = state_in[119:112] == 7'b1001100;
  assign _0439_ = state_in[119:112] == 7'b1001011;
  assign _0440_ = state_in[119:112] == 7'b1001010;
  assign _0441_ = state_in[119:112] == 7'b1001001;
  assign _0442_ = state_in[119:112] == 7'b1001000;
  assign _0443_ = state_in[119:112] == 7'b1000111;
  assign _0444_ = state_in[119:112] == 7'b1000110;
  assign _0445_ = state_in[119:112] == 7'b1000101;
  assign _0446_ = state_in[119:112] == 7'b1000100;
  assign _0447_ = state_in[119:112] == 7'b1000011;
  assign _0448_ = state_in[119:112] == 7'b1000010;
  assign _0449_ = state_in[119:112] == 7'b1000001;
  assign _0450_ = state_in[119:112] == 7'b1000000;
  assign _0451_ = state_in[119:112] == 6'b111111;
  assign _0452_ = state_in[119:112] == 6'b111110;
  assign _0453_ = state_in[119:112] == 6'b111101;
  assign _0454_ = state_in[119:112] == 6'b111100;
  assign _0455_ = state_in[119:112] == 6'b111011;
  assign _0456_ = state_in[119:112] == 6'b111010;
  assign _0457_ = state_in[119:112] == 6'b111001;
  assign _0458_ = state_in[119:112] == 6'b111000;
  assign _0459_ = state_in[119:112] == 6'b110111;
  assign _0460_ = state_in[119:112] == 6'b110110;
  assign _0461_ = state_in[119:112] == 6'b110101;
  assign _0462_ = state_in[119:112] == 6'b110100;
  assign _0463_ = state_in[119:112] == 6'b110011;
  assign _0464_ = state_in[119:112] == 6'b110010;
  assign _0465_ = state_in[119:112] == 6'b110001;
  assign _0466_ = state_in[119:112] == 6'b110000;
  assign _0467_ = state_in[119:112] == 6'b101111;
  assign _0468_ = state_in[119:112] == 6'b101110;
  assign _0469_ = state_in[119:112] == 6'b101101;
  assign _0470_ = state_in[119:112] == 6'b101100;
  assign _0471_ = state_in[119:112] == 6'b101011;
  assign _0472_ = state_in[119:112] == 6'b101010;
  assign _0473_ = state_in[119:112] == 6'b101001;
  assign _0474_ = state_in[119:112] == 6'b101000;
  assign _0475_ = state_in[119:112] == 6'b100111;
  assign _0476_ = state_in[119:112] == 6'b100110;
  assign _0477_ = state_in[119:112] == 6'b100101;
  assign _0478_ = state_in[119:112] == 6'b100100;
  assign _0479_ = state_in[119:112] == 6'b100011;
  assign _0480_ = state_in[119:112] == 6'b100010;
  assign _0481_ = state_in[119:112] == 6'b100001;
  assign _0482_ = state_in[119:112] == 6'b100000;
  assign _0483_ = state_in[119:112] == 5'b11111;
  assign _0484_ = state_in[119:112] == 5'b11110;
  assign _0485_ = state_in[119:112] == 5'b11101;
  assign _0486_ = state_in[119:112] == 5'b11100;
  assign _0487_ = state_in[119:112] == 5'b11011;
  assign _0488_ = state_in[119:112] == 5'b11010;
  assign _0489_ = state_in[119:112] == 5'b11001;
  assign _0490_ = state_in[119:112] == 5'b11000;
  assign _0491_ = state_in[119:112] == 5'b10111;
  assign _0492_ = state_in[119:112] == 5'b10110;
  assign _0493_ = state_in[119:112] == 5'b10101;
  assign _0494_ = state_in[119:112] == 5'b10100;
  assign _0495_ = state_in[119:112] == 5'b10011;
  assign _0496_ = state_in[119:112] == 5'b10010;
  assign _0497_ = state_in[119:112] == 5'b10001;
  assign _0498_ = state_in[119:112] == 5'b10000;
  assign _0499_ = state_in[119:112] == 4'b1111;
  assign _0500_ = state_in[119:112] == 4'b1110;
  assign _0501_ = state_in[119:112] == 4'b1101;
  assign _0502_ = state_in[119:112] == 4'b1100;
  assign _0503_ = state_in[119:112] == 4'b1011;
  assign _0504_ = state_in[119:112] == 4'b1010;
  assign _0505_ = state_in[119:112] == 4'b1001;
  assign _0506_ = state_in[119:112] == 4'b1000;
  assign _0507_ = state_in[119:112] == 3'b111;
  assign _0508_ = state_in[119:112] == 3'b110;
  assign _0509_ = state_in[119:112] == 3'b101;
  assign _0510_ = state_in[119:112] == 3'b100;
  assign _0511_ = state_in[119:112] == 2'b11;
  assign _0512_ = state_in[119:112] == 2'b10;
  assign _0513_ = state_in[119:112] == 1'b1;
  assign _0514_ = ! state_in[119:112];
  always @(posedge clk)
      \t0.t1.s4.out <= _0515_;
  wire [255:0] fangyuan4;
  assign fangyuan4 = { _0514_, _0513_, _0512_, _0511_, _0510_, _0509_, _0508_, _0507_, _0506_, _0505_, _0504_, _0503_, _0502_, _0501_, _0500_, _0499_, _0498_, _0497_, _0496_, _0495_, _0494_, _0493_, _0492_, _0491_, _0490_, _0489_, _0488_, _0487_, _0486_, _0485_, _0484_, _0483_, _0482_, _0481_, _0480_, _0479_, _0478_, _0477_, _0476_, _0475_, _0474_, _0473_, _0472_, _0471_, _0470_, _0469_, _0468_, _0467_, _0466_, _0465_, _0464_, _0463_, _0462_, _0461_, _0460_, _0459_, _0458_, _0457_, _0456_, _0455_, _0454_, _0453_, _0452_, _0451_, _0450_, _0449_, _0448_, _0447_, _0446_, _0445_, _0444_, _0443_, _0442_, _0441_, _0440_, _0439_, _0438_, _0437_, _0436_, _0435_, _0434_, _0433_, _0432_, _0431_, _0430_, _0429_, _0428_, _0427_, _0426_, _0425_, _0424_, _0423_, _0422_, _0421_, _0420_, _0419_, _0418_, _0417_, _0416_, _0415_, _0414_, _0413_, _0412_, _0411_, _0410_, _0409_, _0408_, _0407_, _0406_, _0405_, _0404_, _0403_, _0402_, _0401_, _0400_, _0399_, _0398_, _0397_, _0396_, _0395_, _0394_, _0393_, _0392_, _0391_, _0390_, _0389_, _0388_, _0387_, _0386_, _0385_, _0384_, _0383_, _0382_, _0381_, _0380_, _0379_, _0378_, _0377_, _0376_, _0375_, _0374_, _0373_, _0372_, _0371_, _0370_, _0369_, _0368_, _0367_, _0366_, _0365_, _0364_, _0363_, _0362_, _0361_, _0360_, _0359_, _0358_, _0357_, _0356_, _0355_, _0354_, _0353_, _0352_, _0351_, _0350_, _0349_, _0348_, _0347_, _0346_, _0345_, _0344_, _0343_, _0342_, _0341_, _0340_, _0339_, _0338_, _0337_, _0336_, _0335_, _0334_, _0333_, _0332_, _0331_, _0330_, _0329_, _0328_, _0327_, _0326_, _0325_, _0324_, _0323_, _0322_, _0321_, _0320_, _0319_, _0318_, _0317_, _0316_, _0315_, _0314_, _0313_, _0312_, _0311_, _0310_, _0309_, _0308_, _0307_, _0306_, _0305_, _0304_, _0303_, _0302_, _0301_, _0300_, _0299_, _0298_, _0297_, _0296_, _0295_, _0294_, _0293_, _0292_, _0291_, _0290_, _0289_, _0288_, _0287_, _0286_, _0285_, _0284_, _0283_, _0282_, _0281_, _0280_, _0279_, _0278_, _0277_, _0276_, _0275_, _0274_, _0273_, _0272_, _0271_, _0270_, _0269_, _0268_, _0267_, _0266_, _0265_, _0264_, _0263_, _0262_, _0261_, _0260_, _0259_ };

  always @(\t0.t1.s4.out or fangyuan4) begin
    casez (fangyuan4)
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1 :
        _0515_ = 8'b00101100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1? :
        _0515_ = 8'b01101101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?? :
        _0515_ = 8'b10101000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??? :
        _0515_ = 8'b01111011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???? :
        _0515_ = 8'b00011110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????? :
        _0515_ = 8'b01011010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????? :
        _0515_ = 8'b00101001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????? :
        _0515_ = 8'b10000010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????? :
        _0515_ = 8'b11010000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????? :
        _0515_ = 8'b10000100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????? :
        _0515_ = 8'b11010111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????? :
        _0515_ = 8'b01100101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????? :
        _0515_ = 8'b00011010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????? :
        _0515_ = 8'b00001001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????? :
        _0515_ = 8'b01011001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????? :
        _0515_ = 8'b00000011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????? :
        _0515_ = 8'b10100101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????? :
        _0515_ = 8'b01010000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????? :
        _0515_ = 8'b10101010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????? :
        _0515_ = 8'b10000111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????? :
        _0515_ = 8'b11001001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????? :
        _0515_ = 8'b00010101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????? :
        _0515_ = 8'b00111100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????? :
        _0515_ = 8'b00101101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????? :
        _0515_ = 8'b00110011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????? :
        _0515_ = 8'b00000111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????? :
        _0515_ = 8'b10101001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????? :
        _0515_ = 8'b11010010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????? :
        _0515_ = 8'b00100010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????? :
        _0515_ = 8'b00101011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????? :
        _0515_ = 8'b11101011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????? :
        _0515_ = 8'b11011001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????? :
        _0515_ = 8'b00100111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????? :
        _0515_ = 8'b00111010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????? :
        _0515_ = 8'b10011001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????? :
        _0515_ = 8'b00010111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????? :
        _0515_ = 8'b01101001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????? :
        _0515_ = 8'b10101110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????? :
        _0515_ = 8'b01101010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????? :
        _0515_ = 8'b11000010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????? :
        _0515_ = 8'b00011100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????? :
        _0515_ = 8'b11110111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????? :
        _0515_ = 8'b00000110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????? :
        _0515_ = 8'b10010000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????? :
        _0515_ = 8'b11001100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????? :
        _0515_ = 8'b01110001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????? :
        _0515_ = 8'b01111100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????? :
        _0515_ = 8'b11100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????? :
        _0515_ = 8'b00001111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????? :
        _0515_ = 8'b00001101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????? :
        _0515_ = 8'b01100001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????? :
        _0515_ = 8'b10010110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????? :
        _0515_ = 8'b00111110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????? :
        _0515_ = 8'b11101000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????? :
        _0515_ = 8'b10100001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????? :
        _0515_ = 8'b11001011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????? :
        _0515_ = 8'b10010111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????? :
        _0515_ = 8'b01110011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????? :
        _0515_ = 8'b01010111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????? :
        _0515_ = 8'b00111000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????? :
        _0515_ = 8'b01011100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????? :
        _0515_ = 8'b01001010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????? :
        _0515_ = 8'b11110000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????? :
        _0515_ = 8'b01101111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????? :
        _0515_ = 8'b00010000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b01000111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b11110100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b11001010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b11001111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b11110011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b10101100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b11011000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b01001001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b10011100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b10110001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b00000001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b11011010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b01101110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b10001011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b11010101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b11110010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b11010011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b00110001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b00111001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b11000100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b01000011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b10111101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b10011111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b10111000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b01001000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b00001100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b10010010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b00010100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b01110100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b01100100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b11011011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b10101101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b00010110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b10111100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b10100111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b00101000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b01101011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b11000111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b10001100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b00001011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b00111011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b01010100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b01000100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b10100011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b10011110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b00011001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b11000000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b11100110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b00110010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b10111010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b11001000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b01111010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b11111100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b01010101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b10010011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b00101110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b10001000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b00110101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b10111110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b11000011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b00100110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b00011000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b10000001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b10111111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b11111101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b11100101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b00100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b01000010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b10101111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b01110111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b01100011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b11110001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b01110000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b00100001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b00111111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b00000101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b10000000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b01011101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b10100010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b01001011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b00100101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b01111000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b10100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b11111110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b00000100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b11101001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b10001010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b00010001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b01100110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b10011010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b10000110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b11101101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b01001111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b11000101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b10111011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b10000101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b10110000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b10011000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b10010100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b01110010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b01100111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b10001101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b11010100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b10110110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b01111001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b11100011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b01000000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b11000001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b00000000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b10111001 ;
      256'b????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b10100110 ;
      256'b???????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b00010011 ;
      256'b??????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b01011110 ;
      256'b?????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b11011101 ;
      256'b????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b01010010 ;
      256'b???????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b01111101 ;
      256'b??????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b10110111 ;
      256'b?????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b01110110 ;
      256'b????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b10100100 ;
      256'b???????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b01011011 ;
      256'b??????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b10110100 ;
      256'b?????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b11011100 ;
      256'b????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b00110110 ;
      256'b???????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b00110100 ;
      256'b??????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b01011000 ;
      256'b?????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b00011101 ;
      256'b????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b00010010 ;
      256'b???????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b11101010 ;
      256'b??????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b01111111 ;
      256'b?????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b01001110 ;
      256'b????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b11001101 ;
      256'b???????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b11011111 ;
      256'b??????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b00011011 ;
      256'b?????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b00100100 ;
      256'b????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b00001110 ;
      256'b???????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b00101111 ;
      256'b??????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b00001010 ;
      256'b?????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b00110111 ;
      256'b????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b00110000 ;
      256'b???????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b10011101 ;
      256'b??????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b01000110 ;
      256'b?????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b10010101 ;
      256'b????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b00001000 ;
      256'b???????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b00101010 ;
      256'b??????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b01100010 ;
      256'b?????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b10101011 ;
      256'b????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b11100010 ;
      256'b???????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b11111001 ;
      256'b??????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b11010001 ;
      256'b?????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b01010001 ;
      256'b????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b01101000 ;
      256'b???????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b10000011 ;
      256'b??????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b11110101 ;
      256'b?????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b01111110 ;
      256'b????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b01101100 ;
      256'b???????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b01001100 ;
      256'b??????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b00111101 ;
      256'b?????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b11100001 ;
      256'b????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b01110101 ;
      256'b???????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b10011011 ;
      256'b??????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b11100100 ;
      256'b?????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b01010011 ;
      256'b????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b00100011 ;
      256'b???????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b01000101 ;
      256'b??????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b01011111 ;
      256'b?????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b10110011 ;
      256'b????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b01000001 ;
      256'b???????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b11111011 ;
      256'b??????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b10001110 ;
      256'b?????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b10110010 ;
      256'b????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b11101111 ;
      256'b???????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b11111010 ;
      256'b??????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b10001001 ;
      256'b?????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b00011111 ;
      256'b????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b10001111 ;
      256'b???????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b11101100 ;
      256'b??????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b01001101 ;
      256'b?????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b10110101 ;
      256'b????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b11100111 ;
      256'b???????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b01010110 ;
      256'b??????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b11001110 ;
      256'b?????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b00000010 ;
      256'b????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b01100000 ;
      256'b???????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b10010001 ;
      256'b??????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b11011110 ;
      256'b?????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b11010110 ;
      256'b????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b11111111 ;
      256'b???1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b11110110 ;
      256'b??1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b11101110 ;
      256'b?1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b11111000 ;
      256'b1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b11000110 ;
      default:
        _0515_ = \t0.t1.s4.out ;
    endcase
  end
  assign p02[23:16] = \t0.t2.s0.out ^ \t0.t2.s4.out ;
  always @(posedge clk)
      \t0.t2.s0.out <= _0516_;
  wire [255:0] fangyuan5;
  assign fangyuan5 = { _0772_, _0771_, _0770_, _0769_, _0768_, _0767_, _0766_, _0765_, _0764_, _0763_, _0762_, _0761_, _0760_, _0759_, _0758_, _0757_, _0756_, _0755_, _0754_, _0753_, _0752_, _0751_, _0750_, _0749_, _0748_, _0747_, _0746_, _0745_, _0744_, _0743_, _0742_, _0741_, _0740_, _0739_, _0738_, _0737_, _0736_, _0735_, _0734_, _0733_, _0732_, _0731_, _0730_, _0729_, _0728_, _0727_, _0726_, _0725_, _0724_, _0723_, _0722_, _0721_, _0720_, _0719_, _0718_, _0717_, _0716_, _0715_, _0714_, _0713_, _0712_, _0711_, _0710_, _0709_, _0708_, _0707_, _0706_, _0705_, _0704_, _0703_, _0702_, _0701_, _0700_, _0699_, _0698_, _0697_, _0696_, _0695_, _0694_, _0693_, _0692_, _0691_, _0690_, _0689_, _0688_, _0687_, _0686_, _0685_, _0684_, _0683_, _0682_, _0681_, _0680_, _0679_, _0678_, _0677_, _0676_, _0675_, _0674_, _0673_, _0672_, _0671_, _0670_, _0669_, _0668_, _0667_, _0666_, _0665_, _0664_, _0663_, _0662_, _0661_, _0660_, _0659_, _0658_, _0657_, _0656_, _0655_, _0654_, _0653_, _0652_, _0651_, _0650_, _0649_, _0648_, _0647_, _0646_, _0645_, _0644_, _0643_, _0642_, _0641_, _0640_, _0639_, _0638_, _0637_, _0636_, _0635_, _0634_, _0633_, _0632_, _0631_, _0630_, _0629_, _0628_, _0627_, _0626_, _0625_, _0624_, _0623_, _0622_, _0621_, _0620_, _0619_, _0618_, _0617_, _0616_, _0615_, _0614_, _0613_, _0612_, _0611_, _0610_, _0609_, _0608_, _0607_, _0606_, _0605_, _0604_, _0603_, _0602_, _0601_, _0600_, _0599_, _0598_, _0597_, _0596_, _0595_, _0594_, _0593_, _0592_, _0591_, _0590_, _0589_, _0588_, _0587_, _0586_, _0585_, _0584_, _0583_, _0582_, _0581_, _0580_, _0579_, _0578_, _0577_, _0576_, _0575_, _0574_, _0573_, _0572_, _0571_, _0570_, _0569_, _0568_, _0567_, _0566_, _0565_, _0564_, _0563_, _0562_, _0561_, _0560_, _0559_, _0558_, _0557_, _0556_, _0555_, _0554_, _0553_, _0552_, _0551_, _0550_, _0549_, _0548_, _0547_, _0546_, _0545_, _0544_, _0543_, _0542_, _0541_, _0540_, _0539_, _0538_, _0537_, _0536_, _0535_, _0534_, _0533_, _0532_, _0531_, _0530_, _0529_, _0528_, _0527_, _0526_, _0525_, _0524_, _0523_, _0522_, _0521_, _0520_, _0519_, _0518_, _0517_ };

  always @(\t0.t2.s0.out or fangyuan5) begin
    casez (fangyuan5)
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1 :
        _0516_ = 8'b00010110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1? :
        _0516_ = 8'b10111011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?? :
        _0516_ = 8'b01010100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??? :
        _0516_ = 8'b10110000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???? :
        _0516_ = 8'b00001111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????? :
        _0516_ = 8'b00101101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????? :
        _0516_ = 8'b10011001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????? :
        _0516_ = 8'b01000001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????? :
        _0516_ = 8'b01101000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????? :
        _0516_ = 8'b01000010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????? :
        _0516_ = 8'b11100110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????? :
        _0516_ = 8'b10111111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????? :
        _0516_ = 8'b00001101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????? :
        _0516_ = 8'b10001001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????? :
        _0516_ = 8'b10100001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????? :
        _0516_ = 8'b10001100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????? :
        _0516_ = 8'b11011111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????? :
        _0516_ = 8'b00101000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????? :
        _0516_ = 8'b01010101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????? :
        _0516_ = 8'b11001110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????? :
        _0516_ = 8'b11101001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????? :
        _0516_ = 8'b10000111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????? :
        _0516_ = 8'b00011110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????? :
        _0516_ = 8'b10011011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????? :
        _0516_ = 8'b10010100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????? :
        _0516_ = 8'b10001110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????? :
        _0516_ = 8'b11011001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????? :
        _0516_ = 8'b01101001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????? :
        _0516_ = 8'b00010001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????? :
        _0516_ = 8'b10011000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????? :
        _0516_ = 8'b11111000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????? :
        _0516_ = 8'b11100001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????? :
        _0516_ = 8'b10011110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????? :
        _0516_ = 8'b00011101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????? :
        _0516_ = 8'b11000001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????? :
        _0516_ = 8'b10000110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????? :
        _0516_ = 8'b10111001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????? :
        _0516_ = 8'b01010111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????? :
        _0516_ = 8'b00110101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????? :
        _0516_ = 8'b01100001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????? :
        _0516_ = 8'b00001110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????? :
        _0516_ = 8'b11110110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????? :
        _0516_ = 8'b00000011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????? :
        _0516_ = 8'b01001000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????? :
        _0516_ = 8'b01100110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????? :
        _0516_ = 8'b10110101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????? :
        _0516_ = 8'b00111110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????? :
        _0516_ = 8'b01110000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????? :
        _0516_ = 8'b10001010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????? :
        _0516_ = 8'b10001011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????? :
        _0516_ = 8'b10111101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????? :
        _0516_ = 8'b01001011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????? :
        _0516_ = 8'b00011111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????? :
        _0516_ = 8'b01110100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????? :
        _0516_ = 8'b11011101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????? :
        _0516_ = 8'b11101000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????? :
        _0516_ = 8'b11000110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????? :
        _0516_ = 8'b10110100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????? :
        _0516_ = 8'b10100110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????? :
        _0516_ = 8'b00011100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????? :
        _0516_ = 8'b00101110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????? :
        _0516_ = 8'b00100101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????? :
        _0516_ = 8'b01111000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????? :
        _0516_ = 8'b10111010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????? :
        _0516_ = 8'b00001000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b10101110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b01111010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b01100101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b11101010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b11110100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b01010110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b01101100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b10101001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b01001110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b11010101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b10001101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b01101101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b00110111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b11001000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b11100111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b01111001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b11100100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b10010101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b10010001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b01100010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b10101100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b11010011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b11000010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b01011100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b00100100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b00000110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b01001001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b00001010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b00111010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b00110010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b11100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b11011011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b00001011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b01011110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b11011110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b00010100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b10111000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b11101110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b01000110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b10001000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b10010000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b00101010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b00100010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b11011100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b01001111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b10000001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b01100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b01110011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b00011001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b01011101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b01100100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b00111101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b01111110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b10100111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b11000100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b00010111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b01000100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b10010111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b01011111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b11101100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b00010011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b00001100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b11001101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b11010010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b11110011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b11111111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b00010000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b00100001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b11011010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b10110110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b10111100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b11110101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b00111000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b10011101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b10010010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b10001111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b01000000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b10100011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b01010001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b10101000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b10011111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b00111100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b01010000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b01111111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b00000010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b11111001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b01000101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b10000101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b00110011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b01001101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b01000011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b11111011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b10101010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b11101111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b11010000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b11001111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b01011000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b01001100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b01001010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b00111001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b10111110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b11001011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b01101010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b01011011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b10110001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b11111100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b00100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b11101101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b00000000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b11010001 ;
      256'b????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b01010011 ;
      256'b???????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b10000100 ;
      256'b??????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b00101111 ;
      256'b?????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b11100011 ;
      256'b????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b00101001 ;
      256'b???????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b10110011 ;
      256'b??????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b11010110 ;
      256'b?????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b00111011 ;
      256'b????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b01010010 ;
      256'b???????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b10100000 ;
      256'b??????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b01011010 ;
      256'b?????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b01101110 ;
      256'b????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b00011011 ;
      256'b???????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b00011010 ;
      256'b??????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b00101100 ;
      256'b?????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b10000011 ;
      256'b????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b00001001 ;
      256'b???????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b01110101 ;
      256'b??????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b10110010 ;
      256'b?????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b00100111 ;
      256'b????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b11101011 ;
      256'b???????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b11100010 ;
      256'b??????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b10000000 ;
      256'b?????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b00010010 ;
      256'b????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b00000111 ;
      256'b???????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b10011010 ;
      256'b??????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b00000101 ;
      256'b?????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b10010110 ;
      256'b????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b00011000 ;
      256'b???????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b11000011 ;
      256'b??????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b00100011 ;
      256'b?????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b11000111 ;
      256'b????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b00000100 ;
      256'b???????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b00010101 ;
      256'b??????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b00110001 ;
      256'b?????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b11011000 ;
      256'b????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b01110001 ;
      256'b???????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b11110001 ;
      256'b??????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b11100101 ;
      256'b?????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b10100101 ;
      256'b????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b00110100 ;
      256'b???????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b11001100 ;
      256'b??????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b11110111 ;
      256'b?????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b00111111 ;
      256'b????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b00110110 ;
      256'b???????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b00100110 ;
      256'b??????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b10010011 ;
      256'b?????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b11111101 ;
      256'b????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b10110111 ;
      256'b???????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b11000000 ;
      256'b??????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b01110010 ;
      256'b?????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b10100100 ;
      256'b????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b10011100 ;
      256'b???????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b10101111 ;
      256'b??????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b10100010 ;
      256'b?????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b11010100 ;
      256'b????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b10101101 ;
      256'b???????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b11110000 ;
      256'b??????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b01000111 ;
      256'b?????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b01011001 ;
      256'b????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b11111010 ;
      256'b???????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b01111101 ;
      256'b??????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b11001001 ;
      256'b?????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b10000010 ;
      256'b????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b11001010 ;
      256'b???????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b01110110 ;
      256'b??????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b10101011 ;
      256'b?????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b11010111 ;
      256'b????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b11111110 ;
      256'b???????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b00101011 ;
      256'b??????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b01100111 ;
      256'b?????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b00000001 ;
      256'b????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b00110000 ;
      256'b???????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b11000101 ;
      256'b??????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b01101111 ;
      256'b?????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b01101011 ;
      256'b????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b11110010 ;
      256'b???1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b01111011 ;
      256'b??1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b01110111 ;
      256'b?1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b01111100 ;
      256'b1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b01100011 ;
      default:
        _0516_ = \t0.t2.s0.out ;
    endcase
  end
  assign _0517_ = state_in[111:104] == 8'b11111111;
  assign _0518_ = state_in[111:104] == 8'b11111110;
  assign _0519_ = state_in[111:104] == 8'b11111101;
  assign _0520_ = state_in[111:104] == 8'b11111100;
  assign _0521_ = state_in[111:104] == 8'b11111011;
  assign _0522_ = state_in[111:104] == 8'b11111010;
  assign _0523_ = state_in[111:104] == 8'b11111001;
  assign _0524_ = state_in[111:104] == 8'b11111000;
  assign _0525_ = state_in[111:104] == 8'b11110111;
  assign _0526_ = state_in[111:104] == 8'b11110110;
  assign _0527_ = state_in[111:104] == 8'b11110101;
  assign _0528_ = state_in[111:104] == 8'b11110100;
  assign _0529_ = state_in[111:104] == 8'b11110011;
  assign _0530_ = state_in[111:104] == 8'b11110010;
  assign _0531_ = state_in[111:104] == 8'b11110001;
  assign _0532_ = state_in[111:104] == 8'b11110000;
  assign _0533_ = state_in[111:104] == 8'b11101111;
  assign _0534_ = state_in[111:104] == 8'b11101110;
  assign _0535_ = state_in[111:104] == 8'b11101101;
  assign _0536_ = state_in[111:104] == 8'b11101100;
  assign _0537_ = state_in[111:104] == 8'b11101011;
  assign _0538_ = state_in[111:104] == 8'b11101010;
  assign _0539_ = state_in[111:104] == 8'b11101001;
  assign _0540_ = state_in[111:104] == 8'b11101000;
  assign _0541_ = state_in[111:104] == 8'b11100111;
  assign _0542_ = state_in[111:104] == 8'b11100110;
  assign _0543_ = state_in[111:104] == 8'b11100101;
  assign _0544_ = state_in[111:104] == 8'b11100100;
  assign _0545_ = state_in[111:104] == 8'b11100011;
  assign _0546_ = state_in[111:104] == 8'b11100010;
  assign _0547_ = state_in[111:104] == 8'b11100001;
  assign _0548_ = state_in[111:104] == 8'b11100000;
  assign _0549_ = state_in[111:104] == 8'b11011111;
  assign _0550_ = state_in[111:104] == 8'b11011110;
  assign _0551_ = state_in[111:104] == 8'b11011101;
  assign _0552_ = state_in[111:104] == 8'b11011100;
  assign _0553_ = state_in[111:104] == 8'b11011011;
  assign _0554_ = state_in[111:104] == 8'b11011010;
  assign _0555_ = state_in[111:104] == 8'b11011001;
  assign _0556_ = state_in[111:104] == 8'b11011000;
  assign _0557_ = state_in[111:104] == 8'b11010111;
  assign _0558_ = state_in[111:104] == 8'b11010110;
  assign _0559_ = state_in[111:104] == 8'b11010101;
  assign _0560_ = state_in[111:104] == 8'b11010100;
  assign _0561_ = state_in[111:104] == 8'b11010011;
  assign _0562_ = state_in[111:104] == 8'b11010010;
  assign _0563_ = state_in[111:104] == 8'b11010001;
  assign _0564_ = state_in[111:104] == 8'b11010000;
  assign _0565_ = state_in[111:104] == 8'b11001111;
  assign _0566_ = state_in[111:104] == 8'b11001110;
  assign _0567_ = state_in[111:104] == 8'b11001101;
  assign _0568_ = state_in[111:104] == 8'b11001100;
  assign _0569_ = state_in[111:104] == 8'b11001011;
  assign _0570_ = state_in[111:104] == 8'b11001010;
  assign _0571_ = state_in[111:104] == 8'b11001001;
  assign _0572_ = state_in[111:104] == 8'b11001000;
  assign _0573_ = state_in[111:104] == 8'b11000111;
  assign _0574_ = state_in[111:104] == 8'b11000110;
  assign _0575_ = state_in[111:104] == 8'b11000101;
  assign _0576_ = state_in[111:104] == 8'b11000100;
  assign _0577_ = state_in[111:104] == 8'b11000011;
  assign _0578_ = state_in[111:104] == 8'b11000010;
  assign _0579_ = state_in[111:104] == 8'b11000001;
  assign _0580_ = state_in[111:104] == 8'b11000000;
  assign _0581_ = state_in[111:104] == 8'b10111111;
  assign _0582_ = state_in[111:104] == 8'b10111110;
  assign _0583_ = state_in[111:104] == 8'b10111101;
  assign _0584_ = state_in[111:104] == 8'b10111100;
  assign _0585_ = state_in[111:104] == 8'b10111011;
  assign _0586_ = state_in[111:104] == 8'b10111010;
  assign _0587_ = state_in[111:104] == 8'b10111001;
  assign _0588_ = state_in[111:104] == 8'b10111000;
  assign _0589_ = state_in[111:104] == 8'b10110111;
  assign _0590_ = state_in[111:104] == 8'b10110110;
  assign _0591_ = state_in[111:104] == 8'b10110101;
  assign _0592_ = state_in[111:104] == 8'b10110100;
  assign _0593_ = state_in[111:104] == 8'b10110011;
  assign _0594_ = state_in[111:104] == 8'b10110010;
  assign _0595_ = state_in[111:104] == 8'b10110001;
  assign _0596_ = state_in[111:104] == 8'b10110000;
  assign _0597_ = state_in[111:104] == 8'b10101111;
  assign _0598_ = state_in[111:104] == 8'b10101110;
  assign _0599_ = state_in[111:104] == 8'b10101101;
  assign _0600_ = state_in[111:104] == 8'b10101100;
  assign _0601_ = state_in[111:104] == 8'b10101011;
  assign _0602_ = state_in[111:104] == 8'b10101010;
  assign _0603_ = state_in[111:104] == 8'b10101001;
  assign _0604_ = state_in[111:104] == 8'b10101000;
  assign _0605_ = state_in[111:104] == 8'b10100111;
  assign _0606_ = state_in[111:104] == 8'b10100110;
  assign _0607_ = state_in[111:104] == 8'b10100101;
  assign _0608_ = state_in[111:104] == 8'b10100100;
  assign _0609_ = state_in[111:104] == 8'b10100011;
  assign _0610_ = state_in[111:104] == 8'b10100010;
  assign _0611_ = state_in[111:104] == 8'b10100001;
  assign _0612_ = state_in[111:104] == 8'b10100000;
  assign _0613_ = state_in[111:104] == 8'b10011111;
  assign _0614_ = state_in[111:104] == 8'b10011110;
  assign _0615_ = state_in[111:104] == 8'b10011101;
  assign _0616_ = state_in[111:104] == 8'b10011100;
  assign _0617_ = state_in[111:104] == 8'b10011011;
  assign _0618_ = state_in[111:104] == 8'b10011010;
  assign _0619_ = state_in[111:104] == 8'b10011001;
  assign _0620_ = state_in[111:104] == 8'b10011000;
  assign _0621_ = state_in[111:104] == 8'b10010111;
  assign _0622_ = state_in[111:104] == 8'b10010110;
  assign _0623_ = state_in[111:104] == 8'b10010101;
  assign _0624_ = state_in[111:104] == 8'b10010100;
  assign _0625_ = state_in[111:104] == 8'b10010011;
  assign _0626_ = state_in[111:104] == 8'b10010010;
  assign _0627_ = state_in[111:104] == 8'b10010001;
  assign _0628_ = state_in[111:104] == 8'b10010000;
  assign _0629_ = state_in[111:104] == 8'b10001111;
  assign _0630_ = state_in[111:104] == 8'b10001110;
  assign _0631_ = state_in[111:104] == 8'b10001101;
  assign _0632_ = state_in[111:104] == 8'b10001100;
  assign _0633_ = state_in[111:104] == 8'b10001011;
  assign _0634_ = state_in[111:104] == 8'b10001010;
  assign _0635_ = state_in[111:104] == 8'b10001001;
  assign _0636_ = state_in[111:104] == 8'b10001000;
  assign _0637_ = state_in[111:104] == 8'b10000111;
  assign _0638_ = state_in[111:104] == 8'b10000110;
  assign _0639_ = state_in[111:104] == 8'b10000101;
  assign _0640_ = state_in[111:104] == 8'b10000100;
  assign _0641_ = state_in[111:104] == 8'b10000011;
  assign _0642_ = state_in[111:104] == 8'b10000010;
  assign _0643_ = state_in[111:104] == 8'b10000001;
  assign _0644_ = state_in[111:104] == 8'b10000000;
  assign _0645_ = state_in[111:104] == 7'b1111111;
  assign _0646_ = state_in[111:104] == 7'b1111110;
  assign _0647_ = state_in[111:104] == 7'b1111101;
  assign _0648_ = state_in[111:104] == 7'b1111100;
  assign _0649_ = state_in[111:104] == 7'b1111011;
  assign _0650_ = state_in[111:104] == 7'b1111010;
  assign _0651_ = state_in[111:104] == 7'b1111001;
  assign _0652_ = state_in[111:104] == 7'b1111000;
  assign _0653_ = state_in[111:104] == 7'b1110111;
  assign _0654_ = state_in[111:104] == 7'b1110110;
  assign _0655_ = state_in[111:104] == 7'b1110101;
  assign _0656_ = state_in[111:104] == 7'b1110100;
  assign _0657_ = state_in[111:104] == 7'b1110011;
  assign _0658_ = state_in[111:104] == 7'b1110010;
  assign _0659_ = state_in[111:104] == 7'b1110001;
  assign _0660_ = state_in[111:104] == 7'b1110000;
  assign _0661_ = state_in[111:104] == 7'b1101111;
  assign _0662_ = state_in[111:104] == 7'b1101110;
  assign _0663_ = state_in[111:104] == 7'b1101101;
  assign _0664_ = state_in[111:104] == 7'b1101100;
  assign _0665_ = state_in[111:104] == 7'b1101011;
  assign _0666_ = state_in[111:104] == 7'b1101010;
  assign _0667_ = state_in[111:104] == 7'b1101001;
  assign _0668_ = state_in[111:104] == 7'b1101000;
  assign _0669_ = state_in[111:104] == 7'b1100111;
  assign _0670_ = state_in[111:104] == 7'b1100110;
  assign _0671_ = state_in[111:104] == 7'b1100101;
  assign _0672_ = state_in[111:104] == 7'b1100100;
  assign _0673_ = state_in[111:104] == 7'b1100011;
  assign _0674_ = state_in[111:104] == 7'b1100010;
  assign _0675_ = state_in[111:104] == 7'b1100001;
  assign _0676_ = state_in[111:104] == 7'b1100000;
  assign _0677_ = state_in[111:104] == 7'b1011111;
  assign _0678_ = state_in[111:104] == 7'b1011110;
  assign _0679_ = state_in[111:104] == 7'b1011101;
  assign _0680_ = state_in[111:104] == 7'b1011100;
  assign _0681_ = state_in[111:104] == 7'b1011011;
  assign _0682_ = state_in[111:104] == 7'b1011010;
  assign _0683_ = state_in[111:104] == 7'b1011001;
  assign _0684_ = state_in[111:104] == 7'b1011000;
  assign _0685_ = state_in[111:104] == 7'b1010111;
  assign _0686_ = state_in[111:104] == 7'b1010110;
  assign _0687_ = state_in[111:104] == 7'b1010101;
  assign _0688_ = state_in[111:104] == 7'b1010100;
  assign _0689_ = state_in[111:104] == 7'b1010011;
  assign _0690_ = state_in[111:104] == 7'b1010010;
  assign _0691_ = state_in[111:104] == 7'b1010001;
  assign _0692_ = state_in[111:104] == 7'b1010000;
  assign _0693_ = state_in[111:104] == 7'b1001111;
  assign _0694_ = state_in[111:104] == 7'b1001110;
  assign _0695_ = state_in[111:104] == 7'b1001101;
  assign _0696_ = state_in[111:104] == 7'b1001100;
  assign _0697_ = state_in[111:104] == 7'b1001011;
  assign _0698_ = state_in[111:104] == 7'b1001010;
  assign _0699_ = state_in[111:104] == 7'b1001001;
  assign _0700_ = state_in[111:104] == 7'b1001000;
  assign _0701_ = state_in[111:104] == 7'b1000111;
  assign _0702_ = state_in[111:104] == 7'b1000110;
  assign _0703_ = state_in[111:104] == 7'b1000101;
  assign _0704_ = state_in[111:104] == 7'b1000100;
  assign _0705_ = state_in[111:104] == 7'b1000011;
  assign _0706_ = state_in[111:104] == 7'b1000010;
  assign _0707_ = state_in[111:104] == 7'b1000001;
  assign _0708_ = state_in[111:104] == 7'b1000000;
  assign _0709_ = state_in[111:104] == 6'b111111;
  assign _0710_ = state_in[111:104] == 6'b111110;
  assign _0711_ = state_in[111:104] == 6'b111101;
  assign _0712_ = state_in[111:104] == 6'b111100;
  assign _0713_ = state_in[111:104] == 6'b111011;
  assign _0714_ = state_in[111:104] == 6'b111010;
  assign _0715_ = state_in[111:104] == 6'b111001;
  assign _0716_ = state_in[111:104] == 6'b111000;
  assign _0717_ = state_in[111:104] == 6'b110111;
  assign _0718_ = state_in[111:104] == 6'b110110;
  assign _0719_ = state_in[111:104] == 6'b110101;
  assign _0720_ = state_in[111:104] == 6'b110100;
  assign _0721_ = state_in[111:104] == 6'b110011;
  assign _0722_ = state_in[111:104] == 6'b110010;
  assign _0723_ = state_in[111:104] == 6'b110001;
  assign _0724_ = state_in[111:104] == 6'b110000;
  assign _0725_ = state_in[111:104] == 6'b101111;
  assign _0726_ = state_in[111:104] == 6'b101110;
  assign _0727_ = state_in[111:104] == 6'b101101;
  assign _0728_ = state_in[111:104] == 6'b101100;
  assign _0729_ = state_in[111:104] == 6'b101011;
  assign _0730_ = state_in[111:104] == 6'b101010;
  assign _0731_ = state_in[111:104] == 6'b101001;
  assign _0732_ = state_in[111:104] == 6'b101000;
  assign _0733_ = state_in[111:104] == 6'b100111;
  assign _0734_ = state_in[111:104] == 6'b100110;
  assign _0735_ = state_in[111:104] == 6'b100101;
  assign _0736_ = state_in[111:104] == 6'b100100;
  assign _0737_ = state_in[111:104] == 6'b100011;
  assign _0738_ = state_in[111:104] == 6'b100010;
  assign _0739_ = state_in[111:104] == 6'b100001;
  assign _0740_ = state_in[111:104] == 6'b100000;
  assign _0741_ = state_in[111:104] == 5'b11111;
  assign _0742_ = state_in[111:104] == 5'b11110;
  assign _0743_ = state_in[111:104] == 5'b11101;
  assign _0744_ = state_in[111:104] == 5'b11100;
  assign _0745_ = state_in[111:104] == 5'b11011;
  assign _0746_ = state_in[111:104] == 5'b11010;
  assign _0747_ = state_in[111:104] == 5'b11001;
  assign _0748_ = state_in[111:104] == 5'b11000;
  assign _0749_ = state_in[111:104] == 5'b10111;
  assign _0750_ = state_in[111:104] == 5'b10110;
  assign _0751_ = state_in[111:104] == 5'b10101;
  assign _0752_ = state_in[111:104] == 5'b10100;
  assign _0753_ = state_in[111:104] == 5'b10011;
  assign _0754_ = state_in[111:104] == 5'b10010;
  assign _0755_ = state_in[111:104] == 5'b10001;
  assign _0756_ = state_in[111:104] == 5'b10000;
  assign _0757_ = state_in[111:104] == 4'b1111;
  assign _0758_ = state_in[111:104] == 4'b1110;
  assign _0759_ = state_in[111:104] == 4'b1101;
  assign _0760_ = state_in[111:104] == 4'b1100;
  assign _0761_ = state_in[111:104] == 4'b1011;
  assign _0762_ = state_in[111:104] == 4'b1010;
  assign _0763_ = state_in[111:104] == 4'b1001;
  assign _0764_ = state_in[111:104] == 4'b1000;
  assign _0765_ = state_in[111:104] == 3'b111;
  assign _0766_ = state_in[111:104] == 3'b110;
  assign _0767_ = state_in[111:104] == 3'b101;
  assign _0768_ = state_in[111:104] == 3'b100;
  assign _0769_ = state_in[111:104] == 2'b11;
  assign _0770_ = state_in[111:104] == 2'b10;
  assign _0771_ = state_in[111:104] == 1'b1;
  assign _0772_ = ! state_in[111:104];
  always @(posedge clk)
      \t0.t2.s4.out <= _0773_;
  wire [255:0] fangyuan6;
  assign fangyuan6 = { _0772_, _0771_, _0770_, _0769_, _0768_, _0767_, _0766_, _0765_, _0764_, _0763_, _0762_, _0761_, _0760_, _0759_, _0758_, _0757_, _0756_, _0755_, _0754_, _0753_, _0752_, _0751_, _0750_, _0749_, _0748_, _0747_, _0746_, _0745_, _0744_, _0743_, _0742_, _0741_, _0740_, _0739_, _0738_, _0737_, _0736_, _0735_, _0734_, _0733_, _0732_, _0731_, _0730_, _0729_, _0728_, _0727_, _0726_, _0725_, _0724_, _0723_, _0722_, _0721_, _0720_, _0719_, _0718_, _0717_, _0716_, _0715_, _0714_, _0713_, _0712_, _0711_, _0710_, _0709_, _0708_, _0707_, _0706_, _0705_, _0704_, _0703_, _0702_, _0701_, _0700_, _0699_, _0698_, _0697_, _0696_, _0695_, _0694_, _0693_, _0692_, _0691_, _0690_, _0689_, _0688_, _0687_, _0686_, _0685_, _0684_, _0683_, _0682_, _0681_, _0680_, _0679_, _0678_, _0677_, _0676_, _0675_, _0674_, _0673_, _0672_, _0671_, _0670_, _0669_, _0668_, _0667_, _0666_, _0665_, _0664_, _0663_, _0662_, _0661_, _0660_, _0659_, _0658_, _0657_, _0656_, _0655_, _0654_, _0653_, _0652_, _0651_, _0650_, _0649_, _0648_, _0647_, _0646_, _0645_, _0644_, _0643_, _0642_, _0641_, _0640_, _0639_, _0638_, _0637_, _0636_, _0635_, _0634_, _0633_, _0632_, _0631_, _0630_, _0629_, _0628_, _0627_, _0626_, _0625_, _0624_, _0623_, _0622_, _0621_, _0620_, _0619_, _0618_, _0617_, _0616_, _0615_, _0614_, _0613_, _0612_, _0611_, _0610_, _0609_, _0608_, _0607_, _0606_, _0605_, _0604_, _0603_, _0602_, _0601_, _0600_, _0599_, _0598_, _0597_, _0596_, _0595_, _0594_, _0593_, _0592_, _0591_, _0590_, _0589_, _0588_, _0587_, _0586_, _0585_, _0584_, _0583_, _0582_, _0581_, _0580_, _0579_, _0578_, _0577_, _0576_, _0575_, _0574_, _0573_, _0572_, _0571_, _0570_, _0569_, _0568_, _0567_, _0566_, _0565_, _0564_, _0563_, _0562_, _0561_, _0560_, _0559_, _0558_, _0557_, _0556_, _0555_, _0554_, _0553_, _0552_, _0551_, _0550_, _0549_, _0548_, _0547_, _0546_, _0545_, _0544_, _0543_, _0542_, _0541_, _0540_, _0539_, _0538_, _0537_, _0536_, _0535_, _0534_, _0533_, _0532_, _0531_, _0530_, _0529_, _0528_, _0527_, _0526_, _0525_, _0524_, _0523_, _0522_, _0521_, _0520_, _0519_, _0518_, _0517_ };

  always @(\t0.t2.s4.out or fangyuan6) begin
    casez (fangyuan6)
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1 :
        _0773_ = 8'b00101100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1? :
        _0773_ = 8'b01101101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?? :
        _0773_ = 8'b10101000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??? :
        _0773_ = 8'b01111011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???? :
        _0773_ = 8'b00011110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????? :
        _0773_ = 8'b01011010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????? :
        _0773_ = 8'b00101001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????? :
        _0773_ = 8'b10000010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????? :
        _0773_ = 8'b11010000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????? :
        _0773_ = 8'b10000100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????? :
        _0773_ = 8'b11010111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????? :
        _0773_ = 8'b01100101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????? :
        _0773_ = 8'b00011010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????? :
        _0773_ = 8'b00001001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????? :
        _0773_ = 8'b01011001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????? :
        _0773_ = 8'b00000011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????? :
        _0773_ = 8'b10100101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????? :
        _0773_ = 8'b01010000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????? :
        _0773_ = 8'b10101010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????? :
        _0773_ = 8'b10000111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????? :
        _0773_ = 8'b11001001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????? :
        _0773_ = 8'b00010101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????? :
        _0773_ = 8'b00111100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????? :
        _0773_ = 8'b00101101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????? :
        _0773_ = 8'b00110011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????? :
        _0773_ = 8'b00000111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????? :
        _0773_ = 8'b10101001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????? :
        _0773_ = 8'b11010010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????? :
        _0773_ = 8'b00100010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????? :
        _0773_ = 8'b00101011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????? :
        _0773_ = 8'b11101011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????? :
        _0773_ = 8'b11011001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????? :
        _0773_ = 8'b00100111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????? :
        _0773_ = 8'b00111010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????? :
        _0773_ = 8'b10011001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????? :
        _0773_ = 8'b00010111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????? :
        _0773_ = 8'b01101001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????? :
        _0773_ = 8'b10101110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????? :
        _0773_ = 8'b01101010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????? :
        _0773_ = 8'b11000010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????? :
        _0773_ = 8'b00011100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????? :
        _0773_ = 8'b11110111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????? :
        _0773_ = 8'b00000110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????? :
        _0773_ = 8'b10010000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????? :
        _0773_ = 8'b11001100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????? :
        _0773_ = 8'b01110001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????? :
        _0773_ = 8'b01111100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????? :
        _0773_ = 8'b11100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????? :
        _0773_ = 8'b00001111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????? :
        _0773_ = 8'b00001101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????? :
        _0773_ = 8'b01100001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????? :
        _0773_ = 8'b10010110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????? :
        _0773_ = 8'b00111110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????? :
        _0773_ = 8'b11101000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????? :
        _0773_ = 8'b10100001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????? :
        _0773_ = 8'b11001011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????? :
        _0773_ = 8'b10010111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????? :
        _0773_ = 8'b01110011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????? :
        _0773_ = 8'b01010111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????? :
        _0773_ = 8'b00111000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????? :
        _0773_ = 8'b01011100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????? :
        _0773_ = 8'b01001010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????? :
        _0773_ = 8'b11110000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????? :
        _0773_ = 8'b01101111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????? :
        _0773_ = 8'b00010000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b01000111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b11110100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b11001010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b11001111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b11110011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b10101100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b11011000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b01001001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b10011100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b10110001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b00000001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b11011010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b01101110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b10001011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b11010101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b11110010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b11010011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b00110001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b00111001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b11000100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b01000011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b10111101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b10011111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b10111000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b01001000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b00001100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b10010010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b00010100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b01110100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b01100100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b11011011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b10101101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b00010110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b10111100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b10100111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b00101000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b01101011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b11000111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b10001100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b00001011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b00111011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b01010100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b01000100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b10100011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b10011110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b00011001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b11000000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b11100110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b00110010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b10111010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b11001000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b01111010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b11111100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b01010101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b10010011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b00101110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b10001000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b00110101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b10111110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b11000011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b00100110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b00011000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b10000001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b10111111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b11111101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b11100101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b00100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b01000010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b10101111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b01110111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b01100011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b11110001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b01110000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b00100001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b00111111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b00000101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b10000000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b01011101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b10100010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b01001011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b00100101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b01111000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b10100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b11111110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b00000100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b11101001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b10001010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b00010001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b01100110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b10011010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b10000110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b11101101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b01001111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b11000101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b10111011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b10000101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b10110000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b10011000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b10010100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b01110010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b01100111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b10001101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b11010100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b10110110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b01111001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b11100011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b01000000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b11000001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b00000000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b10111001 ;
      256'b????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b10100110 ;
      256'b???????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b00010011 ;
      256'b??????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b01011110 ;
      256'b?????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b11011101 ;
      256'b????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b01010010 ;
      256'b???????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b01111101 ;
      256'b??????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b10110111 ;
      256'b?????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b01110110 ;
      256'b????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b10100100 ;
      256'b???????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b01011011 ;
      256'b??????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b10110100 ;
      256'b?????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b11011100 ;
      256'b????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b00110110 ;
      256'b???????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b00110100 ;
      256'b??????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b01011000 ;
      256'b?????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b00011101 ;
      256'b????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b00010010 ;
      256'b???????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b11101010 ;
      256'b??????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b01111111 ;
      256'b?????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b01001110 ;
      256'b????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b11001101 ;
      256'b???????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b11011111 ;
      256'b??????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b00011011 ;
      256'b?????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b00100100 ;
      256'b????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b00001110 ;
      256'b???????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b00101111 ;
      256'b??????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b00001010 ;
      256'b?????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b00110111 ;
      256'b????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b00110000 ;
      256'b???????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b10011101 ;
      256'b??????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b01000110 ;
      256'b?????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b10010101 ;
      256'b????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b00001000 ;
      256'b???????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b00101010 ;
      256'b??????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b01100010 ;
      256'b?????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b10101011 ;
      256'b????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b11100010 ;
      256'b???????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b11111001 ;
      256'b??????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b11010001 ;
      256'b?????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b01010001 ;
      256'b????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b01101000 ;
      256'b???????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b10000011 ;
      256'b??????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b11110101 ;
      256'b?????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b01111110 ;
      256'b????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b01101100 ;
      256'b???????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b01001100 ;
      256'b??????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b00111101 ;
      256'b?????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b11100001 ;
      256'b????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b01110101 ;
      256'b???????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b10011011 ;
      256'b??????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b11100100 ;
      256'b?????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b01010011 ;
      256'b????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b00100011 ;
      256'b???????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b01000101 ;
      256'b??????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b01011111 ;
      256'b?????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b10110011 ;
      256'b????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b01000001 ;
      256'b???????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b11111011 ;
      256'b??????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b10001110 ;
      256'b?????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b10110010 ;
      256'b????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b11101111 ;
      256'b???????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b11111010 ;
      256'b??????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b10001001 ;
      256'b?????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b00011111 ;
      256'b????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b10001111 ;
      256'b???????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b11101100 ;
      256'b??????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b01001101 ;
      256'b?????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b10110101 ;
      256'b????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b11100111 ;
      256'b???????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b01010110 ;
      256'b??????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b11001110 ;
      256'b?????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b00000010 ;
      256'b????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b01100000 ;
      256'b???????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b10010001 ;
      256'b??????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b11011110 ;
      256'b?????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b11010110 ;
      256'b????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b11111111 ;
      256'b???1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b11110110 ;
      256'b??1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b11101110 ;
      256'b?1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b11111000 ;
      256'b1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b11000110 ;
      default:
        _0773_ = \t0.t2.s4.out ;
    endcase
  end
  assign p03[15:8] = \t0.t3.s0.out ^ \t0.t3.s4.out ;
  always @(posedge clk)
      \t0.t3.s0.out <= _0774_;
  wire [255:0] fangyuan7;
  assign fangyuan7 = { _1030_, _1029_, _1028_, _1027_, _1026_, _1025_, _1024_, _1023_, _1022_, _1021_, _1020_, _1019_, _1018_, _1017_, _1016_, _1015_, _1014_, _1013_, _1012_, _1011_, _1010_, _1009_, _1008_, _1007_, _1006_, _1005_, _1004_, _1003_, _1002_, _1001_, _1000_, _0999_, _0998_, _0997_, _0996_, _0995_, _0994_, _0993_, _0992_, _0991_, _0990_, _0989_, _0988_, _0987_, _0986_, _0985_, _0984_, _0983_, _0982_, _0981_, _0980_, _0979_, _0978_, _0977_, _0976_, _0975_, _0974_, _0973_, _0972_, _0971_, _0970_, _0969_, _0968_, _0967_, _0966_, _0965_, _0964_, _0963_, _0962_, _0961_, _0960_, _0959_, _0958_, _0957_, _0956_, _0955_, _0954_, _0953_, _0952_, _0951_, _0950_, _0949_, _0948_, _0947_, _0946_, _0945_, _0944_, _0943_, _0942_, _0941_, _0940_, _0939_, _0938_, _0937_, _0936_, _0935_, _0934_, _0933_, _0932_, _0931_, _0930_, _0929_, _0928_, _0927_, _0926_, _0925_, _0924_, _0923_, _0922_, _0921_, _0920_, _0919_, _0918_, _0917_, _0916_, _0915_, _0914_, _0913_, _0912_, _0911_, _0910_, _0909_, _0908_, _0907_, _0906_, _0905_, _0904_, _0903_, _0902_, _0901_, _0900_, _0899_, _0898_, _0897_, _0896_, _0895_, _0894_, _0893_, _0892_, _0891_, _0890_, _0889_, _0888_, _0887_, _0886_, _0885_, _0884_, _0883_, _0882_, _0881_, _0880_, _0879_, _0878_, _0877_, _0876_, _0875_, _0874_, _0873_, _0872_, _0871_, _0870_, _0869_, _0868_, _0867_, _0866_, _0865_, _0864_, _0863_, _0862_, _0861_, _0860_, _0859_, _0858_, _0857_, _0856_, _0855_, _0854_, _0853_, _0852_, _0851_, _0850_, _0849_, _0848_, _0847_, _0846_, _0845_, _0844_, _0843_, _0842_, _0841_, _0840_, _0839_, _0838_, _0837_, _0836_, _0835_, _0834_, _0833_, _0832_, _0831_, _0830_, _0829_, _0828_, _0827_, _0826_, _0825_, _0824_, _0823_, _0822_, _0821_, _0820_, _0819_, _0818_, _0817_, _0816_, _0815_, _0814_, _0813_, _0812_, _0811_, _0810_, _0809_, _0808_, _0807_, _0806_, _0805_, _0804_, _0803_, _0802_, _0801_, _0800_, _0799_, _0798_, _0797_, _0796_, _0795_, _0794_, _0793_, _0792_, _0791_, _0790_, _0789_, _0788_, _0787_, _0786_, _0785_, _0784_, _0783_, _0782_, _0781_, _0780_, _0779_, _0778_, _0777_, _0776_, _0775_ };

  always @(\t0.t3.s0.out or fangyuan7) begin
    casez (fangyuan7)
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1 :
        _0774_ = 8'b00010110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1? :
        _0774_ = 8'b10111011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?? :
        _0774_ = 8'b01010100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??? :
        _0774_ = 8'b10110000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???? :
        _0774_ = 8'b00001111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????? :
        _0774_ = 8'b00101101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????? :
        _0774_ = 8'b10011001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????? :
        _0774_ = 8'b01000001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????? :
        _0774_ = 8'b01101000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????? :
        _0774_ = 8'b01000010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????? :
        _0774_ = 8'b11100110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????? :
        _0774_ = 8'b10111111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????? :
        _0774_ = 8'b00001101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????? :
        _0774_ = 8'b10001001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????? :
        _0774_ = 8'b10100001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????? :
        _0774_ = 8'b10001100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????? :
        _0774_ = 8'b11011111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????? :
        _0774_ = 8'b00101000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????? :
        _0774_ = 8'b01010101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????? :
        _0774_ = 8'b11001110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????? :
        _0774_ = 8'b11101001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????? :
        _0774_ = 8'b10000111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????? :
        _0774_ = 8'b00011110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????? :
        _0774_ = 8'b10011011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????? :
        _0774_ = 8'b10010100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????? :
        _0774_ = 8'b10001110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????? :
        _0774_ = 8'b11011001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????? :
        _0774_ = 8'b01101001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????? :
        _0774_ = 8'b00010001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????? :
        _0774_ = 8'b10011000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????? :
        _0774_ = 8'b11111000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????? :
        _0774_ = 8'b11100001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????? :
        _0774_ = 8'b10011110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????? :
        _0774_ = 8'b00011101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????? :
        _0774_ = 8'b11000001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????? :
        _0774_ = 8'b10000110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????? :
        _0774_ = 8'b10111001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????? :
        _0774_ = 8'b01010111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????? :
        _0774_ = 8'b00110101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????? :
        _0774_ = 8'b01100001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????? :
        _0774_ = 8'b00001110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????? :
        _0774_ = 8'b11110110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????? :
        _0774_ = 8'b00000011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????? :
        _0774_ = 8'b01001000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????? :
        _0774_ = 8'b01100110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????? :
        _0774_ = 8'b10110101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????? :
        _0774_ = 8'b00111110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????? :
        _0774_ = 8'b01110000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????? :
        _0774_ = 8'b10001010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????? :
        _0774_ = 8'b10001011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????? :
        _0774_ = 8'b10111101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????? :
        _0774_ = 8'b01001011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????? :
        _0774_ = 8'b00011111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????? :
        _0774_ = 8'b01110100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????? :
        _0774_ = 8'b11011101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????? :
        _0774_ = 8'b11101000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????? :
        _0774_ = 8'b11000110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????? :
        _0774_ = 8'b10110100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????? :
        _0774_ = 8'b10100110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????? :
        _0774_ = 8'b00011100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????? :
        _0774_ = 8'b00101110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????? :
        _0774_ = 8'b00100101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????? :
        _0774_ = 8'b01111000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????? :
        _0774_ = 8'b10111010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????? :
        _0774_ = 8'b00001000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b10101110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b01111010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b01100101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b11101010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b11110100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b01010110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b01101100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b10101001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b01001110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b11010101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b10001101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b01101101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b00110111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b11001000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b11100111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b01111001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b11100100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b10010101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b10010001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b01100010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b10101100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b11010011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b11000010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b01011100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b00100100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b00000110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b01001001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b00001010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b00111010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b00110010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b11100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b11011011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b00001011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b01011110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b11011110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b00010100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b10111000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b11101110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b01000110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b10001000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b10010000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b00101010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b00100010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b11011100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b01001111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b10000001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b01100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b01110011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b00011001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b01011101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b01100100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b00111101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b01111110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b10100111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b11000100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b00010111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b01000100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b10010111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b01011111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b11101100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b00010011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b00001100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b11001101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b11010010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b11110011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b11111111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b00010000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b00100001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b11011010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b10110110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b10111100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b11110101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b00111000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b10011101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b10010010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b10001111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b01000000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b10100011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b01010001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b10101000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b10011111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b00111100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b01010000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b01111111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b00000010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b11111001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b01000101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b10000101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b00110011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b01001101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b01000011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b11111011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b10101010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b11101111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b11010000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b11001111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b01011000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b01001100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b01001010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b00111001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b10111110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b11001011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b01101010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b01011011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b10110001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b11111100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b00100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b11101101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b00000000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b11010001 ;
      256'b????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b01010011 ;
      256'b???????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b10000100 ;
      256'b??????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b00101111 ;
      256'b?????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b11100011 ;
      256'b????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b00101001 ;
      256'b???????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b10110011 ;
      256'b??????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b11010110 ;
      256'b?????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b00111011 ;
      256'b????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b01010010 ;
      256'b???????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b10100000 ;
      256'b??????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b01011010 ;
      256'b?????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b01101110 ;
      256'b????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b00011011 ;
      256'b???????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b00011010 ;
      256'b??????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b00101100 ;
      256'b?????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b10000011 ;
      256'b????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b00001001 ;
      256'b???????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b01110101 ;
      256'b??????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b10110010 ;
      256'b?????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b00100111 ;
      256'b????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b11101011 ;
      256'b???????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b11100010 ;
      256'b??????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b10000000 ;
      256'b?????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b00010010 ;
      256'b????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b00000111 ;
      256'b???????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b10011010 ;
      256'b??????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b00000101 ;
      256'b?????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b10010110 ;
      256'b????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b00011000 ;
      256'b???????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b11000011 ;
      256'b??????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b00100011 ;
      256'b?????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b11000111 ;
      256'b????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b00000100 ;
      256'b???????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b00010101 ;
      256'b??????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b00110001 ;
      256'b?????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b11011000 ;
      256'b????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b01110001 ;
      256'b???????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b11110001 ;
      256'b??????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b11100101 ;
      256'b?????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b10100101 ;
      256'b????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b00110100 ;
      256'b???????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b11001100 ;
      256'b??????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b11110111 ;
      256'b?????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b00111111 ;
      256'b????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b00110110 ;
      256'b???????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b00100110 ;
      256'b??????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b10010011 ;
      256'b?????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b11111101 ;
      256'b????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b10110111 ;
      256'b???????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b11000000 ;
      256'b??????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b01110010 ;
      256'b?????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b10100100 ;
      256'b????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b10011100 ;
      256'b???????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b10101111 ;
      256'b??????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b10100010 ;
      256'b?????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b11010100 ;
      256'b????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b10101101 ;
      256'b???????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b11110000 ;
      256'b??????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b01000111 ;
      256'b?????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b01011001 ;
      256'b????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b11111010 ;
      256'b???????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b01111101 ;
      256'b??????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b11001001 ;
      256'b?????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b10000010 ;
      256'b????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b11001010 ;
      256'b???????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b01110110 ;
      256'b??????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b10101011 ;
      256'b?????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b11010111 ;
      256'b????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b11111110 ;
      256'b???????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b00101011 ;
      256'b??????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b01100111 ;
      256'b?????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b00000001 ;
      256'b????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b00110000 ;
      256'b???????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b11000101 ;
      256'b??????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b01101111 ;
      256'b?????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b01101011 ;
      256'b????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b11110010 ;
      256'b???1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b01111011 ;
      256'b??1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b01110111 ;
      256'b?1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b01111100 ;
      256'b1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b01100011 ;
      default:
        _0774_ = \t0.t3.s0.out ;
    endcase
  end
  assign _0775_ = state_in[103:96] == 8'b11111111;
  assign _0776_ = state_in[103:96] == 8'b11111110;
  assign _0777_ = state_in[103:96] == 8'b11111101;
  assign _0778_ = state_in[103:96] == 8'b11111100;
  assign _0779_ = state_in[103:96] == 8'b11111011;
  assign _0780_ = state_in[103:96] == 8'b11111010;
  assign _0781_ = state_in[103:96] == 8'b11111001;
  assign _0782_ = state_in[103:96] == 8'b11111000;
  assign _0783_ = state_in[103:96] == 8'b11110111;
  assign _0784_ = state_in[103:96] == 8'b11110110;
  assign _0785_ = state_in[103:96] == 8'b11110101;
  assign _0786_ = state_in[103:96] == 8'b11110100;
  assign _0787_ = state_in[103:96] == 8'b11110011;
  assign _0788_ = state_in[103:96] == 8'b11110010;
  assign _0789_ = state_in[103:96] == 8'b11110001;
  assign _0790_ = state_in[103:96] == 8'b11110000;
  assign _0791_ = state_in[103:96] == 8'b11101111;
  assign _0792_ = state_in[103:96] == 8'b11101110;
  assign _0793_ = state_in[103:96] == 8'b11101101;
  assign _0794_ = state_in[103:96] == 8'b11101100;
  assign _0795_ = state_in[103:96] == 8'b11101011;
  assign _0796_ = state_in[103:96] == 8'b11101010;
  assign _0797_ = state_in[103:96] == 8'b11101001;
  assign _0798_ = state_in[103:96] == 8'b11101000;
  assign _0799_ = state_in[103:96] == 8'b11100111;
  assign _0800_ = state_in[103:96] == 8'b11100110;
  assign _0801_ = state_in[103:96] == 8'b11100101;
  assign _0802_ = state_in[103:96] == 8'b11100100;
  assign _0803_ = state_in[103:96] == 8'b11100011;
  assign _0804_ = state_in[103:96] == 8'b11100010;
  assign _0805_ = state_in[103:96] == 8'b11100001;
  assign _0806_ = state_in[103:96] == 8'b11100000;
  assign _0807_ = state_in[103:96] == 8'b11011111;
  assign _0808_ = state_in[103:96] == 8'b11011110;
  assign _0809_ = state_in[103:96] == 8'b11011101;
  assign _0810_ = state_in[103:96] == 8'b11011100;
  assign _0811_ = state_in[103:96] == 8'b11011011;
  assign _0812_ = state_in[103:96] == 8'b11011010;
  assign _0813_ = state_in[103:96] == 8'b11011001;
  assign _0814_ = state_in[103:96] == 8'b11011000;
  assign _0815_ = state_in[103:96] == 8'b11010111;
  assign _0816_ = state_in[103:96] == 8'b11010110;
  assign _0817_ = state_in[103:96] == 8'b11010101;
  assign _0818_ = state_in[103:96] == 8'b11010100;
  assign _0819_ = state_in[103:96] == 8'b11010011;
  assign _0820_ = state_in[103:96] == 8'b11010010;
  assign _0821_ = state_in[103:96] == 8'b11010001;
  assign _0822_ = state_in[103:96] == 8'b11010000;
  assign _0823_ = state_in[103:96] == 8'b11001111;
  assign _0824_ = state_in[103:96] == 8'b11001110;
  assign _0825_ = state_in[103:96] == 8'b11001101;
  assign _0826_ = state_in[103:96] == 8'b11001100;
  assign _0827_ = state_in[103:96] == 8'b11001011;
  assign _0828_ = state_in[103:96] == 8'b11001010;
  assign _0829_ = state_in[103:96] == 8'b11001001;
  assign _0830_ = state_in[103:96] == 8'b11001000;
  assign _0831_ = state_in[103:96] == 8'b11000111;
  assign _0832_ = state_in[103:96] == 8'b11000110;
  assign _0833_ = state_in[103:96] == 8'b11000101;
  assign _0834_ = state_in[103:96] == 8'b11000100;
  assign _0835_ = state_in[103:96] == 8'b11000011;
  assign _0836_ = state_in[103:96] == 8'b11000010;
  assign _0837_ = state_in[103:96] == 8'b11000001;
  assign _0838_ = state_in[103:96] == 8'b11000000;
  assign _0839_ = state_in[103:96] == 8'b10111111;
  assign _0840_ = state_in[103:96] == 8'b10111110;
  assign _0841_ = state_in[103:96] == 8'b10111101;
  assign _0842_ = state_in[103:96] == 8'b10111100;
  assign _0843_ = state_in[103:96] == 8'b10111011;
  assign _0844_ = state_in[103:96] == 8'b10111010;
  assign _0845_ = state_in[103:96] == 8'b10111001;
  assign _0846_ = state_in[103:96] == 8'b10111000;
  assign _0847_ = state_in[103:96] == 8'b10110111;
  assign _0848_ = state_in[103:96] == 8'b10110110;
  assign _0849_ = state_in[103:96] == 8'b10110101;
  assign _0850_ = state_in[103:96] == 8'b10110100;
  assign _0851_ = state_in[103:96] == 8'b10110011;
  assign _0852_ = state_in[103:96] == 8'b10110010;
  assign _0853_ = state_in[103:96] == 8'b10110001;
  assign _0854_ = state_in[103:96] == 8'b10110000;
  assign _0855_ = state_in[103:96] == 8'b10101111;
  assign _0856_ = state_in[103:96] == 8'b10101110;
  assign _0857_ = state_in[103:96] == 8'b10101101;
  assign _0858_ = state_in[103:96] == 8'b10101100;
  assign _0859_ = state_in[103:96] == 8'b10101011;
  assign _0860_ = state_in[103:96] == 8'b10101010;
  assign _0861_ = state_in[103:96] == 8'b10101001;
  assign _0862_ = state_in[103:96] == 8'b10101000;
  assign _0863_ = state_in[103:96] == 8'b10100111;
  assign _0864_ = state_in[103:96] == 8'b10100110;
  assign _0865_ = state_in[103:96] == 8'b10100101;
  assign _0866_ = state_in[103:96] == 8'b10100100;
  assign _0867_ = state_in[103:96] == 8'b10100011;
  assign _0868_ = state_in[103:96] == 8'b10100010;
  assign _0869_ = state_in[103:96] == 8'b10100001;
  assign _0870_ = state_in[103:96] == 8'b10100000;
  assign _0871_ = state_in[103:96] == 8'b10011111;
  assign _0872_ = state_in[103:96] == 8'b10011110;
  assign _0873_ = state_in[103:96] == 8'b10011101;
  assign _0874_ = state_in[103:96] == 8'b10011100;
  assign _0875_ = state_in[103:96] == 8'b10011011;
  assign _0876_ = state_in[103:96] == 8'b10011010;
  assign _0877_ = state_in[103:96] == 8'b10011001;
  assign _0878_ = state_in[103:96] == 8'b10011000;
  assign _0879_ = state_in[103:96] == 8'b10010111;
  assign _0880_ = state_in[103:96] == 8'b10010110;
  assign _0881_ = state_in[103:96] == 8'b10010101;
  assign _0882_ = state_in[103:96] == 8'b10010100;
  assign _0883_ = state_in[103:96] == 8'b10010011;
  assign _0884_ = state_in[103:96] == 8'b10010010;
  assign _0885_ = state_in[103:96] == 8'b10010001;
  assign _0886_ = state_in[103:96] == 8'b10010000;
  assign _0887_ = state_in[103:96] == 8'b10001111;
  assign _0888_ = state_in[103:96] == 8'b10001110;
  assign _0889_ = state_in[103:96] == 8'b10001101;
  assign _0890_ = state_in[103:96] == 8'b10001100;
  assign _0891_ = state_in[103:96] == 8'b10001011;
  assign _0892_ = state_in[103:96] == 8'b10001010;
  assign _0893_ = state_in[103:96] == 8'b10001001;
  assign _0894_ = state_in[103:96] == 8'b10001000;
  assign _0895_ = state_in[103:96] == 8'b10000111;
  assign _0896_ = state_in[103:96] == 8'b10000110;
  assign _0897_ = state_in[103:96] == 8'b10000101;
  assign _0898_ = state_in[103:96] == 8'b10000100;
  assign _0899_ = state_in[103:96] == 8'b10000011;
  assign _0900_ = state_in[103:96] == 8'b10000010;
  assign _0901_ = state_in[103:96] == 8'b10000001;
  assign _0902_ = state_in[103:96] == 8'b10000000;
  assign _0903_ = state_in[103:96] == 7'b1111111;
  assign _0904_ = state_in[103:96] == 7'b1111110;
  assign _0905_ = state_in[103:96] == 7'b1111101;
  assign _0906_ = state_in[103:96] == 7'b1111100;
  assign _0907_ = state_in[103:96] == 7'b1111011;
  assign _0908_ = state_in[103:96] == 7'b1111010;
  assign _0909_ = state_in[103:96] == 7'b1111001;
  assign _0910_ = state_in[103:96] == 7'b1111000;
  assign _0911_ = state_in[103:96] == 7'b1110111;
  assign _0912_ = state_in[103:96] == 7'b1110110;
  assign _0913_ = state_in[103:96] == 7'b1110101;
  assign _0914_ = state_in[103:96] == 7'b1110100;
  assign _0915_ = state_in[103:96] == 7'b1110011;
  assign _0916_ = state_in[103:96] == 7'b1110010;
  assign _0917_ = state_in[103:96] == 7'b1110001;
  assign _0918_ = state_in[103:96] == 7'b1110000;
  assign _0919_ = state_in[103:96] == 7'b1101111;
  assign _0920_ = state_in[103:96] == 7'b1101110;
  assign _0921_ = state_in[103:96] == 7'b1101101;
  assign _0922_ = state_in[103:96] == 7'b1101100;
  assign _0923_ = state_in[103:96] == 7'b1101011;
  assign _0924_ = state_in[103:96] == 7'b1101010;
  assign _0925_ = state_in[103:96] == 7'b1101001;
  assign _0926_ = state_in[103:96] == 7'b1101000;
  assign _0927_ = state_in[103:96] == 7'b1100111;
  assign _0928_ = state_in[103:96] == 7'b1100110;
  assign _0929_ = state_in[103:96] == 7'b1100101;
  assign _0930_ = state_in[103:96] == 7'b1100100;
  assign _0931_ = state_in[103:96] == 7'b1100011;
  assign _0932_ = state_in[103:96] == 7'b1100010;
  assign _0933_ = state_in[103:96] == 7'b1100001;
  assign _0934_ = state_in[103:96] == 7'b1100000;
  assign _0935_ = state_in[103:96] == 7'b1011111;
  assign _0936_ = state_in[103:96] == 7'b1011110;
  assign _0937_ = state_in[103:96] == 7'b1011101;
  assign _0938_ = state_in[103:96] == 7'b1011100;
  assign _0939_ = state_in[103:96] == 7'b1011011;
  assign _0940_ = state_in[103:96] == 7'b1011010;
  assign _0941_ = state_in[103:96] == 7'b1011001;
  assign _0942_ = state_in[103:96] == 7'b1011000;
  assign _0943_ = state_in[103:96] == 7'b1010111;
  assign _0944_ = state_in[103:96] == 7'b1010110;
  assign _0945_ = state_in[103:96] == 7'b1010101;
  assign _0946_ = state_in[103:96] == 7'b1010100;
  assign _0947_ = state_in[103:96] == 7'b1010011;
  assign _0948_ = state_in[103:96] == 7'b1010010;
  assign _0949_ = state_in[103:96] == 7'b1010001;
  assign _0950_ = state_in[103:96] == 7'b1010000;
  assign _0951_ = state_in[103:96] == 7'b1001111;
  assign _0952_ = state_in[103:96] == 7'b1001110;
  assign _0953_ = state_in[103:96] == 7'b1001101;
  assign _0954_ = state_in[103:96] == 7'b1001100;
  assign _0955_ = state_in[103:96] == 7'b1001011;
  assign _0956_ = state_in[103:96] == 7'b1001010;
  assign _0957_ = state_in[103:96] == 7'b1001001;
  assign _0958_ = state_in[103:96] == 7'b1001000;
  assign _0959_ = state_in[103:96] == 7'b1000111;
  assign _0960_ = state_in[103:96] == 7'b1000110;
  assign _0961_ = state_in[103:96] == 7'b1000101;
  assign _0962_ = state_in[103:96] == 7'b1000100;
  assign _0963_ = state_in[103:96] == 7'b1000011;
  assign _0964_ = state_in[103:96] == 7'b1000010;
  assign _0965_ = state_in[103:96] == 7'b1000001;
  assign _0966_ = state_in[103:96] == 7'b1000000;
  assign _0967_ = state_in[103:96] == 6'b111111;
  assign _0968_ = state_in[103:96] == 6'b111110;
  assign _0969_ = state_in[103:96] == 6'b111101;
  assign _0970_ = state_in[103:96] == 6'b111100;
  assign _0971_ = state_in[103:96] == 6'b111011;
  assign _0972_ = state_in[103:96] == 6'b111010;
  assign _0973_ = state_in[103:96] == 6'b111001;
  assign _0974_ = state_in[103:96] == 6'b111000;
  assign _0975_ = state_in[103:96] == 6'b110111;
  assign _0976_ = state_in[103:96] == 6'b110110;
  assign _0977_ = state_in[103:96] == 6'b110101;
  assign _0978_ = state_in[103:96] == 6'b110100;
  assign _0979_ = state_in[103:96] == 6'b110011;
  assign _0980_ = state_in[103:96] == 6'b110010;
  assign _0981_ = state_in[103:96] == 6'b110001;
  assign _0982_ = state_in[103:96] == 6'b110000;
  assign _0983_ = state_in[103:96] == 6'b101111;
  assign _0984_ = state_in[103:96] == 6'b101110;
  assign _0985_ = state_in[103:96] == 6'b101101;
  assign _0986_ = state_in[103:96] == 6'b101100;
  assign _0987_ = state_in[103:96] == 6'b101011;
  assign _0988_ = state_in[103:96] == 6'b101010;
  assign _0989_ = state_in[103:96] == 6'b101001;
  assign _0990_ = state_in[103:96] == 6'b101000;
  assign _0991_ = state_in[103:96] == 6'b100111;
  assign _0992_ = state_in[103:96] == 6'b100110;
  assign _0993_ = state_in[103:96] == 6'b100101;
  assign _0994_ = state_in[103:96] == 6'b100100;
  assign _0995_ = state_in[103:96] == 6'b100011;
  assign _0996_ = state_in[103:96] == 6'b100010;
  assign _0997_ = state_in[103:96] == 6'b100001;
  assign _0998_ = state_in[103:96] == 6'b100000;
  assign _0999_ = state_in[103:96] == 5'b11111;
  assign _1000_ = state_in[103:96] == 5'b11110;
  assign _1001_ = state_in[103:96] == 5'b11101;
  assign _1002_ = state_in[103:96] == 5'b11100;
  assign _1003_ = state_in[103:96] == 5'b11011;
  assign _1004_ = state_in[103:96] == 5'b11010;
  assign _1005_ = state_in[103:96] == 5'b11001;
  assign _1006_ = state_in[103:96] == 5'b11000;
  assign _1007_ = state_in[103:96] == 5'b10111;
  assign _1008_ = state_in[103:96] == 5'b10110;
  assign _1009_ = state_in[103:96] == 5'b10101;
  assign _1010_ = state_in[103:96] == 5'b10100;
  assign _1011_ = state_in[103:96] == 5'b10011;
  assign _1012_ = state_in[103:96] == 5'b10010;
  assign _1013_ = state_in[103:96] == 5'b10001;
  assign _1014_ = state_in[103:96] == 5'b10000;
  assign _1015_ = state_in[103:96] == 4'b1111;
  assign _1016_ = state_in[103:96] == 4'b1110;
  assign _1017_ = state_in[103:96] == 4'b1101;
  assign _1018_ = state_in[103:96] == 4'b1100;
  assign _1019_ = state_in[103:96] == 4'b1011;
  assign _1020_ = state_in[103:96] == 4'b1010;
  assign _1021_ = state_in[103:96] == 4'b1001;
  assign _1022_ = state_in[103:96] == 4'b1000;
  assign _1023_ = state_in[103:96] == 3'b111;
  assign _1024_ = state_in[103:96] == 3'b110;
  assign _1025_ = state_in[103:96] == 3'b101;
  assign _1026_ = state_in[103:96] == 3'b100;
  assign _1027_ = state_in[103:96] == 2'b11;
  assign _1028_ = state_in[103:96] == 2'b10;
  assign _1029_ = state_in[103:96] == 1'b1;
  assign _1030_ = ! state_in[103:96];
  always @(posedge clk)
      \t0.t3.s4.out <= _1031_;
  wire [255:0] fangyuan8;
  assign fangyuan8 = { _1030_, _1029_, _1028_, _1027_, _1026_, _1025_, _1024_, _1023_, _1022_, _1021_, _1020_, _1019_, _1018_, _1017_, _1016_, _1015_, _1014_, _1013_, _1012_, _1011_, _1010_, _1009_, _1008_, _1007_, _1006_, _1005_, _1004_, _1003_, _1002_, _1001_, _1000_, _0999_, _0998_, _0997_, _0996_, _0995_, _0994_, _0993_, _0992_, _0991_, _0990_, _0989_, _0988_, _0987_, _0986_, _0985_, _0984_, _0983_, _0982_, _0981_, _0980_, _0979_, _0978_, _0977_, _0976_, _0975_, _0974_, _0973_, _0972_, _0971_, _0970_, _0969_, _0968_, _0967_, _0966_, _0965_, _0964_, _0963_, _0962_, _0961_, _0960_, _0959_, _0958_, _0957_, _0956_, _0955_, _0954_, _0953_, _0952_, _0951_, _0950_, _0949_, _0948_, _0947_, _0946_, _0945_, _0944_, _0943_, _0942_, _0941_, _0940_, _0939_, _0938_, _0937_, _0936_, _0935_, _0934_, _0933_, _0932_, _0931_, _0930_, _0929_, _0928_, _0927_, _0926_, _0925_, _0924_, _0923_, _0922_, _0921_, _0920_, _0919_, _0918_, _0917_, _0916_, _0915_, _0914_, _0913_, _0912_, _0911_, _0910_, _0909_, _0908_, _0907_, _0906_, _0905_, _0904_, _0903_, _0902_, _0901_, _0900_, _0899_, _0898_, _0897_, _0896_, _0895_, _0894_, _0893_, _0892_, _0891_, _0890_, _0889_, _0888_, _0887_, _0886_, _0885_, _0884_, _0883_, _0882_, _0881_, _0880_, _0879_, _0878_, _0877_, _0876_, _0875_, _0874_, _0873_, _0872_, _0871_, _0870_, _0869_, _0868_, _0867_, _0866_, _0865_, _0864_, _0863_, _0862_, _0861_, _0860_, _0859_, _0858_, _0857_, _0856_, _0855_, _0854_, _0853_, _0852_, _0851_, _0850_, _0849_, _0848_, _0847_, _0846_, _0845_, _0844_, _0843_, _0842_, _0841_, _0840_, _0839_, _0838_, _0837_, _0836_, _0835_, _0834_, _0833_, _0832_, _0831_, _0830_, _0829_, _0828_, _0827_, _0826_, _0825_, _0824_, _0823_, _0822_, _0821_, _0820_, _0819_, _0818_, _0817_, _0816_, _0815_, _0814_, _0813_, _0812_, _0811_, _0810_, _0809_, _0808_, _0807_, _0806_, _0805_, _0804_, _0803_, _0802_, _0801_, _0800_, _0799_, _0798_, _0797_, _0796_, _0795_, _0794_, _0793_, _0792_, _0791_, _0790_, _0789_, _0788_, _0787_, _0786_, _0785_, _0784_, _0783_, _0782_, _0781_, _0780_, _0779_, _0778_, _0777_, _0776_, _0775_ };

  always @(\t0.t3.s4.out or fangyuan8) begin
    casez (fangyuan8)
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1 :
        _1031_ = 8'b00101100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1? :
        _1031_ = 8'b01101101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?? :
        _1031_ = 8'b10101000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??? :
        _1031_ = 8'b01111011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???? :
        _1031_ = 8'b00011110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????? :
        _1031_ = 8'b01011010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????? :
        _1031_ = 8'b00101001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????? :
        _1031_ = 8'b10000010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????? :
        _1031_ = 8'b11010000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????? :
        _1031_ = 8'b10000100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????? :
        _1031_ = 8'b11010111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????? :
        _1031_ = 8'b01100101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????? :
        _1031_ = 8'b00011010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????? :
        _1031_ = 8'b00001001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????? :
        _1031_ = 8'b01011001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????? :
        _1031_ = 8'b00000011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????? :
        _1031_ = 8'b10100101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????? :
        _1031_ = 8'b01010000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????? :
        _1031_ = 8'b10101010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????? :
        _1031_ = 8'b10000111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????? :
        _1031_ = 8'b11001001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????? :
        _1031_ = 8'b00010101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????? :
        _1031_ = 8'b00111100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????? :
        _1031_ = 8'b00101101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????? :
        _1031_ = 8'b00110011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????? :
        _1031_ = 8'b00000111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????? :
        _1031_ = 8'b10101001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????? :
        _1031_ = 8'b11010010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????? :
        _1031_ = 8'b00100010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????? :
        _1031_ = 8'b00101011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????? :
        _1031_ = 8'b11101011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????? :
        _1031_ = 8'b11011001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????? :
        _1031_ = 8'b00100111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????? :
        _1031_ = 8'b00111010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????? :
        _1031_ = 8'b10011001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????? :
        _1031_ = 8'b00010111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????? :
        _1031_ = 8'b01101001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????? :
        _1031_ = 8'b10101110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????? :
        _1031_ = 8'b01101010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????? :
        _1031_ = 8'b11000010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????? :
        _1031_ = 8'b00011100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????? :
        _1031_ = 8'b11110111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????? :
        _1031_ = 8'b00000110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????? :
        _1031_ = 8'b10010000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????? :
        _1031_ = 8'b11001100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????? :
        _1031_ = 8'b01110001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????? :
        _1031_ = 8'b01111100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????? :
        _1031_ = 8'b11100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????? :
        _1031_ = 8'b00001111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????? :
        _1031_ = 8'b00001101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????? :
        _1031_ = 8'b01100001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????? :
        _1031_ = 8'b10010110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????? :
        _1031_ = 8'b00111110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????? :
        _1031_ = 8'b11101000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????? :
        _1031_ = 8'b10100001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????? :
        _1031_ = 8'b11001011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????? :
        _1031_ = 8'b10010111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????? :
        _1031_ = 8'b01110011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????? :
        _1031_ = 8'b01010111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????? :
        _1031_ = 8'b00111000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????? :
        _1031_ = 8'b01011100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????? :
        _1031_ = 8'b01001010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????? :
        _1031_ = 8'b11110000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????? :
        _1031_ = 8'b01101111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????? :
        _1031_ = 8'b00010000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b01000111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b11110100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b11001010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b11001111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b11110011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b10101100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b11011000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b01001001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b10011100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b10110001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b00000001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b11011010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b01101110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b10001011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b11010101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b11110010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b11010011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b00110001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b00111001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b11000100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b01000011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b10111101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b10011111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b10111000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b01001000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b00001100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b10010010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b00010100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b01110100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b01100100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b11011011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b10101101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b00010110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b10111100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b10100111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b00101000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b01101011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b11000111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b10001100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b00001011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b00111011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b01010100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b01000100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b10100011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b10011110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b00011001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b11000000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b11100110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b00110010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b10111010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b11001000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b01111010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b11111100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b01010101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b10010011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b00101110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b10001000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b00110101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b10111110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b11000011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b00100110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b00011000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b10000001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b10111111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b11111101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b11100101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b00100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b01000010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b10101111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b01110111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b01100011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b11110001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b01110000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b00100001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b00111111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b00000101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b10000000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b01011101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b10100010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b01001011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b00100101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b01111000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b10100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b11111110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b00000100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b11101001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b10001010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b00010001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b01100110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b10011010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b10000110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b11101101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b01001111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b11000101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b10111011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b10000101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b10110000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b10011000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b10010100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b01110010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b01100111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b10001101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b11010100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b10110110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b01111001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b11100011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b01000000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b11000001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b00000000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b10111001 ;
      256'b????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b10100110 ;
      256'b???????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b00010011 ;
      256'b??????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b01011110 ;
      256'b?????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b11011101 ;
      256'b????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b01010010 ;
      256'b???????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b01111101 ;
      256'b??????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b10110111 ;
      256'b?????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b01110110 ;
      256'b????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b10100100 ;
      256'b???????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b01011011 ;
      256'b??????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b10110100 ;
      256'b?????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b11011100 ;
      256'b????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b00110110 ;
      256'b???????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b00110100 ;
      256'b??????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b01011000 ;
      256'b?????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b00011101 ;
      256'b????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b00010010 ;
      256'b???????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b11101010 ;
      256'b??????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b01111111 ;
      256'b?????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b01001110 ;
      256'b????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b11001101 ;
      256'b???????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b11011111 ;
      256'b??????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b00011011 ;
      256'b?????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b00100100 ;
      256'b????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b00001110 ;
      256'b???????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b00101111 ;
      256'b??????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b00001010 ;
      256'b?????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b00110111 ;
      256'b????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b00110000 ;
      256'b???????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b10011101 ;
      256'b??????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b01000110 ;
      256'b?????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b10010101 ;
      256'b????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b00001000 ;
      256'b???????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b00101010 ;
      256'b??????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b01100010 ;
      256'b?????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b10101011 ;
      256'b????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b11100010 ;
      256'b???????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b11111001 ;
      256'b??????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b11010001 ;
      256'b?????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b01010001 ;
      256'b????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b01101000 ;
      256'b???????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b10000011 ;
      256'b??????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b11110101 ;
      256'b?????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b01111110 ;
      256'b????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b01101100 ;
      256'b???????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b01001100 ;
      256'b??????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b00111101 ;
      256'b?????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b11100001 ;
      256'b????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b01110101 ;
      256'b???????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b10011011 ;
      256'b??????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b11100100 ;
      256'b?????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b01010011 ;
      256'b????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b00100011 ;
      256'b???????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b01000101 ;
      256'b??????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b01011111 ;
      256'b?????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b10110011 ;
      256'b????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b01000001 ;
      256'b???????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b11111011 ;
      256'b??????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b10001110 ;
      256'b?????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b10110010 ;
      256'b????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b11101111 ;
      256'b???????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b11111010 ;
      256'b??????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b10001001 ;
      256'b?????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b00011111 ;
      256'b????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b10001111 ;
      256'b???????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b11101100 ;
      256'b??????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b01001101 ;
      256'b?????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b10110101 ;
      256'b????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b11100111 ;
      256'b???????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b01010110 ;
      256'b??????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b11001110 ;
      256'b?????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b00000010 ;
      256'b????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b01100000 ;
      256'b???????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b10010001 ;
      256'b??????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b11011110 ;
      256'b?????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b11010110 ;
      256'b????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b11111111 ;
      256'b???1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b11110110 ;
      256'b??1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b11101110 ;
      256'b?1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b11111000 ;
      256'b1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b11000110 ;
      default:
        _1031_ = \t0.t3.s4.out ;
    endcase
  end
  assign p10[7:0] = \t1.t0.s0.out ^ \t1.t0.s4.out ;
  always @(posedge clk)
      \t1.t0.s0.out <= _1032_;
  wire [255:0] fangyuan9;
  assign fangyuan9 = { _1288_, _1287_, _1286_, _1285_, _1284_, _1283_, _1282_, _1281_, _1280_, _1279_, _1278_, _1277_, _1276_, _1275_, _1274_, _1273_, _1272_, _1271_, _1270_, _1269_, _1268_, _1267_, _1266_, _1265_, _1264_, _1263_, _1262_, _1261_, _1260_, _1259_, _1258_, _1257_, _1256_, _1255_, _1254_, _1253_, _1252_, _1251_, _1250_, _1249_, _1248_, _1247_, _1246_, _1245_, _1244_, _1243_, _1242_, _1241_, _1240_, _1239_, _1238_, _1237_, _1236_, _1235_, _1234_, _1233_, _1232_, _1231_, _1230_, _1229_, _1228_, _1227_, _1226_, _1225_, _1224_, _1223_, _1222_, _1221_, _1220_, _1219_, _1218_, _1217_, _1216_, _1215_, _1214_, _1213_, _1212_, _1211_, _1210_, _1209_, _1208_, _1207_, _1206_, _1205_, _1204_, _1203_, _1202_, _1201_, _1200_, _1199_, _1198_, _1197_, _1196_, _1195_, _1194_, _1193_, _1192_, _1191_, _1190_, _1189_, _1188_, _1187_, _1186_, _1185_, _1184_, _1183_, _1182_, _1181_, _1180_, _1179_, _1178_, _1177_, _1176_, _1175_, _1174_, _1173_, _1172_, _1171_, _1170_, _1169_, _1168_, _1167_, _1166_, _1165_, _1164_, _1163_, _1162_, _1161_, _1160_, _1159_, _1158_, _1157_, _1156_, _1155_, _1154_, _1153_, _1152_, _1151_, _1150_, _1149_, _1148_, _1147_, _1146_, _1145_, _1144_, _1143_, _1142_, _1141_, _1140_, _1139_, _1138_, _1137_, _1136_, _1135_, _1134_, _1133_, _1132_, _1131_, _1130_, _1129_, _1128_, _1127_, _1126_, _1125_, _1124_, _1123_, _1122_, _1121_, _1120_, _1119_, _1118_, _1117_, _1116_, _1115_, _1114_, _1113_, _1112_, _1111_, _1110_, _1109_, _1108_, _1107_, _1106_, _1105_, _1104_, _1103_, _1102_, _1101_, _1100_, _1099_, _1098_, _1097_, _1096_, _1095_, _1094_, _1093_, _1092_, _1091_, _1090_, _1089_, _1088_, _1087_, _1086_, _1085_, _1084_, _1083_, _1082_, _1081_, _1080_, _1079_, _1078_, _1077_, _1076_, _1075_, _1074_, _1073_, _1072_, _1071_, _1070_, _1069_, _1068_, _1067_, _1066_, _1065_, _1064_, _1063_, _1062_, _1061_, _1060_, _1059_, _1058_, _1057_, _1056_, _1055_, _1054_, _1053_, _1052_, _1051_, _1050_, _1049_, _1048_, _1047_, _1046_, _1045_, _1044_, _1043_, _1042_, _1041_, _1040_, _1039_, _1038_, _1037_, _1036_, _1035_, _1034_, _1033_ };

  always @(\t1.t0.s0.out or fangyuan9) begin
    casez (fangyuan9)
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1 :
        _1032_ = 8'b00010110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1? :
        _1032_ = 8'b10111011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?? :
        _1032_ = 8'b01010100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??? :
        _1032_ = 8'b10110000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???? :
        _1032_ = 8'b00001111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????? :
        _1032_ = 8'b00101101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????? :
        _1032_ = 8'b10011001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????? :
        _1032_ = 8'b01000001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????? :
        _1032_ = 8'b01101000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????? :
        _1032_ = 8'b01000010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????? :
        _1032_ = 8'b11100110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????? :
        _1032_ = 8'b10111111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????? :
        _1032_ = 8'b00001101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????? :
        _1032_ = 8'b10001001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????? :
        _1032_ = 8'b10100001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????? :
        _1032_ = 8'b10001100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????? :
        _1032_ = 8'b11011111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????? :
        _1032_ = 8'b00101000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????? :
        _1032_ = 8'b01010101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????? :
        _1032_ = 8'b11001110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????? :
        _1032_ = 8'b11101001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????? :
        _1032_ = 8'b10000111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????? :
        _1032_ = 8'b00011110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????? :
        _1032_ = 8'b10011011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????? :
        _1032_ = 8'b10010100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????? :
        _1032_ = 8'b10001110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????? :
        _1032_ = 8'b11011001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????? :
        _1032_ = 8'b01101001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????? :
        _1032_ = 8'b00010001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????? :
        _1032_ = 8'b10011000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????? :
        _1032_ = 8'b11111000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????? :
        _1032_ = 8'b11100001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????? :
        _1032_ = 8'b10011110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????? :
        _1032_ = 8'b00011101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????? :
        _1032_ = 8'b11000001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????? :
        _1032_ = 8'b10000110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????? :
        _1032_ = 8'b10111001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????? :
        _1032_ = 8'b01010111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????? :
        _1032_ = 8'b00110101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????? :
        _1032_ = 8'b01100001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????? :
        _1032_ = 8'b00001110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????? :
        _1032_ = 8'b11110110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????? :
        _1032_ = 8'b00000011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????? :
        _1032_ = 8'b01001000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????? :
        _1032_ = 8'b01100110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????? :
        _1032_ = 8'b10110101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????? :
        _1032_ = 8'b00111110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????? :
        _1032_ = 8'b01110000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????? :
        _1032_ = 8'b10001010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????? :
        _1032_ = 8'b10001011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????? :
        _1032_ = 8'b10111101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????? :
        _1032_ = 8'b01001011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????? :
        _1032_ = 8'b00011111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????? :
        _1032_ = 8'b01110100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????? :
        _1032_ = 8'b11011101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????? :
        _1032_ = 8'b11101000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????? :
        _1032_ = 8'b11000110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????? :
        _1032_ = 8'b10110100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????? :
        _1032_ = 8'b10100110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????? :
        _1032_ = 8'b00011100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????? :
        _1032_ = 8'b00101110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????? :
        _1032_ = 8'b00100101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????? :
        _1032_ = 8'b01111000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????? :
        _1032_ = 8'b10111010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????? :
        _1032_ = 8'b00001000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b10101110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b01111010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b01100101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b11101010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b11110100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b01010110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b01101100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b10101001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b01001110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b11010101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b10001101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b01101101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b00110111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b11001000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b11100111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b01111001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b11100100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b10010101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b10010001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b01100010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b10101100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b11010011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b11000010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b01011100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b00100100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b00000110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b01001001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b00001010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b00111010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b00110010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b11100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b11011011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b00001011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b01011110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b11011110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b00010100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b10111000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b11101110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b01000110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b10001000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b10010000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b00101010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b00100010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b11011100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b01001111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b10000001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b01100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b01110011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b00011001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b01011101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b01100100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b00111101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b01111110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b10100111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b11000100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b00010111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b01000100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b10010111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b01011111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b11101100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b00010011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b00001100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b11001101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b11010010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b11110011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b11111111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b00010000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b00100001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b11011010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b10110110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b10111100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b11110101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b00111000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b10011101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b10010010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b10001111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b01000000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b10100011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b01010001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b10101000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b10011111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b00111100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b01010000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b01111111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b00000010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b11111001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b01000101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b10000101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b00110011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b01001101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b01000011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b11111011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b10101010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b11101111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b11010000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b11001111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b01011000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b01001100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b01001010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b00111001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b10111110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b11001011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b01101010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b01011011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b10110001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b11111100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b00100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b11101101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b00000000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b11010001 ;
      256'b????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b01010011 ;
      256'b???????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b10000100 ;
      256'b??????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b00101111 ;
      256'b?????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b11100011 ;
      256'b????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b00101001 ;
      256'b???????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b10110011 ;
      256'b??????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b11010110 ;
      256'b?????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b00111011 ;
      256'b????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b01010010 ;
      256'b???????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b10100000 ;
      256'b??????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b01011010 ;
      256'b?????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b01101110 ;
      256'b????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b00011011 ;
      256'b???????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b00011010 ;
      256'b??????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b00101100 ;
      256'b?????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b10000011 ;
      256'b????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b00001001 ;
      256'b???????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b01110101 ;
      256'b??????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b10110010 ;
      256'b?????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b00100111 ;
      256'b????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b11101011 ;
      256'b???????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b11100010 ;
      256'b??????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b10000000 ;
      256'b?????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b00010010 ;
      256'b????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b00000111 ;
      256'b???????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b10011010 ;
      256'b??????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b00000101 ;
      256'b?????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b10010110 ;
      256'b????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b00011000 ;
      256'b???????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b11000011 ;
      256'b??????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b00100011 ;
      256'b?????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b11000111 ;
      256'b????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b00000100 ;
      256'b???????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b00010101 ;
      256'b??????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b00110001 ;
      256'b?????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b11011000 ;
      256'b????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b01110001 ;
      256'b???????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b11110001 ;
      256'b??????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b11100101 ;
      256'b?????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b10100101 ;
      256'b????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b00110100 ;
      256'b???????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b11001100 ;
      256'b??????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b11110111 ;
      256'b?????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b00111111 ;
      256'b????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b00110110 ;
      256'b???????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b00100110 ;
      256'b??????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b10010011 ;
      256'b?????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b11111101 ;
      256'b????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b10110111 ;
      256'b???????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b11000000 ;
      256'b??????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b01110010 ;
      256'b?????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b10100100 ;
      256'b????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b10011100 ;
      256'b???????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b10101111 ;
      256'b??????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b10100010 ;
      256'b?????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b11010100 ;
      256'b????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b10101101 ;
      256'b???????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b11110000 ;
      256'b??????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b01000111 ;
      256'b?????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b01011001 ;
      256'b????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b11111010 ;
      256'b???????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b01111101 ;
      256'b??????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b11001001 ;
      256'b?????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b10000010 ;
      256'b????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b11001010 ;
      256'b???????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b01110110 ;
      256'b??????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b10101011 ;
      256'b?????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b11010111 ;
      256'b????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b11111110 ;
      256'b???????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b00101011 ;
      256'b??????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b01100111 ;
      256'b?????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b00000001 ;
      256'b????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b00110000 ;
      256'b???????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b11000101 ;
      256'b??????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b01101111 ;
      256'b?????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b01101011 ;
      256'b????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b11110010 ;
      256'b???1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b01111011 ;
      256'b??1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b01110111 ;
      256'b?1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b01111100 ;
      256'b1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b01100011 ;
      default:
        _1032_ = \t1.t0.s0.out ;
    endcase
  end
  assign _1033_ = state_in[95:88] == 8'b11111111;
  assign _1034_ = state_in[95:88] == 8'b11111110;
  assign _1035_ = state_in[95:88] == 8'b11111101;
  assign _1036_ = state_in[95:88] == 8'b11111100;
  assign _1037_ = state_in[95:88] == 8'b11111011;
  assign _1038_ = state_in[95:88] == 8'b11111010;
  assign _1039_ = state_in[95:88] == 8'b11111001;
  assign _1040_ = state_in[95:88] == 8'b11111000;
  assign _1041_ = state_in[95:88] == 8'b11110111;
  assign _1042_ = state_in[95:88] == 8'b11110110;
  assign _1043_ = state_in[95:88] == 8'b11110101;
  assign _1044_ = state_in[95:88] == 8'b11110100;
  assign _1045_ = state_in[95:88] == 8'b11110011;
  assign _1046_ = state_in[95:88] == 8'b11110010;
  assign _1047_ = state_in[95:88] == 8'b11110001;
  assign _1048_ = state_in[95:88] == 8'b11110000;
  assign _1049_ = state_in[95:88] == 8'b11101111;
  assign _1050_ = state_in[95:88] == 8'b11101110;
  assign _1051_ = state_in[95:88] == 8'b11101101;
  assign _1052_ = state_in[95:88] == 8'b11101100;
  assign _1053_ = state_in[95:88] == 8'b11101011;
  assign _1054_ = state_in[95:88] == 8'b11101010;
  assign _1055_ = state_in[95:88] == 8'b11101001;
  assign _1056_ = state_in[95:88] == 8'b11101000;
  assign _1057_ = state_in[95:88] == 8'b11100111;
  assign _1058_ = state_in[95:88] == 8'b11100110;
  assign _1059_ = state_in[95:88] == 8'b11100101;
  assign _1060_ = state_in[95:88] == 8'b11100100;
  assign _1061_ = state_in[95:88] == 8'b11100011;
  assign _1062_ = state_in[95:88] == 8'b11100010;
  assign _1063_ = state_in[95:88] == 8'b11100001;
  assign _1064_ = state_in[95:88] == 8'b11100000;
  assign _1065_ = state_in[95:88] == 8'b11011111;
  assign _1066_ = state_in[95:88] == 8'b11011110;
  assign _1067_ = state_in[95:88] == 8'b11011101;
  assign _1068_ = state_in[95:88] == 8'b11011100;
  assign _1069_ = state_in[95:88] == 8'b11011011;
  assign _1070_ = state_in[95:88] == 8'b11011010;
  assign _1071_ = state_in[95:88] == 8'b11011001;
  assign _1072_ = state_in[95:88] == 8'b11011000;
  assign _1073_ = state_in[95:88] == 8'b11010111;
  assign _1074_ = state_in[95:88] == 8'b11010110;
  assign _1075_ = state_in[95:88] == 8'b11010101;
  assign _1076_ = state_in[95:88] == 8'b11010100;
  assign _1077_ = state_in[95:88] == 8'b11010011;
  assign _1078_ = state_in[95:88] == 8'b11010010;
  assign _1079_ = state_in[95:88] == 8'b11010001;
  assign _1080_ = state_in[95:88] == 8'b11010000;
  assign _1081_ = state_in[95:88] == 8'b11001111;
  assign _1082_ = state_in[95:88] == 8'b11001110;
  assign _1083_ = state_in[95:88] == 8'b11001101;
  assign _1084_ = state_in[95:88] == 8'b11001100;
  assign _1085_ = state_in[95:88] == 8'b11001011;
  assign _1086_ = state_in[95:88] == 8'b11001010;
  assign _1087_ = state_in[95:88] == 8'b11001001;
  assign _1088_ = state_in[95:88] == 8'b11001000;
  assign _1089_ = state_in[95:88] == 8'b11000111;
  assign _1090_ = state_in[95:88] == 8'b11000110;
  assign _1091_ = state_in[95:88] == 8'b11000101;
  assign _1092_ = state_in[95:88] == 8'b11000100;
  assign _1093_ = state_in[95:88] == 8'b11000011;
  assign _1094_ = state_in[95:88] == 8'b11000010;
  assign _1095_ = state_in[95:88] == 8'b11000001;
  assign _1096_ = state_in[95:88] == 8'b11000000;
  assign _1097_ = state_in[95:88] == 8'b10111111;
  assign _1098_ = state_in[95:88] == 8'b10111110;
  assign _1099_ = state_in[95:88] == 8'b10111101;
  assign _1100_ = state_in[95:88] == 8'b10111100;
  assign _1101_ = state_in[95:88] == 8'b10111011;
  assign _1102_ = state_in[95:88] == 8'b10111010;
  assign _1103_ = state_in[95:88] == 8'b10111001;
  assign _1104_ = state_in[95:88] == 8'b10111000;
  assign _1105_ = state_in[95:88] == 8'b10110111;
  assign _1106_ = state_in[95:88] == 8'b10110110;
  assign _1107_ = state_in[95:88] == 8'b10110101;
  assign _1108_ = state_in[95:88] == 8'b10110100;
  assign _1109_ = state_in[95:88] == 8'b10110011;
  assign _1110_ = state_in[95:88] == 8'b10110010;
  assign _1111_ = state_in[95:88] == 8'b10110001;
  assign _1112_ = state_in[95:88] == 8'b10110000;
  assign _1113_ = state_in[95:88] == 8'b10101111;
  assign _1114_ = state_in[95:88] == 8'b10101110;
  assign _1115_ = state_in[95:88] == 8'b10101101;
  assign _1116_ = state_in[95:88] == 8'b10101100;
  assign _1117_ = state_in[95:88] == 8'b10101011;
  assign _1118_ = state_in[95:88] == 8'b10101010;
  assign _1119_ = state_in[95:88] == 8'b10101001;
  assign _1120_ = state_in[95:88] == 8'b10101000;
  assign _1121_ = state_in[95:88] == 8'b10100111;
  assign _1122_ = state_in[95:88] == 8'b10100110;
  assign _1123_ = state_in[95:88] == 8'b10100101;
  assign _1124_ = state_in[95:88] == 8'b10100100;
  assign _1125_ = state_in[95:88] == 8'b10100011;
  assign _1126_ = state_in[95:88] == 8'b10100010;
  assign _1127_ = state_in[95:88] == 8'b10100001;
  assign _1128_ = state_in[95:88] == 8'b10100000;
  assign _1129_ = state_in[95:88] == 8'b10011111;
  assign _1130_ = state_in[95:88] == 8'b10011110;
  assign _1131_ = state_in[95:88] == 8'b10011101;
  assign _1132_ = state_in[95:88] == 8'b10011100;
  assign _1133_ = state_in[95:88] == 8'b10011011;
  assign _1134_ = state_in[95:88] == 8'b10011010;
  assign _1135_ = state_in[95:88] == 8'b10011001;
  assign _1136_ = state_in[95:88] == 8'b10011000;
  assign _1137_ = state_in[95:88] == 8'b10010111;
  assign _1138_ = state_in[95:88] == 8'b10010110;
  assign _1139_ = state_in[95:88] == 8'b10010101;
  assign _1140_ = state_in[95:88] == 8'b10010100;
  assign _1141_ = state_in[95:88] == 8'b10010011;
  assign _1142_ = state_in[95:88] == 8'b10010010;
  assign _1143_ = state_in[95:88] == 8'b10010001;
  assign _1144_ = state_in[95:88] == 8'b10010000;
  assign _1145_ = state_in[95:88] == 8'b10001111;
  assign _1146_ = state_in[95:88] == 8'b10001110;
  assign _1147_ = state_in[95:88] == 8'b10001101;
  assign _1148_ = state_in[95:88] == 8'b10001100;
  assign _1149_ = state_in[95:88] == 8'b10001011;
  assign _1150_ = state_in[95:88] == 8'b10001010;
  assign _1151_ = state_in[95:88] == 8'b10001001;
  assign _1152_ = state_in[95:88] == 8'b10001000;
  assign _1153_ = state_in[95:88] == 8'b10000111;
  assign _1154_ = state_in[95:88] == 8'b10000110;
  assign _1155_ = state_in[95:88] == 8'b10000101;
  assign _1156_ = state_in[95:88] == 8'b10000100;
  assign _1157_ = state_in[95:88] == 8'b10000011;
  assign _1158_ = state_in[95:88] == 8'b10000010;
  assign _1159_ = state_in[95:88] == 8'b10000001;
  assign _1160_ = state_in[95:88] == 8'b10000000;
  assign _1161_ = state_in[95:88] == 7'b1111111;
  assign _1162_ = state_in[95:88] == 7'b1111110;
  assign _1163_ = state_in[95:88] == 7'b1111101;
  assign _1164_ = state_in[95:88] == 7'b1111100;
  assign _1165_ = state_in[95:88] == 7'b1111011;
  assign _1166_ = state_in[95:88] == 7'b1111010;
  assign _1167_ = state_in[95:88] == 7'b1111001;
  assign _1168_ = state_in[95:88] == 7'b1111000;
  assign _1169_ = state_in[95:88] == 7'b1110111;
  assign _1170_ = state_in[95:88] == 7'b1110110;
  assign _1171_ = state_in[95:88] == 7'b1110101;
  assign _1172_ = state_in[95:88] == 7'b1110100;
  assign _1173_ = state_in[95:88] == 7'b1110011;
  assign _1174_ = state_in[95:88] == 7'b1110010;
  assign _1175_ = state_in[95:88] == 7'b1110001;
  assign _1176_ = state_in[95:88] == 7'b1110000;
  assign _1177_ = state_in[95:88] == 7'b1101111;
  assign _1178_ = state_in[95:88] == 7'b1101110;
  assign _1179_ = state_in[95:88] == 7'b1101101;
  assign _1180_ = state_in[95:88] == 7'b1101100;
  assign _1181_ = state_in[95:88] == 7'b1101011;
  assign _1182_ = state_in[95:88] == 7'b1101010;
  assign _1183_ = state_in[95:88] == 7'b1101001;
  assign _1184_ = state_in[95:88] == 7'b1101000;
  assign _1185_ = state_in[95:88] == 7'b1100111;
  assign _1186_ = state_in[95:88] == 7'b1100110;
  assign _1187_ = state_in[95:88] == 7'b1100101;
  assign _1188_ = state_in[95:88] == 7'b1100100;
  assign _1189_ = state_in[95:88] == 7'b1100011;
  assign _1190_ = state_in[95:88] == 7'b1100010;
  assign _1191_ = state_in[95:88] == 7'b1100001;
  assign _1192_ = state_in[95:88] == 7'b1100000;
  assign _1193_ = state_in[95:88] == 7'b1011111;
  assign _1194_ = state_in[95:88] == 7'b1011110;
  assign _1195_ = state_in[95:88] == 7'b1011101;
  assign _1196_ = state_in[95:88] == 7'b1011100;
  assign _1197_ = state_in[95:88] == 7'b1011011;
  assign _1198_ = state_in[95:88] == 7'b1011010;
  assign _1199_ = state_in[95:88] == 7'b1011001;
  assign _1200_ = state_in[95:88] == 7'b1011000;
  assign _1201_ = state_in[95:88] == 7'b1010111;
  assign _1202_ = state_in[95:88] == 7'b1010110;
  assign _1203_ = state_in[95:88] == 7'b1010101;
  assign _1204_ = state_in[95:88] == 7'b1010100;
  assign _1205_ = state_in[95:88] == 7'b1010011;
  assign _1206_ = state_in[95:88] == 7'b1010010;
  assign _1207_ = state_in[95:88] == 7'b1010001;
  assign _1208_ = state_in[95:88] == 7'b1010000;
  assign _1209_ = state_in[95:88] == 7'b1001111;
  assign _1210_ = state_in[95:88] == 7'b1001110;
  assign _1211_ = state_in[95:88] == 7'b1001101;
  assign _1212_ = state_in[95:88] == 7'b1001100;
  assign _1213_ = state_in[95:88] == 7'b1001011;
  assign _1214_ = state_in[95:88] == 7'b1001010;
  assign _1215_ = state_in[95:88] == 7'b1001001;
  assign _1216_ = state_in[95:88] == 7'b1001000;
  assign _1217_ = state_in[95:88] == 7'b1000111;
  assign _1218_ = state_in[95:88] == 7'b1000110;
  assign _1219_ = state_in[95:88] == 7'b1000101;
  assign _1220_ = state_in[95:88] == 7'b1000100;
  assign _1221_ = state_in[95:88] == 7'b1000011;
  assign _1222_ = state_in[95:88] == 7'b1000010;
  assign _1223_ = state_in[95:88] == 7'b1000001;
  assign _1224_ = state_in[95:88] == 7'b1000000;
  assign _1225_ = state_in[95:88] == 6'b111111;
  assign _1226_ = state_in[95:88] == 6'b111110;
  assign _1227_ = state_in[95:88] == 6'b111101;
  assign _1228_ = state_in[95:88] == 6'b111100;
  assign _1229_ = state_in[95:88] == 6'b111011;
  assign _1230_ = state_in[95:88] == 6'b111010;
  assign _1231_ = state_in[95:88] == 6'b111001;
  assign _1232_ = state_in[95:88] == 6'b111000;
  assign _1233_ = state_in[95:88] == 6'b110111;
  assign _1234_ = state_in[95:88] == 6'b110110;
  assign _1235_ = state_in[95:88] == 6'b110101;
  assign _1236_ = state_in[95:88] == 6'b110100;
  assign _1237_ = state_in[95:88] == 6'b110011;
  assign _1238_ = state_in[95:88] == 6'b110010;
  assign _1239_ = state_in[95:88] == 6'b110001;
  assign _1240_ = state_in[95:88] == 6'b110000;
  assign _1241_ = state_in[95:88] == 6'b101111;
  assign _1242_ = state_in[95:88] == 6'b101110;
  assign _1243_ = state_in[95:88] == 6'b101101;
  assign _1244_ = state_in[95:88] == 6'b101100;
  assign _1245_ = state_in[95:88] == 6'b101011;
  assign _1246_ = state_in[95:88] == 6'b101010;
  assign _1247_ = state_in[95:88] == 6'b101001;
  assign _1248_ = state_in[95:88] == 6'b101000;
  assign _1249_ = state_in[95:88] == 6'b100111;
  assign _1250_ = state_in[95:88] == 6'b100110;
  assign _1251_ = state_in[95:88] == 6'b100101;
  assign _1252_ = state_in[95:88] == 6'b100100;
  assign _1253_ = state_in[95:88] == 6'b100011;
  assign _1254_ = state_in[95:88] == 6'b100010;
  assign _1255_ = state_in[95:88] == 6'b100001;
  assign _1256_ = state_in[95:88] == 6'b100000;
  assign _1257_ = state_in[95:88] == 5'b11111;
  assign _1258_ = state_in[95:88] == 5'b11110;
  assign _1259_ = state_in[95:88] == 5'b11101;
  assign _1260_ = state_in[95:88] == 5'b11100;
  assign _1261_ = state_in[95:88] == 5'b11011;
  assign _1262_ = state_in[95:88] == 5'b11010;
  assign _1263_ = state_in[95:88] == 5'b11001;
  assign _1264_ = state_in[95:88] == 5'b11000;
  assign _1265_ = state_in[95:88] == 5'b10111;
  assign _1266_ = state_in[95:88] == 5'b10110;
  assign _1267_ = state_in[95:88] == 5'b10101;
  assign _1268_ = state_in[95:88] == 5'b10100;
  assign _1269_ = state_in[95:88] == 5'b10011;
  assign _1270_ = state_in[95:88] == 5'b10010;
  assign _1271_ = state_in[95:88] == 5'b10001;
  assign _1272_ = state_in[95:88] == 5'b10000;
  assign _1273_ = state_in[95:88] == 4'b1111;
  assign _1274_ = state_in[95:88] == 4'b1110;
  assign _1275_ = state_in[95:88] == 4'b1101;
  assign _1276_ = state_in[95:88] == 4'b1100;
  assign _1277_ = state_in[95:88] == 4'b1011;
  assign _1278_ = state_in[95:88] == 4'b1010;
  assign _1279_ = state_in[95:88] == 4'b1001;
  assign _1280_ = state_in[95:88] == 4'b1000;
  assign _1281_ = state_in[95:88] == 3'b111;
  assign _1282_ = state_in[95:88] == 3'b110;
  assign _1283_ = state_in[95:88] == 3'b101;
  assign _1284_ = state_in[95:88] == 3'b100;
  assign _1285_ = state_in[95:88] == 2'b11;
  assign _1286_ = state_in[95:88] == 2'b10;
  assign _1287_ = state_in[95:88] == 1'b1;
  assign _1288_ = ! state_in[95:88];
  always @(posedge clk)
      \t1.t0.s4.out <= _1289_;
  wire [255:0] fangyuan10;
  assign fangyuan10 = { _1288_, _1287_, _1286_, _1285_, _1284_, _1283_, _1282_, _1281_, _1280_, _1279_, _1278_, _1277_, _1276_, _1275_, _1274_, _1273_, _1272_, _1271_, _1270_, _1269_, _1268_, _1267_, _1266_, _1265_, _1264_, _1263_, _1262_, _1261_, _1260_, _1259_, _1258_, _1257_, _1256_, _1255_, _1254_, _1253_, _1252_, _1251_, _1250_, _1249_, _1248_, _1247_, _1246_, _1245_, _1244_, _1243_, _1242_, _1241_, _1240_, _1239_, _1238_, _1237_, _1236_, _1235_, _1234_, _1233_, _1232_, _1231_, _1230_, _1229_, _1228_, _1227_, _1226_, _1225_, _1224_, _1223_, _1222_, _1221_, _1220_, _1219_, _1218_, _1217_, _1216_, _1215_, _1214_, _1213_, _1212_, _1211_, _1210_, _1209_, _1208_, _1207_, _1206_, _1205_, _1204_, _1203_, _1202_, _1201_, _1200_, _1199_, _1198_, _1197_, _1196_, _1195_, _1194_, _1193_, _1192_, _1191_, _1190_, _1189_, _1188_, _1187_, _1186_, _1185_, _1184_, _1183_, _1182_, _1181_, _1180_, _1179_, _1178_, _1177_, _1176_, _1175_, _1174_, _1173_, _1172_, _1171_, _1170_, _1169_, _1168_, _1167_, _1166_, _1165_, _1164_, _1163_, _1162_, _1161_, _1160_, _1159_, _1158_, _1157_, _1156_, _1155_, _1154_, _1153_, _1152_, _1151_, _1150_, _1149_, _1148_, _1147_, _1146_, _1145_, _1144_, _1143_, _1142_, _1141_, _1140_, _1139_, _1138_, _1137_, _1136_, _1135_, _1134_, _1133_, _1132_, _1131_, _1130_, _1129_, _1128_, _1127_, _1126_, _1125_, _1124_, _1123_, _1122_, _1121_, _1120_, _1119_, _1118_, _1117_, _1116_, _1115_, _1114_, _1113_, _1112_, _1111_, _1110_, _1109_, _1108_, _1107_, _1106_, _1105_, _1104_, _1103_, _1102_, _1101_, _1100_, _1099_, _1098_, _1097_, _1096_, _1095_, _1094_, _1093_, _1092_, _1091_, _1090_, _1089_, _1088_, _1087_, _1086_, _1085_, _1084_, _1083_, _1082_, _1081_, _1080_, _1079_, _1078_, _1077_, _1076_, _1075_, _1074_, _1073_, _1072_, _1071_, _1070_, _1069_, _1068_, _1067_, _1066_, _1065_, _1064_, _1063_, _1062_, _1061_, _1060_, _1059_, _1058_, _1057_, _1056_, _1055_, _1054_, _1053_, _1052_, _1051_, _1050_, _1049_, _1048_, _1047_, _1046_, _1045_, _1044_, _1043_, _1042_, _1041_, _1040_, _1039_, _1038_, _1037_, _1036_, _1035_, _1034_, _1033_ };

  always @(\t1.t0.s4.out or fangyuan10) begin
    casez (fangyuan10)
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1 :
        _1289_ = 8'b00101100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1? :
        _1289_ = 8'b01101101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?? :
        _1289_ = 8'b10101000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??? :
        _1289_ = 8'b01111011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???? :
        _1289_ = 8'b00011110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????? :
        _1289_ = 8'b01011010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????? :
        _1289_ = 8'b00101001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????? :
        _1289_ = 8'b10000010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????? :
        _1289_ = 8'b11010000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????? :
        _1289_ = 8'b10000100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????? :
        _1289_ = 8'b11010111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????? :
        _1289_ = 8'b01100101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????? :
        _1289_ = 8'b00011010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????? :
        _1289_ = 8'b00001001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????? :
        _1289_ = 8'b01011001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????? :
        _1289_ = 8'b00000011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????? :
        _1289_ = 8'b10100101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????? :
        _1289_ = 8'b01010000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????? :
        _1289_ = 8'b10101010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????? :
        _1289_ = 8'b10000111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????? :
        _1289_ = 8'b11001001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????? :
        _1289_ = 8'b00010101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????? :
        _1289_ = 8'b00111100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????? :
        _1289_ = 8'b00101101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????? :
        _1289_ = 8'b00110011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????? :
        _1289_ = 8'b00000111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????? :
        _1289_ = 8'b10101001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????? :
        _1289_ = 8'b11010010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????? :
        _1289_ = 8'b00100010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????? :
        _1289_ = 8'b00101011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????? :
        _1289_ = 8'b11101011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????? :
        _1289_ = 8'b11011001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????? :
        _1289_ = 8'b00100111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????? :
        _1289_ = 8'b00111010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????? :
        _1289_ = 8'b10011001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????? :
        _1289_ = 8'b00010111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????? :
        _1289_ = 8'b01101001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????? :
        _1289_ = 8'b10101110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????? :
        _1289_ = 8'b01101010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????? :
        _1289_ = 8'b11000010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????? :
        _1289_ = 8'b00011100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????? :
        _1289_ = 8'b11110111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????? :
        _1289_ = 8'b00000110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????? :
        _1289_ = 8'b10010000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????? :
        _1289_ = 8'b11001100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????? :
        _1289_ = 8'b01110001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????? :
        _1289_ = 8'b01111100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????? :
        _1289_ = 8'b11100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????? :
        _1289_ = 8'b00001111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????? :
        _1289_ = 8'b00001101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????? :
        _1289_ = 8'b01100001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????? :
        _1289_ = 8'b10010110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????? :
        _1289_ = 8'b00111110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????? :
        _1289_ = 8'b11101000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????? :
        _1289_ = 8'b10100001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????? :
        _1289_ = 8'b11001011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????? :
        _1289_ = 8'b10010111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????? :
        _1289_ = 8'b01110011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????? :
        _1289_ = 8'b01010111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????? :
        _1289_ = 8'b00111000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????? :
        _1289_ = 8'b01011100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????? :
        _1289_ = 8'b01001010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????? :
        _1289_ = 8'b11110000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????? :
        _1289_ = 8'b01101111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????? :
        _1289_ = 8'b00010000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b01000111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b11110100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b11001010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b11001111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b11110011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b10101100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b11011000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b01001001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b10011100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b10110001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b00000001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b11011010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b01101110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b10001011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b11010101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b11110010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b11010011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b00110001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b00111001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b11000100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b01000011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b10111101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b10011111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b10111000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b01001000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b00001100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b10010010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b00010100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b01110100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b01100100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b11011011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b10101101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b00010110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b10111100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b10100111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b00101000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b01101011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b11000111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b10001100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b00001011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b00111011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b01010100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b01000100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b10100011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b10011110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b00011001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b11000000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b11100110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b00110010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b10111010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b11001000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b01111010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b11111100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b01010101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b10010011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b00101110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b10001000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b00110101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b10111110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b11000011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b00100110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b00011000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b10000001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b10111111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b11111101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b11100101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b00100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b01000010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b10101111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b01110111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b01100011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b11110001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b01110000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b00100001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b00111111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b00000101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b10000000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b01011101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b10100010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b01001011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b00100101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b01111000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b10100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b11111110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b00000100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b11101001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b10001010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b00010001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b01100110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b10011010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b10000110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b11101101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b01001111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b11000101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b10111011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b10000101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b10110000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b10011000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b10010100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b01110010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b01100111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b10001101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b11010100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b10110110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b01111001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b11100011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b01000000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b11000001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b00000000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b10111001 ;
      256'b????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b10100110 ;
      256'b???????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b00010011 ;
      256'b??????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b01011110 ;
      256'b?????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b11011101 ;
      256'b????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b01010010 ;
      256'b???????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b01111101 ;
      256'b??????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b10110111 ;
      256'b?????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b01110110 ;
      256'b????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b10100100 ;
      256'b???????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b01011011 ;
      256'b??????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b10110100 ;
      256'b?????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b11011100 ;
      256'b????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b00110110 ;
      256'b???????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b00110100 ;
      256'b??????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b01011000 ;
      256'b?????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b00011101 ;
      256'b????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b00010010 ;
      256'b???????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b11101010 ;
      256'b??????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b01111111 ;
      256'b?????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b01001110 ;
      256'b????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b11001101 ;
      256'b???????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b11011111 ;
      256'b??????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b00011011 ;
      256'b?????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b00100100 ;
      256'b????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b00001110 ;
      256'b???????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b00101111 ;
      256'b??????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b00001010 ;
      256'b?????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b00110111 ;
      256'b????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b00110000 ;
      256'b???????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b10011101 ;
      256'b??????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b01000110 ;
      256'b?????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b10010101 ;
      256'b????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b00001000 ;
      256'b???????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b00101010 ;
      256'b??????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b01100010 ;
      256'b?????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b10101011 ;
      256'b????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b11100010 ;
      256'b???????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b11111001 ;
      256'b??????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b11010001 ;
      256'b?????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b01010001 ;
      256'b????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b01101000 ;
      256'b???????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b10000011 ;
      256'b??????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b11110101 ;
      256'b?????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b01111110 ;
      256'b????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b01101100 ;
      256'b???????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b01001100 ;
      256'b??????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b00111101 ;
      256'b?????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b11100001 ;
      256'b????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b01110101 ;
      256'b???????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b10011011 ;
      256'b??????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b11100100 ;
      256'b?????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b01010011 ;
      256'b????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b00100011 ;
      256'b???????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b01000101 ;
      256'b??????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b01011111 ;
      256'b?????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b10110011 ;
      256'b????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b01000001 ;
      256'b???????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b11111011 ;
      256'b??????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b10001110 ;
      256'b?????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b10110010 ;
      256'b????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b11101111 ;
      256'b???????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b11111010 ;
      256'b??????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b10001001 ;
      256'b?????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b00011111 ;
      256'b????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b10001111 ;
      256'b???????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b11101100 ;
      256'b??????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b01001101 ;
      256'b?????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b10110101 ;
      256'b????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b11100111 ;
      256'b???????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b01010110 ;
      256'b??????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b11001110 ;
      256'b?????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b00000010 ;
      256'b????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b01100000 ;
      256'b???????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b10010001 ;
      256'b??????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b11011110 ;
      256'b?????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b11010110 ;
      256'b????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b11111111 ;
      256'b???1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b11110110 ;
      256'b??1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b11101110 ;
      256'b?1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b11111000 ;
      256'b1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b11000110 ;
      default:
        _1289_ = \t1.t0.s4.out ;
    endcase
  end
  assign p11[31:24] = \t1.t1.s0.out ^ \t1.t1.s4.out ;
  always @(posedge clk)
      \t1.t1.s0.out <= _1290_;
  wire [255:0] fangyuan11;
  assign fangyuan11 = { _1546_, _1545_, _1544_, _1543_, _1542_, _1541_, _1540_, _1539_, _1538_, _1537_, _1536_, _1535_, _1534_, _1533_, _1532_, _1531_, _1530_, _1529_, _1528_, _1527_, _1526_, _1525_, _1524_, _1523_, _1522_, _1521_, _1520_, _1519_, _1518_, _1517_, _1516_, _1515_, _1514_, _1513_, _1512_, _1511_, _1510_, _1509_, _1508_, _1507_, _1506_, _1505_, _1504_, _1503_, _1502_, _1501_, _1500_, _1499_, _1498_, _1497_, _1496_, _1495_, _1494_, _1493_, _1492_, _1491_, _1490_, _1489_, _1488_, _1487_, _1486_, _1485_, _1484_, _1483_, _1482_, _1481_, _1480_, _1479_, _1478_, _1477_, _1476_, _1475_, _1474_, _1473_, _1472_, _1471_, _1470_, _1469_, _1468_, _1467_, _1466_, _1465_, _1464_, _1463_, _1462_, _1461_, _1460_, _1459_, _1458_, _1457_, _1456_, _1455_, _1454_, _1453_, _1452_, _1451_, _1450_, _1449_, _1448_, _1447_, _1446_, _1445_, _1444_, _1443_, _1442_, _1441_, _1440_, _1439_, _1438_, _1437_, _1436_, _1435_, _1434_, _1433_, _1432_, _1431_, _1430_, _1429_, _1428_, _1427_, _1426_, _1425_, _1424_, _1423_, _1422_, _1421_, _1420_, _1419_, _1418_, _1417_, _1416_, _1415_, _1414_, _1413_, _1412_, _1411_, _1410_, _1409_, _1408_, _1407_, _1406_, _1405_, _1404_, _1403_, _1402_, _1401_, _1400_, _1399_, _1398_, _1397_, _1396_, _1395_, _1394_, _1393_, _1392_, _1391_, _1390_, _1389_, _1388_, _1387_, _1386_, _1385_, _1384_, _1383_, _1382_, _1381_, _1380_, _1379_, _1378_, _1377_, _1376_, _1375_, _1374_, _1373_, _1372_, _1371_, _1370_, _1369_, _1368_, _1367_, _1366_, _1365_, _1364_, _1363_, _1362_, _1361_, _1360_, _1359_, _1358_, _1357_, _1356_, _1355_, _1354_, _1353_, _1352_, _1351_, _1350_, _1349_, _1348_, _1347_, _1346_, _1345_, _1344_, _1343_, _1342_, _1341_, _1340_, _1339_, _1338_, _1337_, _1336_, _1335_, _1334_, _1333_, _1332_, _1331_, _1330_, _1329_, _1328_, _1327_, _1326_, _1325_, _1324_, _1323_, _1322_, _1321_, _1320_, _1319_, _1318_, _1317_, _1316_, _1315_, _1314_, _1313_, _1312_, _1311_, _1310_, _1309_, _1308_, _1307_, _1306_, _1305_, _1304_, _1303_, _1302_, _1301_, _1300_, _1299_, _1298_, _1297_, _1296_, _1295_, _1294_, _1293_, _1292_, _1291_ };

  always @(\t1.t1.s0.out or fangyuan11) begin
    casez (fangyuan11)
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1 :
        _1290_ = 8'b00010110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1? :
        _1290_ = 8'b10111011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?? :
        _1290_ = 8'b01010100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??? :
        _1290_ = 8'b10110000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???? :
        _1290_ = 8'b00001111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????? :
        _1290_ = 8'b00101101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????? :
        _1290_ = 8'b10011001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????? :
        _1290_ = 8'b01000001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????? :
        _1290_ = 8'b01101000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????? :
        _1290_ = 8'b01000010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????? :
        _1290_ = 8'b11100110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????? :
        _1290_ = 8'b10111111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????? :
        _1290_ = 8'b00001101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????? :
        _1290_ = 8'b10001001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????? :
        _1290_ = 8'b10100001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????? :
        _1290_ = 8'b10001100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????? :
        _1290_ = 8'b11011111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????? :
        _1290_ = 8'b00101000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????? :
        _1290_ = 8'b01010101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????? :
        _1290_ = 8'b11001110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????? :
        _1290_ = 8'b11101001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????? :
        _1290_ = 8'b10000111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????? :
        _1290_ = 8'b00011110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????? :
        _1290_ = 8'b10011011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????? :
        _1290_ = 8'b10010100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????? :
        _1290_ = 8'b10001110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????? :
        _1290_ = 8'b11011001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????? :
        _1290_ = 8'b01101001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????? :
        _1290_ = 8'b00010001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????? :
        _1290_ = 8'b10011000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????? :
        _1290_ = 8'b11111000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????? :
        _1290_ = 8'b11100001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????? :
        _1290_ = 8'b10011110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????? :
        _1290_ = 8'b00011101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????? :
        _1290_ = 8'b11000001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????? :
        _1290_ = 8'b10000110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????? :
        _1290_ = 8'b10111001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????? :
        _1290_ = 8'b01010111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????? :
        _1290_ = 8'b00110101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????? :
        _1290_ = 8'b01100001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????? :
        _1290_ = 8'b00001110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????? :
        _1290_ = 8'b11110110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????? :
        _1290_ = 8'b00000011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????? :
        _1290_ = 8'b01001000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????? :
        _1290_ = 8'b01100110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????? :
        _1290_ = 8'b10110101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????? :
        _1290_ = 8'b00111110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????? :
        _1290_ = 8'b01110000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????? :
        _1290_ = 8'b10001010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????? :
        _1290_ = 8'b10001011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????? :
        _1290_ = 8'b10111101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????? :
        _1290_ = 8'b01001011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????? :
        _1290_ = 8'b00011111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????? :
        _1290_ = 8'b01110100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????? :
        _1290_ = 8'b11011101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????? :
        _1290_ = 8'b11101000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????? :
        _1290_ = 8'b11000110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????? :
        _1290_ = 8'b10110100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????? :
        _1290_ = 8'b10100110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????? :
        _1290_ = 8'b00011100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????? :
        _1290_ = 8'b00101110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????? :
        _1290_ = 8'b00100101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????? :
        _1290_ = 8'b01111000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????? :
        _1290_ = 8'b10111010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????? :
        _1290_ = 8'b00001000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b10101110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b01111010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b01100101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b11101010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b11110100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b01010110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b01101100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b10101001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b01001110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b11010101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b10001101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b01101101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b00110111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b11001000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b11100111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b01111001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b11100100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b10010101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b10010001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b01100010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b10101100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b11010011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b11000010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b01011100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b00100100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b00000110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b01001001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b00001010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b00111010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b00110010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b11100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b11011011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b00001011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b01011110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b11011110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b00010100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b10111000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b11101110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b01000110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b10001000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b10010000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b00101010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b00100010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b11011100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b01001111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b10000001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b01100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b01110011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b00011001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b01011101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b01100100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b00111101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b01111110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b10100111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b11000100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b00010111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b01000100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b10010111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b01011111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b11101100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b00010011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b00001100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b11001101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b11010010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b11110011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b11111111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b00010000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b00100001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b11011010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b10110110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b10111100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b11110101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b00111000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b10011101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b10010010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b10001111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b01000000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b10100011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b01010001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b10101000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b10011111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b00111100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b01010000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b01111111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b00000010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b11111001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b01000101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b10000101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b00110011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b01001101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b01000011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b11111011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b10101010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b11101111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b11010000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b11001111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b01011000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b01001100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b01001010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b00111001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b10111110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b11001011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b01101010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b01011011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b10110001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b11111100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b00100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b11101101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b00000000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b11010001 ;
      256'b????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b01010011 ;
      256'b???????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b10000100 ;
      256'b??????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b00101111 ;
      256'b?????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b11100011 ;
      256'b????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b00101001 ;
      256'b???????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b10110011 ;
      256'b??????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b11010110 ;
      256'b?????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b00111011 ;
      256'b????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b01010010 ;
      256'b???????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b10100000 ;
      256'b??????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b01011010 ;
      256'b?????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b01101110 ;
      256'b????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b00011011 ;
      256'b???????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b00011010 ;
      256'b??????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b00101100 ;
      256'b?????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b10000011 ;
      256'b????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b00001001 ;
      256'b???????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b01110101 ;
      256'b??????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b10110010 ;
      256'b?????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b00100111 ;
      256'b????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b11101011 ;
      256'b???????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b11100010 ;
      256'b??????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b10000000 ;
      256'b?????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b00010010 ;
      256'b????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b00000111 ;
      256'b???????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b10011010 ;
      256'b??????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b00000101 ;
      256'b?????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b10010110 ;
      256'b????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b00011000 ;
      256'b???????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b11000011 ;
      256'b??????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b00100011 ;
      256'b?????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b11000111 ;
      256'b????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b00000100 ;
      256'b???????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b00010101 ;
      256'b??????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b00110001 ;
      256'b?????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b11011000 ;
      256'b????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b01110001 ;
      256'b???????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b11110001 ;
      256'b??????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b11100101 ;
      256'b?????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b10100101 ;
      256'b????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b00110100 ;
      256'b???????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b11001100 ;
      256'b??????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b11110111 ;
      256'b?????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b00111111 ;
      256'b????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b00110110 ;
      256'b???????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b00100110 ;
      256'b??????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b10010011 ;
      256'b?????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b11111101 ;
      256'b????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b10110111 ;
      256'b???????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b11000000 ;
      256'b??????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b01110010 ;
      256'b?????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b10100100 ;
      256'b????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b10011100 ;
      256'b???????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b10101111 ;
      256'b??????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b10100010 ;
      256'b?????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b11010100 ;
      256'b????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b10101101 ;
      256'b???????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b11110000 ;
      256'b??????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b01000111 ;
      256'b?????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b01011001 ;
      256'b????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b11111010 ;
      256'b???????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b01111101 ;
      256'b??????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b11001001 ;
      256'b?????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b10000010 ;
      256'b????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b11001010 ;
      256'b???????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b01110110 ;
      256'b??????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b10101011 ;
      256'b?????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b11010111 ;
      256'b????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b11111110 ;
      256'b???????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b00101011 ;
      256'b??????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b01100111 ;
      256'b?????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b00000001 ;
      256'b????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b00110000 ;
      256'b???????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b11000101 ;
      256'b??????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b01101111 ;
      256'b?????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b01101011 ;
      256'b????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b11110010 ;
      256'b???1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b01111011 ;
      256'b??1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b01110111 ;
      256'b?1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b01111100 ;
      256'b1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b01100011 ;
      default:
        _1290_ = \t1.t1.s0.out ;
    endcase
  end
  assign _1291_ = state_in[87:80] == 8'b11111111;
  assign _1292_ = state_in[87:80] == 8'b11111110;
  assign _1293_ = state_in[87:80] == 8'b11111101;
  assign _1294_ = state_in[87:80] == 8'b11111100;
  assign _1295_ = state_in[87:80] == 8'b11111011;
  assign _1296_ = state_in[87:80] == 8'b11111010;
  assign _1297_ = state_in[87:80] == 8'b11111001;
  assign _1298_ = state_in[87:80] == 8'b11111000;
  assign _1299_ = state_in[87:80] == 8'b11110111;
  assign _1300_ = state_in[87:80] == 8'b11110110;
  assign _1301_ = state_in[87:80] == 8'b11110101;
  assign _1302_ = state_in[87:80] == 8'b11110100;
  assign _1303_ = state_in[87:80] == 8'b11110011;
  assign _1304_ = state_in[87:80] == 8'b11110010;
  assign _1305_ = state_in[87:80] == 8'b11110001;
  assign _1306_ = state_in[87:80] == 8'b11110000;
  assign _1307_ = state_in[87:80] == 8'b11101111;
  assign _1308_ = state_in[87:80] == 8'b11101110;
  assign _1309_ = state_in[87:80] == 8'b11101101;
  assign _1310_ = state_in[87:80] == 8'b11101100;
  assign _1311_ = state_in[87:80] == 8'b11101011;
  assign _1312_ = state_in[87:80] == 8'b11101010;
  assign _1313_ = state_in[87:80] == 8'b11101001;
  assign _1314_ = state_in[87:80] == 8'b11101000;
  assign _1315_ = state_in[87:80] == 8'b11100111;
  assign _1316_ = state_in[87:80] == 8'b11100110;
  assign _1317_ = state_in[87:80] == 8'b11100101;
  assign _1318_ = state_in[87:80] == 8'b11100100;
  assign _1319_ = state_in[87:80] == 8'b11100011;
  assign _1320_ = state_in[87:80] == 8'b11100010;
  assign _1321_ = state_in[87:80] == 8'b11100001;
  assign _1322_ = state_in[87:80] == 8'b11100000;
  assign _1323_ = state_in[87:80] == 8'b11011111;
  assign _1324_ = state_in[87:80] == 8'b11011110;
  assign _1325_ = state_in[87:80] == 8'b11011101;
  assign _1326_ = state_in[87:80] == 8'b11011100;
  assign _1327_ = state_in[87:80] == 8'b11011011;
  assign _1328_ = state_in[87:80] == 8'b11011010;
  assign _1329_ = state_in[87:80] == 8'b11011001;
  assign _1330_ = state_in[87:80] == 8'b11011000;
  assign _1331_ = state_in[87:80] == 8'b11010111;
  assign _1332_ = state_in[87:80] == 8'b11010110;
  assign _1333_ = state_in[87:80] == 8'b11010101;
  assign _1334_ = state_in[87:80] == 8'b11010100;
  assign _1335_ = state_in[87:80] == 8'b11010011;
  assign _1336_ = state_in[87:80] == 8'b11010010;
  assign _1337_ = state_in[87:80] == 8'b11010001;
  assign _1338_ = state_in[87:80] == 8'b11010000;
  assign _1339_ = state_in[87:80] == 8'b11001111;
  assign _1340_ = state_in[87:80] == 8'b11001110;
  assign _1341_ = state_in[87:80] == 8'b11001101;
  assign _1342_ = state_in[87:80] == 8'b11001100;
  assign _1343_ = state_in[87:80] == 8'b11001011;
  assign _1344_ = state_in[87:80] == 8'b11001010;
  assign _1345_ = state_in[87:80] == 8'b11001001;
  assign _1346_ = state_in[87:80] == 8'b11001000;
  assign _1347_ = state_in[87:80] == 8'b11000111;
  assign _1348_ = state_in[87:80] == 8'b11000110;
  assign _1349_ = state_in[87:80] == 8'b11000101;
  assign _1350_ = state_in[87:80] == 8'b11000100;
  assign _1351_ = state_in[87:80] == 8'b11000011;
  assign _1352_ = state_in[87:80] == 8'b11000010;
  assign _1353_ = state_in[87:80] == 8'b11000001;
  assign _1354_ = state_in[87:80] == 8'b11000000;
  assign _1355_ = state_in[87:80] == 8'b10111111;
  assign _1356_ = state_in[87:80] == 8'b10111110;
  assign _1357_ = state_in[87:80] == 8'b10111101;
  assign _1358_ = state_in[87:80] == 8'b10111100;
  assign _1359_ = state_in[87:80] == 8'b10111011;
  assign _1360_ = state_in[87:80] == 8'b10111010;
  assign _1361_ = state_in[87:80] == 8'b10111001;
  assign _1362_ = state_in[87:80] == 8'b10111000;
  assign _1363_ = state_in[87:80] == 8'b10110111;
  assign _1364_ = state_in[87:80] == 8'b10110110;
  assign _1365_ = state_in[87:80] == 8'b10110101;
  assign _1366_ = state_in[87:80] == 8'b10110100;
  assign _1367_ = state_in[87:80] == 8'b10110011;
  assign _1368_ = state_in[87:80] == 8'b10110010;
  assign _1369_ = state_in[87:80] == 8'b10110001;
  assign _1370_ = state_in[87:80] == 8'b10110000;
  assign _1371_ = state_in[87:80] == 8'b10101111;
  assign _1372_ = state_in[87:80] == 8'b10101110;
  assign _1373_ = state_in[87:80] == 8'b10101101;
  assign _1374_ = state_in[87:80] == 8'b10101100;
  assign _1375_ = state_in[87:80] == 8'b10101011;
  assign _1376_ = state_in[87:80] == 8'b10101010;
  assign _1377_ = state_in[87:80] == 8'b10101001;
  assign _1378_ = state_in[87:80] == 8'b10101000;
  assign _1379_ = state_in[87:80] == 8'b10100111;
  assign _1380_ = state_in[87:80] == 8'b10100110;
  assign _1381_ = state_in[87:80] == 8'b10100101;
  assign _1382_ = state_in[87:80] == 8'b10100100;
  assign _1383_ = state_in[87:80] == 8'b10100011;
  assign _1384_ = state_in[87:80] == 8'b10100010;
  assign _1385_ = state_in[87:80] == 8'b10100001;
  assign _1386_ = state_in[87:80] == 8'b10100000;
  assign _1387_ = state_in[87:80] == 8'b10011111;
  assign _1388_ = state_in[87:80] == 8'b10011110;
  assign _1389_ = state_in[87:80] == 8'b10011101;
  assign _1390_ = state_in[87:80] == 8'b10011100;
  assign _1391_ = state_in[87:80] == 8'b10011011;
  assign _1392_ = state_in[87:80] == 8'b10011010;
  assign _1393_ = state_in[87:80] == 8'b10011001;
  assign _1394_ = state_in[87:80] == 8'b10011000;
  assign _1395_ = state_in[87:80] == 8'b10010111;
  assign _1396_ = state_in[87:80] == 8'b10010110;
  assign _1397_ = state_in[87:80] == 8'b10010101;
  assign _1398_ = state_in[87:80] == 8'b10010100;
  assign _1399_ = state_in[87:80] == 8'b10010011;
  assign _1400_ = state_in[87:80] == 8'b10010010;
  assign _1401_ = state_in[87:80] == 8'b10010001;
  assign _1402_ = state_in[87:80] == 8'b10010000;
  assign _1403_ = state_in[87:80] == 8'b10001111;
  assign _1404_ = state_in[87:80] == 8'b10001110;
  assign _1405_ = state_in[87:80] == 8'b10001101;
  assign _1406_ = state_in[87:80] == 8'b10001100;
  assign _1407_ = state_in[87:80] == 8'b10001011;
  assign _1408_ = state_in[87:80] == 8'b10001010;
  assign _1409_ = state_in[87:80] == 8'b10001001;
  assign _1410_ = state_in[87:80] == 8'b10001000;
  assign _1411_ = state_in[87:80] == 8'b10000111;
  assign _1412_ = state_in[87:80] == 8'b10000110;
  assign _1413_ = state_in[87:80] == 8'b10000101;
  assign _1414_ = state_in[87:80] == 8'b10000100;
  assign _1415_ = state_in[87:80] == 8'b10000011;
  assign _1416_ = state_in[87:80] == 8'b10000010;
  assign _1417_ = state_in[87:80] == 8'b10000001;
  assign _1418_ = state_in[87:80] == 8'b10000000;
  assign _1419_ = state_in[87:80] == 7'b1111111;
  assign _1420_ = state_in[87:80] == 7'b1111110;
  assign _1421_ = state_in[87:80] == 7'b1111101;
  assign _1422_ = state_in[87:80] == 7'b1111100;
  assign _1423_ = state_in[87:80] == 7'b1111011;
  assign _1424_ = state_in[87:80] == 7'b1111010;
  assign _1425_ = state_in[87:80] == 7'b1111001;
  assign _1426_ = state_in[87:80] == 7'b1111000;
  assign _1427_ = state_in[87:80] == 7'b1110111;
  assign _1428_ = state_in[87:80] == 7'b1110110;
  assign _1429_ = state_in[87:80] == 7'b1110101;
  assign _1430_ = state_in[87:80] == 7'b1110100;
  assign _1431_ = state_in[87:80] == 7'b1110011;
  assign _1432_ = state_in[87:80] == 7'b1110010;
  assign _1433_ = state_in[87:80] == 7'b1110001;
  assign _1434_ = state_in[87:80] == 7'b1110000;
  assign _1435_ = state_in[87:80] == 7'b1101111;
  assign _1436_ = state_in[87:80] == 7'b1101110;
  assign _1437_ = state_in[87:80] == 7'b1101101;
  assign _1438_ = state_in[87:80] == 7'b1101100;
  assign _1439_ = state_in[87:80] == 7'b1101011;
  assign _1440_ = state_in[87:80] == 7'b1101010;
  assign _1441_ = state_in[87:80] == 7'b1101001;
  assign _1442_ = state_in[87:80] == 7'b1101000;
  assign _1443_ = state_in[87:80] == 7'b1100111;
  assign _1444_ = state_in[87:80] == 7'b1100110;
  assign _1445_ = state_in[87:80] == 7'b1100101;
  assign _1446_ = state_in[87:80] == 7'b1100100;
  assign _1447_ = state_in[87:80] == 7'b1100011;
  assign _1448_ = state_in[87:80] == 7'b1100010;
  assign _1449_ = state_in[87:80] == 7'b1100001;
  assign _1450_ = state_in[87:80] == 7'b1100000;
  assign _1451_ = state_in[87:80] == 7'b1011111;
  assign _1452_ = state_in[87:80] == 7'b1011110;
  assign _1453_ = state_in[87:80] == 7'b1011101;
  assign _1454_ = state_in[87:80] == 7'b1011100;
  assign _1455_ = state_in[87:80] == 7'b1011011;
  assign _1456_ = state_in[87:80] == 7'b1011010;
  assign _1457_ = state_in[87:80] == 7'b1011001;
  assign _1458_ = state_in[87:80] == 7'b1011000;
  assign _1459_ = state_in[87:80] == 7'b1010111;
  assign _1460_ = state_in[87:80] == 7'b1010110;
  assign _1461_ = state_in[87:80] == 7'b1010101;
  assign _1462_ = state_in[87:80] == 7'b1010100;
  assign _1463_ = state_in[87:80] == 7'b1010011;
  assign _1464_ = state_in[87:80] == 7'b1010010;
  assign _1465_ = state_in[87:80] == 7'b1010001;
  assign _1466_ = state_in[87:80] == 7'b1010000;
  assign _1467_ = state_in[87:80] == 7'b1001111;
  assign _1468_ = state_in[87:80] == 7'b1001110;
  assign _1469_ = state_in[87:80] == 7'b1001101;
  assign _1470_ = state_in[87:80] == 7'b1001100;
  assign _1471_ = state_in[87:80] == 7'b1001011;
  assign _1472_ = state_in[87:80] == 7'b1001010;
  assign _1473_ = state_in[87:80] == 7'b1001001;
  assign _1474_ = state_in[87:80] == 7'b1001000;
  assign _1475_ = state_in[87:80] == 7'b1000111;
  assign _1476_ = state_in[87:80] == 7'b1000110;
  assign _1477_ = state_in[87:80] == 7'b1000101;
  assign _1478_ = state_in[87:80] == 7'b1000100;
  assign _1479_ = state_in[87:80] == 7'b1000011;
  assign _1480_ = state_in[87:80] == 7'b1000010;
  assign _1481_ = state_in[87:80] == 7'b1000001;
  assign _1482_ = state_in[87:80] == 7'b1000000;
  assign _1483_ = state_in[87:80] == 6'b111111;
  assign _1484_ = state_in[87:80] == 6'b111110;
  assign _1485_ = state_in[87:80] == 6'b111101;
  assign _1486_ = state_in[87:80] == 6'b111100;
  assign _1487_ = state_in[87:80] == 6'b111011;
  assign _1488_ = state_in[87:80] == 6'b111010;
  assign _1489_ = state_in[87:80] == 6'b111001;
  assign _1490_ = state_in[87:80] == 6'b111000;
  assign _1491_ = state_in[87:80] == 6'b110111;
  assign _1492_ = state_in[87:80] == 6'b110110;
  assign _1493_ = state_in[87:80] == 6'b110101;
  assign _1494_ = state_in[87:80] == 6'b110100;
  assign _1495_ = state_in[87:80] == 6'b110011;
  assign _1496_ = state_in[87:80] == 6'b110010;
  assign _1497_ = state_in[87:80] == 6'b110001;
  assign _1498_ = state_in[87:80] == 6'b110000;
  assign _1499_ = state_in[87:80] == 6'b101111;
  assign _1500_ = state_in[87:80] == 6'b101110;
  assign _1501_ = state_in[87:80] == 6'b101101;
  assign _1502_ = state_in[87:80] == 6'b101100;
  assign _1503_ = state_in[87:80] == 6'b101011;
  assign _1504_ = state_in[87:80] == 6'b101010;
  assign _1505_ = state_in[87:80] == 6'b101001;
  assign _1506_ = state_in[87:80] == 6'b101000;
  assign _1507_ = state_in[87:80] == 6'b100111;
  assign _1508_ = state_in[87:80] == 6'b100110;
  assign _1509_ = state_in[87:80] == 6'b100101;
  assign _1510_ = state_in[87:80] == 6'b100100;
  assign _1511_ = state_in[87:80] == 6'b100011;
  assign _1512_ = state_in[87:80] == 6'b100010;
  assign _1513_ = state_in[87:80] == 6'b100001;
  assign _1514_ = state_in[87:80] == 6'b100000;
  assign _1515_ = state_in[87:80] == 5'b11111;
  assign _1516_ = state_in[87:80] == 5'b11110;
  assign _1517_ = state_in[87:80] == 5'b11101;
  assign _1518_ = state_in[87:80] == 5'b11100;
  assign _1519_ = state_in[87:80] == 5'b11011;
  assign _1520_ = state_in[87:80] == 5'b11010;
  assign _1521_ = state_in[87:80] == 5'b11001;
  assign _1522_ = state_in[87:80] == 5'b11000;
  assign _1523_ = state_in[87:80] == 5'b10111;
  assign _1524_ = state_in[87:80] == 5'b10110;
  assign _1525_ = state_in[87:80] == 5'b10101;
  assign _1526_ = state_in[87:80] == 5'b10100;
  assign _1527_ = state_in[87:80] == 5'b10011;
  assign _1528_ = state_in[87:80] == 5'b10010;
  assign _1529_ = state_in[87:80] == 5'b10001;
  assign _1530_ = state_in[87:80] == 5'b10000;
  assign _1531_ = state_in[87:80] == 4'b1111;
  assign _1532_ = state_in[87:80] == 4'b1110;
  assign _1533_ = state_in[87:80] == 4'b1101;
  assign _1534_ = state_in[87:80] == 4'b1100;
  assign _1535_ = state_in[87:80] == 4'b1011;
  assign _1536_ = state_in[87:80] == 4'b1010;
  assign _1537_ = state_in[87:80] == 4'b1001;
  assign _1538_ = state_in[87:80] == 4'b1000;
  assign _1539_ = state_in[87:80] == 3'b111;
  assign _1540_ = state_in[87:80] == 3'b110;
  assign _1541_ = state_in[87:80] == 3'b101;
  assign _1542_ = state_in[87:80] == 3'b100;
  assign _1543_ = state_in[87:80] == 2'b11;
  assign _1544_ = state_in[87:80] == 2'b10;
  assign _1545_ = state_in[87:80] == 1'b1;
  assign _1546_ = ! state_in[87:80];
  always @(posedge clk)
      \t1.t1.s4.out <= _1547_;
  wire [255:0] fangyuan12;
  assign fangyuan12 = { _1546_, _1545_, _1544_, _1543_, _1542_, _1541_, _1540_, _1539_, _1538_, _1537_, _1536_, _1535_, _1534_, _1533_, _1532_, _1531_, _1530_, _1529_, _1528_, _1527_, _1526_, _1525_, _1524_, _1523_, _1522_, _1521_, _1520_, _1519_, _1518_, _1517_, _1516_, _1515_, _1514_, _1513_, _1512_, _1511_, _1510_, _1509_, _1508_, _1507_, _1506_, _1505_, _1504_, _1503_, _1502_, _1501_, _1500_, _1499_, _1498_, _1497_, _1496_, _1495_, _1494_, _1493_, _1492_, _1491_, _1490_, _1489_, _1488_, _1487_, _1486_, _1485_, _1484_, _1483_, _1482_, _1481_, _1480_, _1479_, _1478_, _1477_, _1476_, _1475_, _1474_, _1473_, _1472_, _1471_, _1470_, _1469_, _1468_, _1467_, _1466_, _1465_, _1464_, _1463_, _1462_, _1461_, _1460_, _1459_, _1458_, _1457_, _1456_, _1455_, _1454_, _1453_, _1452_, _1451_, _1450_, _1449_, _1448_, _1447_, _1446_, _1445_, _1444_, _1443_, _1442_, _1441_, _1440_, _1439_, _1438_, _1437_, _1436_, _1435_, _1434_, _1433_, _1432_, _1431_, _1430_, _1429_, _1428_, _1427_, _1426_, _1425_, _1424_, _1423_, _1422_, _1421_, _1420_, _1419_, _1418_, _1417_, _1416_, _1415_, _1414_, _1413_, _1412_, _1411_, _1410_, _1409_, _1408_, _1407_, _1406_, _1405_, _1404_, _1403_, _1402_, _1401_, _1400_, _1399_, _1398_, _1397_, _1396_, _1395_, _1394_, _1393_, _1392_, _1391_, _1390_, _1389_, _1388_, _1387_, _1386_, _1385_, _1384_, _1383_, _1382_, _1381_, _1380_, _1379_, _1378_, _1377_, _1376_, _1375_, _1374_, _1373_, _1372_, _1371_, _1370_, _1369_, _1368_, _1367_, _1366_, _1365_, _1364_, _1363_, _1362_, _1361_, _1360_, _1359_, _1358_, _1357_, _1356_, _1355_, _1354_, _1353_, _1352_, _1351_, _1350_, _1349_, _1348_, _1347_, _1346_, _1345_, _1344_, _1343_, _1342_, _1341_, _1340_, _1339_, _1338_, _1337_, _1336_, _1335_, _1334_, _1333_, _1332_, _1331_, _1330_, _1329_, _1328_, _1327_, _1326_, _1325_, _1324_, _1323_, _1322_, _1321_, _1320_, _1319_, _1318_, _1317_, _1316_, _1315_, _1314_, _1313_, _1312_, _1311_, _1310_, _1309_, _1308_, _1307_, _1306_, _1305_, _1304_, _1303_, _1302_, _1301_, _1300_, _1299_, _1298_, _1297_, _1296_, _1295_, _1294_, _1293_, _1292_, _1291_ };

  always @(\t1.t1.s4.out or fangyuan12) begin
    casez (fangyuan12)
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1 :
        _1547_ = 8'b00101100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1? :
        _1547_ = 8'b01101101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?? :
        _1547_ = 8'b10101000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??? :
        _1547_ = 8'b01111011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???? :
        _1547_ = 8'b00011110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????? :
        _1547_ = 8'b01011010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????? :
        _1547_ = 8'b00101001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????? :
        _1547_ = 8'b10000010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????? :
        _1547_ = 8'b11010000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????? :
        _1547_ = 8'b10000100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????? :
        _1547_ = 8'b11010111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????? :
        _1547_ = 8'b01100101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????? :
        _1547_ = 8'b00011010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????? :
        _1547_ = 8'b00001001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????? :
        _1547_ = 8'b01011001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????? :
        _1547_ = 8'b00000011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????? :
        _1547_ = 8'b10100101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????? :
        _1547_ = 8'b01010000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????? :
        _1547_ = 8'b10101010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????? :
        _1547_ = 8'b10000111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????? :
        _1547_ = 8'b11001001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????? :
        _1547_ = 8'b00010101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????? :
        _1547_ = 8'b00111100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????? :
        _1547_ = 8'b00101101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????? :
        _1547_ = 8'b00110011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????? :
        _1547_ = 8'b00000111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????? :
        _1547_ = 8'b10101001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????? :
        _1547_ = 8'b11010010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????? :
        _1547_ = 8'b00100010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????? :
        _1547_ = 8'b00101011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????? :
        _1547_ = 8'b11101011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????? :
        _1547_ = 8'b11011001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????? :
        _1547_ = 8'b00100111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????? :
        _1547_ = 8'b00111010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????? :
        _1547_ = 8'b10011001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????? :
        _1547_ = 8'b00010111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????? :
        _1547_ = 8'b01101001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????? :
        _1547_ = 8'b10101110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????? :
        _1547_ = 8'b01101010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????? :
        _1547_ = 8'b11000010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????? :
        _1547_ = 8'b00011100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????? :
        _1547_ = 8'b11110111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????? :
        _1547_ = 8'b00000110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????? :
        _1547_ = 8'b10010000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????? :
        _1547_ = 8'b11001100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????? :
        _1547_ = 8'b01110001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????? :
        _1547_ = 8'b01111100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????? :
        _1547_ = 8'b11100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????? :
        _1547_ = 8'b00001111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????? :
        _1547_ = 8'b00001101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????? :
        _1547_ = 8'b01100001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????? :
        _1547_ = 8'b10010110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????? :
        _1547_ = 8'b00111110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????? :
        _1547_ = 8'b11101000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????? :
        _1547_ = 8'b10100001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????? :
        _1547_ = 8'b11001011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????? :
        _1547_ = 8'b10010111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????? :
        _1547_ = 8'b01110011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????? :
        _1547_ = 8'b01010111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????? :
        _1547_ = 8'b00111000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????? :
        _1547_ = 8'b01011100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????? :
        _1547_ = 8'b01001010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????? :
        _1547_ = 8'b11110000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????? :
        _1547_ = 8'b01101111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????? :
        _1547_ = 8'b00010000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b01000111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b11110100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b11001010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b11001111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b11110011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b10101100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b11011000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b01001001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b10011100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b10110001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b00000001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b11011010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b01101110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b10001011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b11010101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b11110010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b11010011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b00110001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b00111001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b11000100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b01000011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b10111101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b10011111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b10111000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b01001000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b00001100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b10010010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b00010100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b01110100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b01100100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b11011011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b10101101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b00010110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b10111100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b10100111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b00101000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b01101011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b11000111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b10001100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b00001011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b00111011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b01010100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b01000100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b10100011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b10011110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b00011001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b11000000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b11100110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b00110010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b10111010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b11001000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b01111010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b11111100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b01010101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b10010011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b00101110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b10001000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b00110101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b10111110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b11000011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b00100110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b00011000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b10000001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b10111111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b11111101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b11100101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b00100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b01000010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b10101111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b01110111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b01100011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b11110001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b01110000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b00100001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b00111111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b00000101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b10000000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b01011101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b10100010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b01001011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b00100101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b01111000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b10100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b11111110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b00000100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b11101001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b10001010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b00010001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b01100110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b10011010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b10000110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b11101101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b01001111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b11000101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b10111011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b10000101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b10110000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b10011000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b10010100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b01110010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b01100111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b10001101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b11010100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b10110110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b01111001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b11100011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b01000000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b11000001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b00000000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b10111001 ;
      256'b????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b10100110 ;
      256'b???????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b00010011 ;
      256'b??????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b01011110 ;
      256'b?????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b11011101 ;
      256'b????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b01010010 ;
      256'b???????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b01111101 ;
      256'b??????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b10110111 ;
      256'b?????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b01110110 ;
      256'b????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b10100100 ;
      256'b???????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b01011011 ;
      256'b??????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b10110100 ;
      256'b?????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b11011100 ;
      256'b????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b00110110 ;
      256'b???????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b00110100 ;
      256'b??????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b01011000 ;
      256'b?????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b00011101 ;
      256'b????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b00010010 ;
      256'b???????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b11101010 ;
      256'b??????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b01111111 ;
      256'b?????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b01001110 ;
      256'b????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b11001101 ;
      256'b???????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b11011111 ;
      256'b??????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b00011011 ;
      256'b?????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b00100100 ;
      256'b????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b00001110 ;
      256'b???????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b00101111 ;
      256'b??????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b00001010 ;
      256'b?????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b00110111 ;
      256'b????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b00110000 ;
      256'b???????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b10011101 ;
      256'b??????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b01000110 ;
      256'b?????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b10010101 ;
      256'b????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b00001000 ;
      256'b???????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b00101010 ;
      256'b??????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b01100010 ;
      256'b?????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b10101011 ;
      256'b????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b11100010 ;
      256'b???????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b11111001 ;
      256'b??????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b11010001 ;
      256'b?????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b01010001 ;
      256'b????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b01101000 ;
      256'b???????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b10000011 ;
      256'b??????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b11110101 ;
      256'b?????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b01111110 ;
      256'b????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b01101100 ;
      256'b???????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b01001100 ;
      256'b??????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b00111101 ;
      256'b?????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b11100001 ;
      256'b????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b01110101 ;
      256'b???????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b10011011 ;
      256'b??????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b11100100 ;
      256'b?????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b01010011 ;
      256'b????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b00100011 ;
      256'b???????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b01000101 ;
      256'b??????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b01011111 ;
      256'b?????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b10110011 ;
      256'b????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b01000001 ;
      256'b???????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b11111011 ;
      256'b??????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b10001110 ;
      256'b?????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b10110010 ;
      256'b????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b11101111 ;
      256'b???????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b11111010 ;
      256'b??????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b10001001 ;
      256'b?????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b00011111 ;
      256'b????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b10001111 ;
      256'b???????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b11101100 ;
      256'b??????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b01001101 ;
      256'b?????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b10110101 ;
      256'b????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b11100111 ;
      256'b???????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b01010110 ;
      256'b??????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b11001110 ;
      256'b?????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b00000010 ;
      256'b????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b01100000 ;
      256'b???????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b10010001 ;
      256'b??????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b11011110 ;
      256'b?????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b11010110 ;
      256'b????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b11111111 ;
      256'b???1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b11110110 ;
      256'b??1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b11101110 ;
      256'b?1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b11111000 ;
      256'b1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b11000110 ;
      default:
        _1547_ = \t1.t1.s4.out ;
    endcase
  end
  assign p12[23:16] = \t1.t2.s0.out ^ \t1.t2.s4.out ;
  always @(posedge clk)
      \t1.t2.s0.out <= _1548_;
  wire [255:0] fangyuan13;
  assign fangyuan13 = { _1804_, _1803_, _1802_, _1801_, _1800_, _1799_, _1798_, _1797_, _1796_, _1795_, _1794_, _1793_, _1792_, _1791_, _1790_, _1789_, _1788_, _1787_, _1786_, _1785_, _1784_, _1783_, _1782_, _1781_, _1780_, _1779_, _1778_, _1777_, _1776_, _1775_, _1774_, _1773_, _1772_, _1771_, _1770_, _1769_, _1768_, _1767_, _1766_, _1765_, _1764_, _1763_, _1762_, _1761_, _1760_, _1759_, _1758_, _1757_, _1756_, _1755_, _1754_, _1753_, _1752_, _1751_, _1750_, _1749_, _1748_, _1747_, _1746_, _1745_, _1744_, _1743_, _1742_, _1741_, _1740_, _1739_, _1738_, _1737_, _1736_, _1735_, _1734_, _1733_, _1732_, _1731_, _1730_, _1729_, _1728_, _1727_, _1726_, _1725_, _1724_, _1723_, _1722_, _1721_, _1720_, _1719_, _1718_, _1717_, _1716_, _1715_, _1714_, _1713_, _1712_, _1711_, _1710_, _1709_, _1708_, _1707_, _1706_, _1705_, _1704_, _1703_, _1702_, _1701_, _1700_, _1699_, _1698_, _1697_, _1696_, _1695_, _1694_, _1693_, _1692_, _1691_, _1690_, _1689_, _1688_, _1687_, _1686_, _1685_, _1684_, _1683_, _1682_, _1681_, _1680_, _1679_, _1678_, _1677_, _1676_, _1675_, _1674_, _1673_, _1672_, _1671_, _1670_, _1669_, _1668_, _1667_, _1666_, _1665_, _1664_, _1663_, _1662_, _1661_, _1660_, _1659_, _1658_, _1657_, _1656_, _1655_, _1654_, _1653_, _1652_, _1651_, _1650_, _1649_, _1648_, _1647_, _1646_, _1645_, _1644_, _1643_, _1642_, _1641_, _1640_, _1639_, _1638_, _1637_, _1636_, _1635_, _1634_, _1633_, _1632_, _1631_, _1630_, _1629_, _1628_, _1627_, _1626_, _1625_, _1624_, _1623_, _1622_, _1621_, _1620_, _1619_, _1618_, _1617_, _1616_, _1615_, _1614_, _1613_, _1612_, _1611_, _1610_, _1609_, _1608_, _1607_, _1606_, _1605_, _1604_, _1603_, _1602_, _1601_, _1600_, _1599_, _1598_, _1597_, _1596_, _1595_, _1594_, _1593_, _1592_, _1591_, _1590_, _1589_, _1588_, _1587_, _1586_, _1585_, _1584_, _1583_, _1582_, _1581_, _1580_, _1579_, _1578_, _1577_, _1576_, _1575_, _1574_, _1573_, _1572_, _1571_, _1570_, _1569_, _1568_, _1567_, _1566_, _1565_, _1564_, _1563_, _1562_, _1561_, _1560_, _1559_, _1558_, _1557_, _1556_, _1555_, _1554_, _1553_, _1552_, _1551_, _1550_, _1549_ };

  always @(\t1.t2.s0.out or fangyuan13) begin
    casez (fangyuan13)
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1 :
        _1548_ = 8'b00010110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1? :
        _1548_ = 8'b10111011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?? :
        _1548_ = 8'b01010100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??? :
        _1548_ = 8'b10110000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???? :
        _1548_ = 8'b00001111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????? :
        _1548_ = 8'b00101101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????? :
        _1548_ = 8'b10011001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????? :
        _1548_ = 8'b01000001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????? :
        _1548_ = 8'b01101000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????? :
        _1548_ = 8'b01000010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????? :
        _1548_ = 8'b11100110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????? :
        _1548_ = 8'b10111111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????? :
        _1548_ = 8'b00001101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????? :
        _1548_ = 8'b10001001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????? :
        _1548_ = 8'b10100001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????? :
        _1548_ = 8'b10001100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????? :
        _1548_ = 8'b11011111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????? :
        _1548_ = 8'b00101000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????? :
        _1548_ = 8'b01010101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????? :
        _1548_ = 8'b11001110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????? :
        _1548_ = 8'b11101001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????? :
        _1548_ = 8'b10000111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????? :
        _1548_ = 8'b00011110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????? :
        _1548_ = 8'b10011011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????? :
        _1548_ = 8'b10010100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????? :
        _1548_ = 8'b10001110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????? :
        _1548_ = 8'b11011001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????? :
        _1548_ = 8'b01101001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????? :
        _1548_ = 8'b00010001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????? :
        _1548_ = 8'b10011000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????? :
        _1548_ = 8'b11111000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????? :
        _1548_ = 8'b11100001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????? :
        _1548_ = 8'b10011110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????? :
        _1548_ = 8'b00011101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????? :
        _1548_ = 8'b11000001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????? :
        _1548_ = 8'b10000110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????? :
        _1548_ = 8'b10111001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????? :
        _1548_ = 8'b01010111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????? :
        _1548_ = 8'b00110101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????? :
        _1548_ = 8'b01100001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????? :
        _1548_ = 8'b00001110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????? :
        _1548_ = 8'b11110110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????? :
        _1548_ = 8'b00000011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????? :
        _1548_ = 8'b01001000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????? :
        _1548_ = 8'b01100110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????? :
        _1548_ = 8'b10110101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????? :
        _1548_ = 8'b00111110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????? :
        _1548_ = 8'b01110000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????? :
        _1548_ = 8'b10001010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????? :
        _1548_ = 8'b10001011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????? :
        _1548_ = 8'b10111101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????? :
        _1548_ = 8'b01001011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????? :
        _1548_ = 8'b00011111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????? :
        _1548_ = 8'b01110100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????? :
        _1548_ = 8'b11011101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????? :
        _1548_ = 8'b11101000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????? :
        _1548_ = 8'b11000110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????? :
        _1548_ = 8'b10110100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????? :
        _1548_ = 8'b10100110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????? :
        _1548_ = 8'b00011100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????? :
        _1548_ = 8'b00101110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????? :
        _1548_ = 8'b00100101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????? :
        _1548_ = 8'b01111000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????? :
        _1548_ = 8'b10111010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????? :
        _1548_ = 8'b00001000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b10101110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b01111010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b01100101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b11101010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b11110100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b01010110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b01101100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b10101001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b01001110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b11010101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b10001101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b01101101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b00110111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b11001000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b11100111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b01111001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b11100100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b10010101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b10010001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b01100010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b10101100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b11010011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b11000010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b01011100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b00100100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b00000110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b01001001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b00001010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b00111010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b00110010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b11100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b11011011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b00001011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b01011110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b11011110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b00010100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b10111000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b11101110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b01000110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b10001000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b10010000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b00101010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b00100010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b11011100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b01001111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b10000001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b01100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b01110011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b00011001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b01011101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b01100100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b00111101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b01111110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b10100111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b11000100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b00010111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b01000100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b10010111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b01011111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b11101100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b00010011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b00001100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b11001101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b11010010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b11110011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b11111111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b00010000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b00100001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b11011010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b10110110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b10111100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b11110101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b00111000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b10011101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b10010010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b10001111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b01000000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b10100011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b01010001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b10101000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b10011111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b00111100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b01010000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b01111111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b00000010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b11111001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b01000101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b10000101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b00110011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b01001101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b01000011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b11111011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b10101010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b11101111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b11010000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b11001111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b01011000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b01001100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b01001010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b00111001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b10111110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b11001011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b01101010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b01011011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b10110001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b11111100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b00100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b11101101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b00000000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b11010001 ;
      256'b????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b01010011 ;
      256'b???????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b10000100 ;
      256'b??????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b00101111 ;
      256'b?????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b11100011 ;
      256'b????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b00101001 ;
      256'b???????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b10110011 ;
      256'b??????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b11010110 ;
      256'b?????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b00111011 ;
      256'b????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b01010010 ;
      256'b???????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b10100000 ;
      256'b??????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b01011010 ;
      256'b?????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b01101110 ;
      256'b????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b00011011 ;
      256'b???????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b00011010 ;
      256'b??????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b00101100 ;
      256'b?????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b10000011 ;
      256'b????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b00001001 ;
      256'b???????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b01110101 ;
      256'b??????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b10110010 ;
      256'b?????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b00100111 ;
      256'b????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b11101011 ;
      256'b???????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b11100010 ;
      256'b??????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b10000000 ;
      256'b?????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b00010010 ;
      256'b????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b00000111 ;
      256'b???????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b10011010 ;
      256'b??????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b00000101 ;
      256'b?????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b10010110 ;
      256'b????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b00011000 ;
      256'b???????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b11000011 ;
      256'b??????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b00100011 ;
      256'b?????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b11000111 ;
      256'b????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b00000100 ;
      256'b???????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b00010101 ;
      256'b??????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b00110001 ;
      256'b?????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b11011000 ;
      256'b????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b01110001 ;
      256'b???????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b11110001 ;
      256'b??????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b11100101 ;
      256'b?????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b10100101 ;
      256'b????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b00110100 ;
      256'b???????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b11001100 ;
      256'b??????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b11110111 ;
      256'b?????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b00111111 ;
      256'b????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b00110110 ;
      256'b???????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b00100110 ;
      256'b??????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b10010011 ;
      256'b?????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b11111101 ;
      256'b????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b10110111 ;
      256'b???????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b11000000 ;
      256'b??????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b01110010 ;
      256'b?????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b10100100 ;
      256'b????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b10011100 ;
      256'b???????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b10101111 ;
      256'b??????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b10100010 ;
      256'b?????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b11010100 ;
      256'b????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b10101101 ;
      256'b???????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b11110000 ;
      256'b??????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b01000111 ;
      256'b?????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b01011001 ;
      256'b????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b11111010 ;
      256'b???????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b01111101 ;
      256'b??????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b11001001 ;
      256'b?????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b10000010 ;
      256'b????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b11001010 ;
      256'b???????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b01110110 ;
      256'b??????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b10101011 ;
      256'b?????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b11010111 ;
      256'b????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b11111110 ;
      256'b???????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b00101011 ;
      256'b??????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b01100111 ;
      256'b?????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b00000001 ;
      256'b????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b00110000 ;
      256'b???????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b11000101 ;
      256'b??????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b01101111 ;
      256'b?????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b01101011 ;
      256'b????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b11110010 ;
      256'b???1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b01111011 ;
      256'b??1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b01110111 ;
      256'b?1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b01111100 ;
      256'b1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b01100011 ;
      default:
        _1548_ = \t1.t2.s0.out ;
    endcase
  end
  assign _1549_ = state_in[79:72] == 8'b11111111;
  assign _1550_ = state_in[79:72] == 8'b11111110;
  assign _1551_ = state_in[79:72] == 8'b11111101;
  assign _1552_ = state_in[79:72] == 8'b11111100;
  assign _1553_ = state_in[79:72] == 8'b11111011;
  assign _1554_ = state_in[79:72] == 8'b11111010;
  assign _1555_ = state_in[79:72] == 8'b11111001;
  assign _1556_ = state_in[79:72] == 8'b11111000;
  assign _1557_ = state_in[79:72] == 8'b11110111;
  assign _1558_ = state_in[79:72] == 8'b11110110;
  assign _1559_ = state_in[79:72] == 8'b11110101;
  assign _1560_ = state_in[79:72] == 8'b11110100;
  assign _1561_ = state_in[79:72] == 8'b11110011;
  assign _1562_ = state_in[79:72] == 8'b11110010;
  assign _1563_ = state_in[79:72] == 8'b11110001;
  assign _1564_ = state_in[79:72] == 8'b11110000;
  assign _1565_ = state_in[79:72] == 8'b11101111;
  assign _1566_ = state_in[79:72] == 8'b11101110;
  assign _1567_ = state_in[79:72] == 8'b11101101;
  assign _1568_ = state_in[79:72] == 8'b11101100;
  assign _1569_ = state_in[79:72] == 8'b11101011;
  assign _1570_ = state_in[79:72] == 8'b11101010;
  assign _1571_ = state_in[79:72] == 8'b11101001;
  assign _1572_ = state_in[79:72] == 8'b11101000;
  assign _1573_ = state_in[79:72] == 8'b11100111;
  assign _1574_ = state_in[79:72] == 8'b11100110;
  assign _1575_ = state_in[79:72] == 8'b11100101;
  assign _1576_ = state_in[79:72] == 8'b11100100;
  assign _1577_ = state_in[79:72] == 8'b11100011;
  assign _1578_ = state_in[79:72] == 8'b11100010;
  assign _1579_ = state_in[79:72] == 8'b11100001;
  assign _1580_ = state_in[79:72] == 8'b11100000;
  assign _1581_ = state_in[79:72] == 8'b11011111;
  assign _1582_ = state_in[79:72] == 8'b11011110;
  assign _1583_ = state_in[79:72] == 8'b11011101;
  assign _1584_ = state_in[79:72] == 8'b11011100;
  assign _1585_ = state_in[79:72] == 8'b11011011;
  assign _1586_ = state_in[79:72] == 8'b11011010;
  assign _1587_ = state_in[79:72] == 8'b11011001;
  assign _1588_ = state_in[79:72] == 8'b11011000;
  assign _1589_ = state_in[79:72] == 8'b11010111;
  assign _1590_ = state_in[79:72] == 8'b11010110;
  assign _1591_ = state_in[79:72] == 8'b11010101;
  assign _1592_ = state_in[79:72] == 8'b11010100;
  assign _1593_ = state_in[79:72] == 8'b11010011;
  assign _1594_ = state_in[79:72] == 8'b11010010;
  assign _1595_ = state_in[79:72] == 8'b11010001;
  assign _1596_ = state_in[79:72] == 8'b11010000;
  assign _1597_ = state_in[79:72] == 8'b11001111;
  assign _1598_ = state_in[79:72] == 8'b11001110;
  assign _1599_ = state_in[79:72] == 8'b11001101;
  assign _1600_ = state_in[79:72] == 8'b11001100;
  assign _1601_ = state_in[79:72] == 8'b11001011;
  assign _1602_ = state_in[79:72] == 8'b11001010;
  assign _1603_ = state_in[79:72] == 8'b11001001;
  assign _1604_ = state_in[79:72] == 8'b11001000;
  assign _1605_ = state_in[79:72] == 8'b11000111;
  assign _1606_ = state_in[79:72] == 8'b11000110;
  assign _1607_ = state_in[79:72] == 8'b11000101;
  assign _1608_ = state_in[79:72] == 8'b11000100;
  assign _1609_ = state_in[79:72] == 8'b11000011;
  assign _1610_ = state_in[79:72] == 8'b11000010;
  assign _1611_ = state_in[79:72] == 8'b11000001;
  assign _1612_ = state_in[79:72] == 8'b11000000;
  assign _1613_ = state_in[79:72] == 8'b10111111;
  assign _1614_ = state_in[79:72] == 8'b10111110;
  assign _1615_ = state_in[79:72] == 8'b10111101;
  assign _1616_ = state_in[79:72] == 8'b10111100;
  assign _1617_ = state_in[79:72] == 8'b10111011;
  assign _1618_ = state_in[79:72] == 8'b10111010;
  assign _1619_ = state_in[79:72] == 8'b10111001;
  assign _1620_ = state_in[79:72] == 8'b10111000;
  assign _1621_ = state_in[79:72] == 8'b10110111;
  assign _1622_ = state_in[79:72] == 8'b10110110;
  assign _1623_ = state_in[79:72] == 8'b10110101;
  assign _1624_ = state_in[79:72] == 8'b10110100;
  assign _1625_ = state_in[79:72] == 8'b10110011;
  assign _1626_ = state_in[79:72] == 8'b10110010;
  assign _1627_ = state_in[79:72] == 8'b10110001;
  assign _1628_ = state_in[79:72] == 8'b10110000;
  assign _1629_ = state_in[79:72] == 8'b10101111;
  assign _1630_ = state_in[79:72] == 8'b10101110;
  assign _1631_ = state_in[79:72] == 8'b10101101;
  assign _1632_ = state_in[79:72] == 8'b10101100;
  assign _1633_ = state_in[79:72] == 8'b10101011;
  assign _1634_ = state_in[79:72] == 8'b10101010;
  assign _1635_ = state_in[79:72] == 8'b10101001;
  assign _1636_ = state_in[79:72] == 8'b10101000;
  assign _1637_ = state_in[79:72] == 8'b10100111;
  assign _1638_ = state_in[79:72] == 8'b10100110;
  assign _1639_ = state_in[79:72] == 8'b10100101;
  assign _1640_ = state_in[79:72] == 8'b10100100;
  assign _1641_ = state_in[79:72] == 8'b10100011;
  assign _1642_ = state_in[79:72] == 8'b10100010;
  assign _1643_ = state_in[79:72] == 8'b10100001;
  assign _1644_ = state_in[79:72] == 8'b10100000;
  assign _1645_ = state_in[79:72] == 8'b10011111;
  assign _1646_ = state_in[79:72] == 8'b10011110;
  assign _1647_ = state_in[79:72] == 8'b10011101;
  assign _1648_ = state_in[79:72] == 8'b10011100;
  assign _1649_ = state_in[79:72] == 8'b10011011;
  assign _1650_ = state_in[79:72] == 8'b10011010;
  assign _1651_ = state_in[79:72] == 8'b10011001;
  assign _1652_ = state_in[79:72] == 8'b10011000;
  assign _1653_ = state_in[79:72] == 8'b10010111;
  assign _1654_ = state_in[79:72] == 8'b10010110;
  assign _1655_ = state_in[79:72] == 8'b10010101;
  assign _1656_ = state_in[79:72] == 8'b10010100;
  assign _1657_ = state_in[79:72] == 8'b10010011;
  assign _1658_ = state_in[79:72] == 8'b10010010;
  assign _1659_ = state_in[79:72] == 8'b10010001;
  assign _1660_ = state_in[79:72] == 8'b10010000;
  assign _1661_ = state_in[79:72] == 8'b10001111;
  assign _1662_ = state_in[79:72] == 8'b10001110;
  assign _1663_ = state_in[79:72] == 8'b10001101;
  assign _1664_ = state_in[79:72] == 8'b10001100;
  assign _1665_ = state_in[79:72] == 8'b10001011;
  assign _1666_ = state_in[79:72] == 8'b10001010;
  assign _1667_ = state_in[79:72] == 8'b10001001;
  assign _1668_ = state_in[79:72] == 8'b10001000;
  assign _1669_ = state_in[79:72] == 8'b10000111;
  assign _1670_ = state_in[79:72] == 8'b10000110;
  assign _1671_ = state_in[79:72] == 8'b10000101;
  assign _1672_ = state_in[79:72] == 8'b10000100;
  assign _1673_ = state_in[79:72] == 8'b10000011;
  assign _1674_ = state_in[79:72] == 8'b10000010;
  assign _1675_ = state_in[79:72] == 8'b10000001;
  assign _1676_ = state_in[79:72] == 8'b10000000;
  assign _1677_ = state_in[79:72] == 7'b1111111;
  assign _1678_ = state_in[79:72] == 7'b1111110;
  assign _1679_ = state_in[79:72] == 7'b1111101;
  assign _1680_ = state_in[79:72] == 7'b1111100;
  assign _1681_ = state_in[79:72] == 7'b1111011;
  assign _1682_ = state_in[79:72] == 7'b1111010;
  assign _1683_ = state_in[79:72] == 7'b1111001;
  assign _1684_ = state_in[79:72] == 7'b1111000;
  assign _1685_ = state_in[79:72] == 7'b1110111;
  assign _1686_ = state_in[79:72] == 7'b1110110;
  assign _1687_ = state_in[79:72] == 7'b1110101;
  assign _1688_ = state_in[79:72] == 7'b1110100;
  assign _1689_ = state_in[79:72] == 7'b1110011;
  assign _1690_ = state_in[79:72] == 7'b1110010;
  assign _1691_ = state_in[79:72] == 7'b1110001;
  assign _1692_ = state_in[79:72] == 7'b1110000;
  assign _1693_ = state_in[79:72] == 7'b1101111;
  assign _1694_ = state_in[79:72] == 7'b1101110;
  assign _1695_ = state_in[79:72] == 7'b1101101;
  assign _1696_ = state_in[79:72] == 7'b1101100;
  assign _1697_ = state_in[79:72] == 7'b1101011;
  assign _1698_ = state_in[79:72] == 7'b1101010;
  assign _1699_ = state_in[79:72] == 7'b1101001;
  assign _1700_ = state_in[79:72] == 7'b1101000;
  assign _1701_ = state_in[79:72] == 7'b1100111;
  assign _1702_ = state_in[79:72] == 7'b1100110;
  assign _1703_ = state_in[79:72] == 7'b1100101;
  assign _1704_ = state_in[79:72] == 7'b1100100;
  assign _1705_ = state_in[79:72] == 7'b1100011;
  assign _1706_ = state_in[79:72] == 7'b1100010;
  assign _1707_ = state_in[79:72] == 7'b1100001;
  assign _1708_ = state_in[79:72] == 7'b1100000;
  assign _1709_ = state_in[79:72] == 7'b1011111;
  assign _1710_ = state_in[79:72] == 7'b1011110;
  assign _1711_ = state_in[79:72] == 7'b1011101;
  assign _1712_ = state_in[79:72] == 7'b1011100;
  assign _1713_ = state_in[79:72] == 7'b1011011;
  assign _1714_ = state_in[79:72] == 7'b1011010;
  assign _1715_ = state_in[79:72] == 7'b1011001;
  assign _1716_ = state_in[79:72] == 7'b1011000;
  assign _1717_ = state_in[79:72] == 7'b1010111;
  assign _1718_ = state_in[79:72] == 7'b1010110;
  assign _1719_ = state_in[79:72] == 7'b1010101;
  assign _1720_ = state_in[79:72] == 7'b1010100;
  assign _1721_ = state_in[79:72] == 7'b1010011;
  assign _1722_ = state_in[79:72] == 7'b1010010;
  assign _1723_ = state_in[79:72] == 7'b1010001;
  assign _1724_ = state_in[79:72] == 7'b1010000;
  assign _1725_ = state_in[79:72] == 7'b1001111;
  assign _1726_ = state_in[79:72] == 7'b1001110;
  assign _1727_ = state_in[79:72] == 7'b1001101;
  assign _1728_ = state_in[79:72] == 7'b1001100;
  assign _1729_ = state_in[79:72] == 7'b1001011;
  assign _1730_ = state_in[79:72] == 7'b1001010;
  assign _1731_ = state_in[79:72] == 7'b1001001;
  assign _1732_ = state_in[79:72] == 7'b1001000;
  assign _1733_ = state_in[79:72] == 7'b1000111;
  assign _1734_ = state_in[79:72] == 7'b1000110;
  assign _1735_ = state_in[79:72] == 7'b1000101;
  assign _1736_ = state_in[79:72] == 7'b1000100;
  assign _1737_ = state_in[79:72] == 7'b1000011;
  assign _1738_ = state_in[79:72] == 7'b1000010;
  assign _1739_ = state_in[79:72] == 7'b1000001;
  assign _1740_ = state_in[79:72] == 7'b1000000;
  assign _1741_ = state_in[79:72] == 6'b111111;
  assign _1742_ = state_in[79:72] == 6'b111110;
  assign _1743_ = state_in[79:72] == 6'b111101;
  assign _1744_ = state_in[79:72] == 6'b111100;
  assign _1745_ = state_in[79:72] == 6'b111011;
  assign _1746_ = state_in[79:72] == 6'b111010;
  assign _1747_ = state_in[79:72] == 6'b111001;
  assign _1748_ = state_in[79:72] == 6'b111000;
  assign _1749_ = state_in[79:72] == 6'b110111;
  assign _1750_ = state_in[79:72] == 6'b110110;
  assign _1751_ = state_in[79:72] == 6'b110101;
  assign _1752_ = state_in[79:72] == 6'b110100;
  assign _1753_ = state_in[79:72] == 6'b110011;
  assign _1754_ = state_in[79:72] == 6'b110010;
  assign _1755_ = state_in[79:72] == 6'b110001;
  assign _1756_ = state_in[79:72] == 6'b110000;
  assign _1757_ = state_in[79:72] == 6'b101111;
  assign _1758_ = state_in[79:72] == 6'b101110;
  assign _1759_ = state_in[79:72] == 6'b101101;
  assign _1760_ = state_in[79:72] == 6'b101100;
  assign _1761_ = state_in[79:72] == 6'b101011;
  assign _1762_ = state_in[79:72] == 6'b101010;
  assign _1763_ = state_in[79:72] == 6'b101001;
  assign _1764_ = state_in[79:72] == 6'b101000;
  assign _1765_ = state_in[79:72] == 6'b100111;
  assign _1766_ = state_in[79:72] == 6'b100110;
  assign _1767_ = state_in[79:72] == 6'b100101;
  assign _1768_ = state_in[79:72] == 6'b100100;
  assign _1769_ = state_in[79:72] == 6'b100011;
  assign _1770_ = state_in[79:72] == 6'b100010;
  assign _1771_ = state_in[79:72] == 6'b100001;
  assign _1772_ = state_in[79:72] == 6'b100000;
  assign _1773_ = state_in[79:72] == 5'b11111;
  assign _1774_ = state_in[79:72] == 5'b11110;
  assign _1775_ = state_in[79:72] == 5'b11101;
  assign _1776_ = state_in[79:72] == 5'b11100;
  assign _1777_ = state_in[79:72] == 5'b11011;
  assign _1778_ = state_in[79:72] == 5'b11010;
  assign _1779_ = state_in[79:72] == 5'b11001;
  assign _1780_ = state_in[79:72] == 5'b11000;
  assign _1781_ = state_in[79:72] == 5'b10111;
  assign _1782_ = state_in[79:72] == 5'b10110;
  assign _1783_ = state_in[79:72] == 5'b10101;
  assign _1784_ = state_in[79:72] == 5'b10100;
  assign _1785_ = state_in[79:72] == 5'b10011;
  assign _1786_ = state_in[79:72] == 5'b10010;
  assign _1787_ = state_in[79:72] == 5'b10001;
  assign _1788_ = state_in[79:72] == 5'b10000;
  assign _1789_ = state_in[79:72] == 4'b1111;
  assign _1790_ = state_in[79:72] == 4'b1110;
  assign _1791_ = state_in[79:72] == 4'b1101;
  assign _1792_ = state_in[79:72] == 4'b1100;
  assign _1793_ = state_in[79:72] == 4'b1011;
  assign _1794_ = state_in[79:72] == 4'b1010;
  assign _1795_ = state_in[79:72] == 4'b1001;
  assign _1796_ = state_in[79:72] == 4'b1000;
  assign _1797_ = state_in[79:72] == 3'b111;
  assign _1798_ = state_in[79:72] == 3'b110;
  assign _1799_ = state_in[79:72] == 3'b101;
  assign _1800_ = state_in[79:72] == 3'b100;
  assign _1801_ = state_in[79:72] == 2'b11;
  assign _1802_ = state_in[79:72] == 2'b10;
  assign _1803_ = state_in[79:72] == 1'b1;
  assign _1804_ = ! state_in[79:72];
  always @(posedge clk)
      \t1.t2.s4.out <= _1805_;
  wire [255:0] fangyuan14;
  assign fangyuan14 = { _1804_, _1803_, _1802_, _1801_, _1800_, _1799_, _1798_, _1797_, _1796_, _1795_, _1794_, _1793_, _1792_, _1791_, _1790_, _1789_, _1788_, _1787_, _1786_, _1785_, _1784_, _1783_, _1782_, _1781_, _1780_, _1779_, _1778_, _1777_, _1776_, _1775_, _1774_, _1773_, _1772_, _1771_, _1770_, _1769_, _1768_, _1767_, _1766_, _1765_, _1764_, _1763_, _1762_, _1761_, _1760_, _1759_, _1758_, _1757_, _1756_, _1755_, _1754_, _1753_, _1752_, _1751_, _1750_, _1749_, _1748_, _1747_, _1746_, _1745_, _1744_, _1743_, _1742_, _1741_, _1740_, _1739_, _1738_, _1737_, _1736_, _1735_, _1734_, _1733_, _1732_, _1731_, _1730_, _1729_, _1728_, _1727_, _1726_, _1725_, _1724_, _1723_, _1722_, _1721_, _1720_, _1719_, _1718_, _1717_, _1716_, _1715_, _1714_, _1713_, _1712_, _1711_, _1710_, _1709_, _1708_, _1707_, _1706_, _1705_, _1704_, _1703_, _1702_, _1701_, _1700_, _1699_, _1698_, _1697_, _1696_, _1695_, _1694_, _1693_, _1692_, _1691_, _1690_, _1689_, _1688_, _1687_, _1686_, _1685_, _1684_, _1683_, _1682_, _1681_, _1680_, _1679_, _1678_, _1677_, _1676_, _1675_, _1674_, _1673_, _1672_, _1671_, _1670_, _1669_, _1668_, _1667_, _1666_, _1665_, _1664_, _1663_, _1662_, _1661_, _1660_, _1659_, _1658_, _1657_, _1656_, _1655_, _1654_, _1653_, _1652_, _1651_, _1650_, _1649_, _1648_, _1647_, _1646_, _1645_, _1644_, _1643_, _1642_, _1641_, _1640_, _1639_, _1638_, _1637_, _1636_, _1635_, _1634_, _1633_, _1632_, _1631_, _1630_, _1629_, _1628_, _1627_, _1626_, _1625_, _1624_, _1623_, _1622_, _1621_, _1620_, _1619_, _1618_, _1617_, _1616_, _1615_, _1614_, _1613_, _1612_, _1611_, _1610_, _1609_, _1608_, _1607_, _1606_, _1605_, _1604_, _1603_, _1602_, _1601_, _1600_, _1599_, _1598_, _1597_, _1596_, _1595_, _1594_, _1593_, _1592_, _1591_, _1590_, _1589_, _1588_, _1587_, _1586_, _1585_, _1584_, _1583_, _1582_, _1581_, _1580_, _1579_, _1578_, _1577_, _1576_, _1575_, _1574_, _1573_, _1572_, _1571_, _1570_, _1569_, _1568_, _1567_, _1566_, _1565_, _1564_, _1563_, _1562_, _1561_, _1560_, _1559_, _1558_, _1557_, _1556_, _1555_, _1554_, _1553_, _1552_, _1551_, _1550_, _1549_ };

  always @(\t1.t2.s4.out or fangyuan14) begin
    casez (fangyuan14)
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1 :
        _1805_ = 8'b00101100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1? :
        _1805_ = 8'b01101101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?? :
        _1805_ = 8'b10101000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??? :
        _1805_ = 8'b01111011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???? :
        _1805_ = 8'b00011110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????? :
        _1805_ = 8'b01011010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????? :
        _1805_ = 8'b00101001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????? :
        _1805_ = 8'b10000010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????? :
        _1805_ = 8'b11010000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????? :
        _1805_ = 8'b10000100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????? :
        _1805_ = 8'b11010111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????? :
        _1805_ = 8'b01100101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????? :
        _1805_ = 8'b00011010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????? :
        _1805_ = 8'b00001001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????? :
        _1805_ = 8'b01011001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????? :
        _1805_ = 8'b00000011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????? :
        _1805_ = 8'b10100101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????? :
        _1805_ = 8'b01010000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????? :
        _1805_ = 8'b10101010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????? :
        _1805_ = 8'b10000111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????? :
        _1805_ = 8'b11001001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????? :
        _1805_ = 8'b00010101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????? :
        _1805_ = 8'b00111100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????? :
        _1805_ = 8'b00101101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????? :
        _1805_ = 8'b00110011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????? :
        _1805_ = 8'b00000111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????? :
        _1805_ = 8'b10101001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????? :
        _1805_ = 8'b11010010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????? :
        _1805_ = 8'b00100010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????? :
        _1805_ = 8'b00101011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????? :
        _1805_ = 8'b11101011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????? :
        _1805_ = 8'b11011001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????? :
        _1805_ = 8'b00100111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????? :
        _1805_ = 8'b00111010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????? :
        _1805_ = 8'b10011001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????? :
        _1805_ = 8'b00010111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????? :
        _1805_ = 8'b01101001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????? :
        _1805_ = 8'b10101110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????? :
        _1805_ = 8'b01101010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????? :
        _1805_ = 8'b11000010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????? :
        _1805_ = 8'b00011100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????? :
        _1805_ = 8'b11110111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????? :
        _1805_ = 8'b00000110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????? :
        _1805_ = 8'b10010000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????? :
        _1805_ = 8'b11001100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????? :
        _1805_ = 8'b01110001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????? :
        _1805_ = 8'b01111100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????? :
        _1805_ = 8'b11100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????? :
        _1805_ = 8'b00001111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????? :
        _1805_ = 8'b00001101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????? :
        _1805_ = 8'b01100001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????? :
        _1805_ = 8'b10010110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????? :
        _1805_ = 8'b00111110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????? :
        _1805_ = 8'b11101000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????? :
        _1805_ = 8'b10100001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????? :
        _1805_ = 8'b11001011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????? :
        _1805_ = 8'b10010111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????? :
        _1805_ = 8'b01110011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????? :
        _1805_ = 8'b01010111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????? :
        _1805_ = 8'b00111000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????? :
        _1805_ = 8'b01011100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????? :
        _1805_ = 8'b01001010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????? :
        _1805_ = 8'b11110000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????? :
        _1805_ = 8'b01101111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????? :
        _1805_ = 8'b00010000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b01000111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b11110100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b11001010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b11001111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b11110011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b10101100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b11011000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b01001001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b10011100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b10110001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b00000001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b11011010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b01101110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b10001011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b11010101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b11110010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b11010011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b00110001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b00111001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b11000100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b01000011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b10111101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b10011111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b10111000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b01001000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b00001100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b10010010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b00010100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b01110100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b01100100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b11011011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b10101101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b00010110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b10111100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b10100111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b00101000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b01101011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b11000111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b10001100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b00001011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b00111011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b01010100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b01000100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b10100011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b10011110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b00011001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b11000000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b11100110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b00110010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b10111010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b11001000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b01111010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b11111100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b01010101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b10010011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b00101110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b10001000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b00110101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b10111110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b11000011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b00100110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b00011000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b10000001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b10111111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b11111101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b11100101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b00100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b01000010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b10101111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b01110111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b01100011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b11110001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b01110000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b00100001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b00111111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b00000101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b10000000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b01011101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b10100010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b01001011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b00100101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b01111000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b10100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b11111110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b00000100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b11101001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b10001010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b00010001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b01100110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b10011010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b10000110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b11101101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b01001111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b11000101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b10111011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b10000101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b10110000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b10011000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b10010100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b01110010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b01100111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b10001101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b11010100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b10110110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b01111001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b11100011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b01000000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b11000001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b00000000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b10111001 ;
      256'b????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b10100110 ;
      256'b???????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b00010011 ;
      256'b??????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b01011110 ;
      256'b?????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b11011101 ;
      256'b????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b01010010 ;
      256'b???????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b01111101 ;
      256'b??????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b10110111 ;
      256'b?????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b01110110 ;
      256'b????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b10100100 ;
      256'b???????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b01011011 ;
      256'b??????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b10110100 ;
      256'b?????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b11011100 ;
      256'b????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b00110110 ;
      256'b???????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b00110100 ;
      256'b??????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b01011000 ;
      256'b?????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b00011101 ;
      256'b????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b00010010 ;
      256'b???????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b11101010 ;
      256'b??????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b01111111 ;
      256'b?????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b01001110 ;
      256'b????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b11001101 ;
      256'b???????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b11011111 ;
      256'b??????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b00011011 ;
      256'b?????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b00100100 ;
      256'b????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b00001110 ;
      256'b???????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b00101111 ;
      256'b??????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b00001010 ;
      256'b?????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b00110111 ;
      256'b????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b00110000 ;
      256'b???????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b10011101 ;
      256'b??????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b01000110 ;
      256'b?????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b10010101 ;
      256'b????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b00001000 ;
      256'b???????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b00101010 ;
      256'b??????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b01100010 ;
      256'b?????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b10101011 ;
      256'b????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b11100010 ;
      256'b???????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b11111001 ;
      256'b??????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b11010001 ;
      256'b?????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b01010001 ;
      256'b????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b01101000 ;
      256'b???????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b10000011 ;
      256'b??????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b11110101 ;
      256'b?????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b01111110 ;
      256'b????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b01101100 ;
      256'b???????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b01001100 ;
      256'b??????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b00111101 ;
      256'b?????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b11100001 ;
      256'b????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b01110101 ;
      256'b???????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b10011011 ;
      256'b??????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b11100100 ;
      256'b?????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b01010011 ;
      256'b????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b00100011 ;
      256'b???????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b01000101 ;
      256'b??????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b01011111 ;
      256'b?????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b10110011 ;
      256'b????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b01000001 ;
      256'b???????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b11111011 ;
      256'b??????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b10001110 ;
      256'b?????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b10110010 ;
      256'b????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b11101111 ;
      256'b???????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b11111010 ;
      256'b??????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b10001001 ;
      256'b?????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b00011111 ;
      256'b????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b10001111 ;
      256'b???????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b11101100 ;
      256'b??????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b01001101 ;
      256'b?????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b10110101 ;
      256'b????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b11100111 ;
      256'b???????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b01010110 ;
      256'b??????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b11001110 ;
      256'b?????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b00000010 ;
      256'b????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b01100000 ;
      256'b???????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b10010001 ;
      256'b??????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b11011110 ;
      256'b?????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b11010110 ;
      256'b????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b11111111 ;
      256'b???1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b11110110 ;
      256'b??1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b11101110 ;
      256'b?1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b11111000 ;
      256'b1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b11000110 ;
      default:
        _1805_ = \t1.t2.s4.out ;
    endcase
  end
  assign p13[15:8] = \t1.t3.s0.out ^ \t1.t3.s4.out ;
  always @(posedge clk)
      \t1.t3.s0.out <= _1806_;
  wire [255:0] fangyuan15;
  assign fangyuan15 = { _2062_, _2061_, _2060_, _2059_, _2058_, _2057_, _2056_, _2055_, _2054_, _2053_, _2052_, _2051_, _2050_, _2049_, _2048_, _2047_, _2046_, _2045_, _2044_, _2043_, _2042_, _2041_, _2040_, _2039_, _2038_, _2037_, _2036_, _2035_, _2034_, _2033_, _2032_, _2031_, _2030_, _2029_, _2028_, _2027_, _2026_, _2025_, _2024_, _2023_, _2022_, _2021_, _2020_, _2019_, _2018_, _2017_, _2016_, _2015_, _2014_, _2013_, _2012_, _2011_, _2010_, _2009_, _2008_, _2007_, _2006_, _2005_, _2004_, _2003_, _2002_, _2001_, _2000_, _1999_, _1998_, _1997_, _1996_, _1995_, _1994_, _1993_, _1992_, _1991_, _1990_, _1989_, _1988_, _1987_, _1986_, _1985_, _1984_, _1983_, _1982_, _1981_, _1980_, _1979_, _1978_, _1977_, _1976_, _1975_, _1974_, _1973_, _1972_, _1971_, _1970_, _1969_, _1968_, _1967_, _1966_, _1965_, _1964_, _1963_, _1962_, _1961_, _1960_, _1959_, _1958_, _1957_, _1956_, _1955_, _1954_, _1953_, _1952_, _1951_, _1950_, _1949_, _1948_, _1947_, _1946_, _1945_, _1944_, _1943_, _1942_, _1941_, _1940_, _1939_, _1938_, _1937_, _1936_, _1935_, _1934_, _1933_, _1932_, _1931_, _1930_, _1929_, _1928_, _1927_, _1926_, _1925_, _1924_, _1923_, _1922_, _1921_, _1920_, _1919_, _1918_, _1917_, _1916_, _1915_, _1914_, _1913_, _1912_, _1911_, _1910_, _1909_, _1908_, _1907_, _1906_, _1905_, _1904_, _1903_, _1902_, _1901_, _1900_, _1899_, _1898_, _1897_, _1896_, _1895_, _1894_, _1893_, _1892_, _1891_, _1890_, _1889_, _1888_, _1887_, _1886_, _1885_, _1884_, _1883_, _1882_, _1881_, _1880_, _1879_, _1878_, _1877_, _1876_, _1875_, _1874_, _1873_, _1872_, _1871_, _1870_, _1869_, _1868_, _1867_, _1866_, _1865_, _1864_, _1863_, _1862_, _1861_, _1860_, _1859_, _1858_, _1857_, _1856_, _1855_, _1854_, _1853_, _1852_, _1851_, _1850_, _1849_, _1848_, _1847_, _1846_, _1845_, _1844_, _1843_, _1842_, _1841_, _1840_, _1839_, _1838_, _1837_, _1836_, _1835_, _1834_, _1833_, _1832_, _1831_, _1830_, _1829_, _1828_, _1827_, _1826_, _1825_, _1824_, _1823_, _1822_, _1821_, _1820_, _1819_, _1818_, _1817_, _1816_, _1815_, _1814_, _1813_, _1812_, _1811_, _1810_, _1809_, _1808_, _1807_ };

  always @(\t1.t3.s0.out or fangyuan15) begin
    casez (fangyuan15)
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1 :
        _1806_ = 8'b00010110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1? :
        _1806_ = 8'b10111011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?? :
        _1806_ = 8'b01010100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??? :
        _1806_ = 8'b10110000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???? :
        _1806_ = 8'b00001111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????? :
        _1806_ = 8'b00101101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????? :
        _1806_ = 8'b10011001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????? :
        _1806_ = 8'b01000001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????? :
        _1806_ = 8'b01101000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????? :
        _1806_ = 8'b01000010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????? :
        _1806_ = 8'b11100110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????? :
        _1806_ = 8'b10111111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????? :
        _1806_ = 8'b00001101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????? :
        _1806_ = 8'b10001001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????? :
        _1806_ = 8'b10100001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????? :
        _1806_ = 8'b10001100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????? :
        _1806_ = 8'b11011111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????? :
        _1806_ = 8'b00101000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????? :
        _1806_ = 8'b01010101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????? :
        _1806_ = 8'b11001110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????? :
        _1806_ = 8'b11101001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????? :
        _1806_ = 8'b10000111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????? :
        _1806_ = 8'b00011110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????? :
        _1806_ = 8'b10011011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????? :
        _1806_ = 8'b10010100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????? :
        _1806_ = 8'b10001110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????? :
        _1806_ = 8'b11011001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????? :
        _1806_ = 8'b01101001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????? :
        _1806_ = 8'b00010001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????? :
        _1806_ = 8'b10011000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????? :
        _1806_ = 8'b11111000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????? :
        _1806_ = 8'b11100001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????? :
        _1806_ = 8'b10011110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????? :
        _1806_ = 8'b00011101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????? :
        _1806_ = 8'b11000001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????? :
        _1806_ = 8'b10000110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????? :
        _1806_ = 8'b10111001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????? :
        _1806_ = 8'b01010111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????? :
        _1806_ = 8'b00110101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????? :
        _1806_ = 8'b01100001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????? :
        _1806_ = 8'b00001110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????? :
        _1806_ = 8'b11110110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????? :
        _1806_ = 8'b00000011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????? :
        _1806_ = 8'b01001000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????? :
        _1806_ = 8'b01100110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????? :
        _1806_ = 8'b10110101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????? :
        _1806_ = 8'b00111110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????? :
        _1806_ = 8'b01110000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????? :
        _1806_ = 8'b10001010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????? :
        _1806_ = 8'b10001011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????? :
        _1806_ = 8'b10111101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????? :
        _1806_ = 8'b01001011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????? :
        _1806_ = 8'b00011111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????? :
        _1806_ = 8'b01110100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????? :
        _1806_ = 8'b11011101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????? :
        _1806_ = 8'b11101000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????? :
        _1806_ = 8'b11000110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????? :
        _1806_ = 8'b10110100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????? :
        _1806_ = 8'b10100110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????? :
        _1806_ = 8'b00011100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????? :
        _1806_ = 8'b00101110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????? :
        _1806_ = 8'b00100101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????? :
        _1806_ = 8'b01111000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????? :
        _1806_ = 8'b10111010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????? :
        _1806_ = 8'b00001000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b10101110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b01111010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b01100101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b11101010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b11110100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b01010110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b01101100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b10101001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b01001110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b11010101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b10001101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b01101101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b00110111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b11001000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b11100111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b01111001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b11100100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b10010101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b10010001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b01100010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b10101100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b11010011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b11000010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b01011100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b00100100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b00000110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b01001001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b00001010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b00111010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b00110010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b11100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b11011011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b00001011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b01011110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b11011110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b00010100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b10111000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b11101110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b01000110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b10001000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b10010000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b00101010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b00100010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b11011100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b01001111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b10000001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b01100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b01110011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b00011001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b01011101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b01100100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b00111101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b01111110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b10100111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b11000100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b00010111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b01000100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b10010111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b01011111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b11101100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b00010011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b00001100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b11001101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b11010010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b11110011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b11111111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b00010000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b00100001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b11011010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b10110110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b10111100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b11110101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b00111000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b10011101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b10010010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b10001111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b01000000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b10100011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b01010001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b10101000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b10011111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b00111100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b01010000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b01111111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b00000010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b11111001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b01000101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b10000101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b00110011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b01001101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b01000011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b11111011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b10101010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b11101111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b11010000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b11001111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b01011000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b01001100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b01001010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b00111001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b10111110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b11001011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b01101010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b01011011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b10110001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b11111100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b00100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b11101101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b00000000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b11010001 ;
      256'b????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b01010011 ;
      256'b???????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b10000100 ;
      256'b??????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b00101111 ;
      256'b?????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b11100011 ;
      256'b????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b00101001 ;
      256'b???????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b10110011 ;
      256'b??????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b11010110 ;
      256'b?????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b00111011 ;
      256'b????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b01010010 ;
      256'b???????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b10100000 ;
      256'b??????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b01011010 ;
      256'b?????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b01101110 ;
      256'b????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b00011011 ;
      256'b???????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b00011010 ;
      256'b??????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b00101100 ;
      256'b?????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b10000011 ;
      256'b????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b00001001 ;
      256'b???????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b01110101 ;
      256'b??????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b10110010 ;
      256'b?????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b00100111 ;
      256'b????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b11101011 ;
      256'b???????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b11100010 ;
      256'b??????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b10000000 ;
      256'b?????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b00010010 ;
      256'b????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b00000111 ;
      256'b???????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b10011010 ;
      256'b??????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b00000101 ;
      256'b?????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b10010110 ;
      256'b????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b00011000 ;
      256'b???????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b11000011 ;
      256'b??????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b00100011 ;
      256'b?????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b11000111 ;
      256'b????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b00000100 ;
      256'b???????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b00010101 ;
      256'b??????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b00110001 ;
      256'b?????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b11011000 ;
      256'b????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b01110001 ;
      256'b???????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b11110001 ;
      256'b??????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b11100101 ;
      256'b?????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b10100101 ;
      256'b????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b00110100 ;
      256'b???????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b11001100 ;
      256'b??????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b11110111 ;
      256'b?????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b00111111 ;
      256'b????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b00110110 ;
      256'b???????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b00100110 ;
      256'b??????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b10010011 ;
      256'b?????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b11111101 ;
      256'b????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b10110111 ;
      256'b???????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b11000000 ;
      256'b??????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b01110010 ;
      256'b?????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b10100100 ;
      256'b????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b10011100 ;
      256'b???????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b10101111 ;
      256'b??????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b10100010 ;
      256'b?????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b11010100 ;
      256'b????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b10101101 ;
      256'b???????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b11110000 ;
      256'b??????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b01000111 ;
      256'b?????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b01011001 ;
      256'b????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b11111010 ;
      256'b???????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b01111101 ;
      256'b??????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b11001001 ;
      256'b?????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b10000010 ;
      256'b????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b11001010 ;
      256'b???????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b01110110 ;
      256'b??????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b10101011 ;
      256'b?????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b11010111 ;
      256'b????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b11111110 ;
      256'b???????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b00101011 ;
      256'b??????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b01100111 ;
      256'b?????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b00000001 ;
      256'b????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b00110000 ;
      256'b???????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b11000101 ;
      256'b??????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b01101111 ;
      256'b?????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b01101011 ;
      256'b????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b11110010 ;
      256'b???1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b01111011 ;
      256'b??1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b01110111 ;
      256'b?1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b01111100 ;
      256'b1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b01100011 ;
      default:
        _1806_ = \t1.t3.s0.out ;
    endcase
  end
  assign _1807_ = state_in[71:64] == 8'b11111111;
  assign _1808_ = state_in[71:64] == 8'b11111110;
  assign _1809_ = state_in[71:64] == 8'b11111101;
  assign _1810_ = state_in[71:64] == 8'b11111100;
  assign _1811_ = state_in[71:64] == 8'b11111011;
  assign _1812_ = state_in[71:64] == 8'b11111010;
  assign _1813_ = state_in[71:64] == 8'b11111001;
  assign _1814_ = state_in[71:64] == 8'b11111000;
  assign _1815_ = state_in[71:64] == 8'b11110111;
  assign _1816_ = state_in[71:64] == 8'b11110110;
  assign _1817_ = state_in[71:64] == 8'b11110101;
  assign _1818_ = state_in[71:64] == 8'b11110100;
  assign _1819_ = state_in[71:64] == 8'b11110011;
  assign _1820_ = state_in[71:64] == 8'b11110010;
  assign _1821_ = state_in[71:64] == 8'b11110001;
  assign _1822_ = state_in[71:64] == 8'b11110000;
  assign _1823_ = state_in[71:64] == 8'b11101111;
  assign _1824_ = state_in[71:64] == 8'b11101110;
  assign _1825_ = state_in[71:64] == 8'b11101101;
  assign _1826_ = state_in[71:64] == 8'b11101100;
  assign _1827_ = state_in[71:64] == 8'b11101011;
  assign _1828_ = state_in[71:64] == 8'b11101010;
  assign _1829_ = state_in[71:64] == 8'b11101001;
  assign _1830_ = state_in[71:64] == 8'b11101000;
  assign _1831_ = state_in[71:64] == 8'b11100111;
  assign _1832_ = state_in[71:64] == 8'b11100110;
  assign _1833_ = state_in[71:64] == 8'b11100101;
  assign _1834_ = state_in[71:64] == 8'b11100100;
  assign _1835_ = state_in[71:64] == 8'b11100011;
  assign _1836_ = state_in[71:64] == 8'b11100010;
  assign _1837_ = state_in[71:64] == 8'b11100001;
  assign _1838_ = state_in[71:64] == 8'b11100000;
  assign _1839_ = state_in[71:64] == 8'b11011111;
  assign _1840_ = state_in[71:64] == 8'b11011110;
  assign _1841_ = state_in[71:64] == 8'b11011101;
  assign _1842_ = state_in[71:64] == 8'b11011100;
  assign _1843_ = state_in[71:64] == 8'b11011011;
  assign _1844_ = state_in[71:64] == 8'b11011010;
  assign _1845_ = state_in[71:64] == 8'b11011001;
  assign _1846_ = state_in[71:64] == 8'b11011000;
  assign _1847_ = state_in[71:64] == 8'b11010111;
  assign _1848_ = state_in[71:64] == 8'b11010110;
  assign _1849_ = state_in[71:64] == 8'b11010101;
  assign _1850_ = state_in[71:64] == 8'b11010100;
  assign _1851_ = state_in[71:64] == 8'b11010011;
  assign _1852_ = state_in[71:64] == 8'b11010010;
  assign _1853_ = state_in[71:64] == 8'b11010001;
  assign _1854_ = state_in[71:64] == 8'b11010000;
  assign _1855_ = state_in[71:64] == 8'b11001111;
  assign _1856_ = state_in[71:64] == 8'b11001110;
  assign _1857_ = state_in[71:64] == 8'b11001101;
  assign _1858_ = state_in[71:64] == 8'b11001100;
  assign _1859_ = state_in[71:64] == 8'b11001011;
  assign _1860_ = state_in[71:64] == 8'b11001010;
  assign _1861_ = state_in[71:64] == 8'b11001001;
  assign _1862_ = state_in[71:64] == 8'b11001000;
  assign _1863_ = state_in[71:64] == 8'b11000111;
  assign _1864_ = state_in[71:64] == 8'b11000110;
  assign _1865_ = state_in[71:64] == 8'b11000101;
  assign _1866_ = state_in[71:64] == 8'b11000100;
  assign _1867_ = state_in[71:64] == 8'b11000011;
  assign _1868_ = state_in[71:64] == 8'b11000010;
  assign _1869_ = state_in[71:64] == 8'b11000001;
  assign _1870_ = state_in[71:64] == 8'b11000000;
  assign _1871_ = state_in[71:64] == 8'b10111111;
  assign _1872_ = state_in[71:64] == 8'b10111110;
  assign _1873_ = state_in[71:64] == 8'b10111101;
  assign _1874_ = state_in[71:64] == 8'b10111100;
  assign _1875_ = state_in[71:64] == 8'b10111011;
  assign _1876_ = state_in[71:64] == 8'b10111010;
  assign _1877_ = state_in[71:64] == 8'b10111001;
  assign _1878_ = state_in[71:64] == 8'b10111000;
  assign _1879_ = state_in[71:64] == 8'b10110111;
  assign _1880_ = state_in[71:64] == 8'b10110110;
  assign _1881_ = state_in[71:64] == 8'b10110101;
  assign _1882_ = state_in[71:64] == 8'b10110100;
  assign _1883_ = state_in[71:64] == 8'b10110011;
  assign _1884_ = state_in[71:64] == 8'b10110010;
  assign _1885_ = state_in[71:64] == 8'b10110001;
  assign _1886_ = state_in[71:64] == 8'b10110000;
  assign _1887_ = state_in[71:64] == 8'b10101111;
  assign _1888_ = state_in[71:64] == 8'b10101110;
  assign _1889_ = state_in[71:64] == 8'b10101101;
  assign _1890_ = state_in[71:64] == 8'b10101100;
  assign _1891_ = state_in[71:64] == 8'b10101011;
  assign _1892_ = state_in[71:64] == 8'b10101010;
  assign _1893_ = state_in[71:64] == 8'b10101001;
  assign _1894_ = state_in[71:64] == 8'b10101000;
  assign _1895_ = state_in[71:64] == 8'b10100111;
  assign _1896_ = state_in[71:64] == 8'b10100110;
  assign _1897_ = state_in[71:64] == 8'b10100101;
  assign _1898_ = state_in[71:64] == 8'b10100100;
  assign _1899_ = state_in[71:64] == 8'b10100011;
  assign _1900_ = state_in[71:64] == 8'b10100010;
  assign _1901_ = state_in[71:64] == 8'b10100001;
  assign _1902_ = state_in[71:64] == 8'b10100000;
  assign _1903_ = state_in[71:64] == 8'b10011111;
  assign _1904_ = state_in[71:64] == 8'b10011110;
  assign _1905_ = state_in[71:64] == 8'b10011101;
  assign _1906_ = state_in[71:64] == 8'b10011100;
  assign _1907_ = state_in[71:64] == 8'b10011011;
  assign _1908_ = state_in[71:64] == 8'b10011010;
  assign _1909_ = state_in[71:64] == 8'b10011001;
  assign _1910_ = state_in[71:64] == 8'b10011000;
  assign _1911_ = state_in[71:64] == 8'b10010111;
  assign _1912_ = state_in[71:64] == 8'b10010110;
  assign _1913_ = state_in[71:64] == 8'b10010101;
  assign _1914_ = state_in[71:64] == 8'b10010100;
  assign _1915_ = state_in[71:64] == 8'b10010011;
  assign _1916_ = state_in[71:64] == 8'b10010010;
  assign _1917_ = state_in[71:64] == 8'b10010001;
  assign _1918_ = state_in[71:64] == 8'b10010000;
  assign _1919_ = state_in[71:64] == 8'b10001111;
  assign _1920_ = state_in[71:64] == 8'b10001110;
  assign _1921_ = state_in[71:64] == 8'b10001101;
  assign _1922_ = state_in[71:64] == 8'b10001100;
  assign _1923_ = state_in[71:64] == 8'b10001011;
  assign _1924_ = state_in[71:64] == 8'b10001010;
  assign _1925_ = state_in[71:64] == 8'b10001001;
  assign _1926_ = state_in[71:64] == 8'b10001000;
  assign _1927_ = state_in[71:64] == 8'b10000111;
  assign _1928_ = state_in[71:64] == 8'b10000110;
  assign _1929_ = state_in[71:64] == 8'b10000101;
  assign _1930_ = state_in[71:64] == 8'b10000100;
  assign _1931_ = state_in[71:64] == 8'b10000011;
  assign _1932_ = state_in[71:64] == 8'b10000010;
  assign _1933_ = state_in[71:64] == 8'b10000001;
  assign _1934_ = state_in[71:64] == 8'b10000000;
  assign _1935_ = state_in[71:64] == 7'b1111111;
  assign _1936_ = state_in[71:64] == 7'b1111110;
  assign _1937_ = state_in[71:64] == 7'b1111101;
  assign _1938_ = state_in[71:64] == 7'b1111100;
  assign _1939_ = state_in[71:64] == 7'b1111011;
  assign _1940_ = state_in[71:64] == 7'b1111010;
  assign _1941_ = state_in[71:64] == 7'b1111001;
  assign _1942_ = state_in[71:64] == 7'b1111000;
  assign _1943_ = state_in[71:64] == 7'b1110111;
  assign _1944_ = state_in[71:64] == 7'b1110110;
  assign _1945_ = state_in[71:64] == 7'b1110101;
  assign _1946_ = state_in[71:64] == 7'b1110100;
  assign _1947_ = state_in[71:64] == 7'b1110011;
  assign _1948_ = state_in[71:64] == 7'b1110010;
  assign _1949_ = state_in[71:64] == 7'b1110001;
  assign _1950_ = state_in[71:64] == 7'b1110000;
  assign _1951_ = state_in[71:64] == 7'b1101111;
  assign _1952_ = state_in[71:64] == 7'b1101110;
  assign _1953_ = state_in[71:64] == 7'b1101101;
  assign _1954_ = state_in[71:64] == 7'b1101100;
  assign _1955_ = state_in[71:64] == 7'b1101011;
  assign _1956_ = state_in[71:64] == 7'b1101010;
  assign _1957_ = state_in[71:64] == 7'b1101001;
  assign _1958_ = state_in[71:64] == 7'b1101000;
  assign _1959_ = state_in[71:64] == 7'b1100111;
  assign _1960_ = state_in[71:64] == 7'b1100110;
  assign _1961_ = state_in[71:64] == 7'b1100101;
  assign _1962_ = state_in[71:64] == 7'b1100100;
  assign _1963_ = state_in[71:64] == 7'b1100011;
  assign _1964_ = state_in[71:64] == 7'b1100010;
  assign _1965_ = state_in[71:64] == 7'b1100001;
  assign _1966_ = state_in[71:64] == 7'b1100000;
  assign _1967_ = state_in[71:64] == 7'b1011111;
  assign _1968_ = state_in[71:64] == 7'b1011110;
  assign _1969_ = state_in[71:64] == 7'b1011101;
  assign _1970_ = state_in[71:64] == 7'b1011100;
  assign _1971_ = state_in[71:64] == 7'b1011011;
  assign _1972_ = state_in[71:64] == 7'b1011010;
  assign _1973_ = state_in[71:64] == 7'b1011001;
  assign _1974_ = state_in[71:64] == 7'b1011000;
  assign _1975_ = state_in[71:64] == 7'b1010111;
  assign _1976_ = state_in[71:64] == 7'b1010110;
  assign _1977_ = state_in[71:64] == 7'b1010101;
  assign _1978_ = state_in[71:64] == 7'b1010100;
  assign _1979_ = state_in[71:64] == 7'b1010011;
  assign _1980_ = state_in[71:64] == 7'b1010010;
  assign _1981_ = state_in[71:64] == 7'b1010001;
  assign _1982_ = state_in[71:64] == 7'b1010000;
  assign _1983_ = state_in[71:64] == 7'b1001111;
  assign _1984_ = state_in[71:64] == 7'b1001110;
  assign _1985_ = state_in[71:64] == 7'b1001101;
  assign _1986_ = state_in[71:64] == 7'b1001100;
  assign _1987_ = state_in[71:64] == 7'b1001011;
  assign _1988_ = state_in[71:64] == 7'b1001010;
  assign _1989_ = state_in[71:64] == 7'b1001001;
  assign _1990_ = state_in[71:64] == 7'b1001000;
  assign _1991_ = state_in[71:64] == 7'b1000111;
  assign _1992_ = state_in[71:64] == 7'b1000110;
  assign _1993_ = state_in[71:64] == 7'b1000101;
  assign _1994_ = state_in[71:64] == 7'b1000100;
  assign _1995_ = state_in[71:64] == 7'b1000011;
  assign _1996_ = state_in[71:64] == 7'b1000010;
  assign _1997_ = state_in[71:64] == 7'b1000001;
  assign _1998_ = state_in[71:64] == 7'b1000000;
  assign _1999_ = state_in[71:64] == 6'b111111;
  assign _2000_ = state_in[71:64] == 6'b111110;
  assign _2001_ = state_in[71:64] == 6'b111101;
  assign _2002_ = state_in[71:64] == 6'b111100;
  assign _2003_ = state_in[71:64] == 6'b111011;
  assign _2004_ = state_in[71:64] == 6'b111010;
  assign _2005_ = state_in[71:64] == 6'b111001;
  assign _2006_ = state_in[71:64] == 6'b111000;
  assign _2007_ = state_in[71:64] == 6'b110111;
  assign _2008_ = state_in[71:64] == 6'b110110;
  assign _2009_ = state_in[71:64] == 6'b110101;
  assign _2010_ = state_in[71:64] == 6'b110100;
  assign _2011_ = state_in[71:64] == 6'b110011;
  assign _2012_ = state_in[71:64] == 6'b110010;
  assign _2013_ = state_in[71:64] == 6'b110001;
  assign _2014_ = state_in[71:64] == 6'b110000;
  assign _2015_ = state_in[71:64] == 6'b101111;
  assign _2016_ = state_in[71:64] == 6'b101110;
  assign _2017_ = state_in[71:64] == 6'b101101;
  assign _2018_ = state_in[71:64] == 6'b101100;
  assign _2019_ = state_in[71:64] == 6'b101011;
  assign _2020_ = state_in[71:64] == 6'b101010;
  assign _2021_ = state_in[71:64] == 6'b101001;
  assign _2022_ = state_in[71:64] == 6'b101000;
  assign _2023_ = state_in[71:64] == 6'b100111;
  assign _2024_ = state_in[71:64] == 6'b100110;
  assign _2025_ = state_in[71:64] == 6'b100101;
  assign _2026_ = state_in[71:64] == 6'b100100;
  assign _2027_ = state_in[71:64] == 6'b100011;
  assign _2028_ = state_in[71:64] == 6'b100010;
  assign _2029_ = state_in[71:64] == 6'b100001;
  assign _2030_ = state_in[71:64] == 6'b100000;
  assign _2031_ = state_in[71:64] == 5'b11111;
  assign _2032_ = state_in[71:64] == 5'b11110;
  assign _2033_ = state_in[71:64] == 5'b11101;
  assign _2034_ = state_in[71:64] == 5'b11100;
  assign _2035_ = state_in[71:64] == 5'b11011;
  assign _2036_ = state_in[71:64] == 5'b11010;
  assign _2037_ = state_in[71:64] == 5'b11001;
  assign _2038_ = state_in[71:64] == 5'b11000;
  assign _2039_ = state_in[71:64] == 5'b10111;
  assign _2040_ = state_in[71:64] == 5'b10110;
  assign _2041_ = state_in[71:64] == 5'b10101;
  assign _2042_ = state_in[71:64] == 5'b10100;
  assign _2043_ = state_in[71:64] == 5'b10011;
  assign _2044_ = state_in[71:64] == 5'b10010;
  assign _2045_ = state_in[71:64] == 5'b10001;
  assign _2046_ = state_in[71:64] == 5'b10000;
  assign _2047_ = state_in[71:64] == 4'b1111;
  assign _2048_ = state_in[71:64] == 4'b1110;
  assign _2049_ = state_in[71:64] == 4'b1101;
  assign _2050_ = state_in[71:64] == 4'b1100;
  assign _2051_ = state_in[71:64] == 4'b1011;
  assign _2052_ = state_in[71:64] == 4'b1010;
  assign _2053_ = state_in[71:64] == 4'b1001;
  assign _2054_ = state_in[71:64] == 4'b1000;
  assign _2055_ = state_in[71:64] == 3'b111;
  assign _2056_ = state_in[71:64] == 3'b110;
  assign _2057_ = state_in[71:64] == 3'b101;
  assign _2058_ = state_in[71:64] == 3'b100;
  assign _2059_ = state_in[71:64] == 2'b11;
  assign _2060_ = state_in[71:64] == 2'b10;
  assign _2061_ = state_in[71:64] == 1'b1;
  assign _2062_ = ! state_in[71:64];
  always @(posedge clk)
      \t1.t3.s4.out <= _2063_;
  wire [255:0] fangyuan16;
  assign fangyuan16 = { _2062_, _2061_, _2060_, _2059_, _2058_, _2057_, _2056_, _2055_, _2054_, _2053_, _2052_, _2051_, _2050_, _2049_, _2048_, _2047_, _2046_, _2045_, _2044_, _2043_, _2042_, _2041_, _2040_, _2039_, _2038_, _2037_, _2036_, _2035_, _2034_, _2033_, _2032_, _2031_, _2030_, _2029_, _2028_, _2027_, _2026_, _2025_, _2024_, _2023_, _2022_, _2021_, _2020_, _2019_, _2018_, _2017_, _2016_, _2015_, _2014_, _2013_, _2012_, _2011_, _2010_, _2009_, _2008_, _2007_, _2006_, _2005_, _2004_, _2003_, _2002_, _2001_, _2000_, _1999_, _1998_, _1997_, _1996_, _1995_, _1994_, _1993_, _1992_, _1991_, _1990_, _1989_, _1988_, _1987_, _1986_, _1985_, _1984_, _1983_, _1982_, _1981_, _1980_, _1979_, _1978_, _1977_, _1976_, _1975_, _1974_, _1973_, _1972_, _1971_, _1970_, _1969_, _1968_, _1967_, _1966_, _1965_, _1964_, _1963_, _1962_, _1961_, _1960_, _1959_, _1958_, _1957_, _1956_, _1955_, _1954_, _1953_, _1952_, _1951_, _1950_, _1949_, _1948_, _1947_, _1946_, _1945_, _1944_, _1943_, _1942_, _1941_, _1940_, _1939_, _1938_, _1937_, _1936_, _1935_, _1934_, _1933_, _1932_, _1931_, _1930_, _1929_, _1928_, _1927_, _1926_, _1925_, _1924_, _1923_, _1922_, _1921_, _1920_, _1919_, _1918_, _1917_, _1916_, _1915_, _1914_, _1913_, _1912_, _1911_, _1910_, _1909_, _1908_, _1907_, _1906_, _1905_, _1904_, _1903_, _1902_, _1901_, _1900_, _1899_, _1898_, _1897_, _1896_, _1895_, _1894_, _1893_, _1892_, _1891_, _1890_, _1889_, _1888_, _1887_, _1886_, _1885_, _1884_, _1883_, _1882_, _1881_, _1880_, _1879_, _1878_, _1877_, _1876_, _1875_, _1874_, _1873_, _1872_, _1871_, _1870_, _1869_, _1868_, _1867_, _1866_, _1865_, _1864_, _1863_, _1862_, _1861_, _1860_, _1859_, _1858_, _1857_, _1856_, _1855_, _1854_, _1853_, _1852_, _1851_, _1850_, _1849_, _1848_, _1847_, _1846_, _1845_, _1844_, _1843_, _1842_, _1841_, _1840_, _1839_, _1838_, _1837_, _1836_, _1835_, _1834_, _1833_, _1832_, _1831_, _1830_, _1829_, _1828_, _1827_, _1826_, _1825_, _1824_, _1823_, _1822_, _1821_, _1820_, _1819_, _1818_, _1817_, _1816_, _1815_, _1814_, _1813_, _1812_, _1811_, _1810_, _1809_, _1808_, _1807_ };

  always @(\t1.t3.s4.out or fangyuan16) begin
    casez (fangyuan16)
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1 :
        _2063_ = 8'b00101100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1? :
        _2063_ = 8'b01101101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?? :
        _2063_ = 8'b10101000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??? :
        _2063_ = 8'b01111011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???? :
        _2063_ = 8'b00011110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????? :
        _2063_ = 8'b01011010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????? :
        _2063_ = 8'b00101001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????? :
        _2063_ = 8'b10000010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????? :
        _2063_ = 8'b11010000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????? :
        _2063_ = 8'b10000100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????? :
        _2063_ = 8'b11010111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????? :
        _2063_ = 8'b01100101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????? :
        _2063_ = 8'b00011010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????? :
        _2063_ = 8'b00001001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????? :
        _2063_ = 8'b01011001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????? :
        _2063_ = 8'b00000011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????? :
        _2063_ = 8'b10100101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????? :
        _2063_ = 8'b01010000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????? :
        _2063_ = 8'b10101010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????? :
        _2063_ = 8'b10000111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????? :
        _2063_ = 8'b11001001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????? :
        _2063_ = 8'b00010101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????? :
        _2063_ = 8'b00111100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????? :
        _2063_ = 8'b00101101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????? :
        _2063_ = 8'b00110011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????? :
        _2063_ = 8'b00000111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????? :
        _2063_ = 8'b10101001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????? :
        _2063_ = 8'b11010010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????? :
        _2063_ = 8'b00100010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????? :
        _2063_ = 8'b00101011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????? :
        _2063_ = 8'b11101011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????? :
        _2063_ = 8'b11011001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????? :
        _2063_ = 8'b00100111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????? :
        _2063_ = 8'b00111010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????? :
        _2063_ = 8'b10011001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????? :
        _2063_ = 8'b00010111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????? :
        _2063_ = 8'b01101001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????? :
        _2063_ = 8'b10101110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????? :
        _2063_ = 8'b01101010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????? :
        _2063_ = 8'b11000010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????? :
        _2063_ = 8'b00011100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????? :
        _2063_ = 8'b11110111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????? :
        _2063_ = 8'b00000110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????? :
        _2063_ = 8'b10010000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????? :
        _2063_ = 8'b11001100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????? :
        _2063_ = 8'b01110001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????? :
        _2063_ = 8'b01111100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????? :
        _2063_ = 8'b11100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????? :
        _2063_ = 8'b00001111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????? :
        _2063_ = 8'b00001101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????? :
        _2063_ = 8'b01100001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????? :
        _2063_ = 8'b10010110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????? :
        _2063_ = 8'b00111110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????? :
        _2063_ = 8'b11101000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????? :
        _2063_ = 8'b10100001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????? :
        _2063_ = 8'b11001011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????? :
        _2063_ = 8'b10010111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????? :
        _2063_ = 8'b01110011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????? :
        _2063_ = 8'b01010111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????? :
        _2063_ = 8'b00111000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????? :
        _2063_ = 8'b01011100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????? :
        _2063_ = 8'b01001010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????? :
        _2063_ = 8'b11110000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????? :
        _2063_ = 8'b01101111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????? :
        _2063_ = 8'b00010000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b01000111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b11110100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b11001010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b11001111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b11110011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b10101100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b11011000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b01001001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b10011100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b10110001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b00000001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b11011010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b01101110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b10001011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b11010101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b11110010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b11010011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b00110001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b00111001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b11000100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b01000011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b10111101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b10011111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b10111000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b01001000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b00001100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b10010010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b00010100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b01110100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b01100100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b11011011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b10101101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b00010110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b10111100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b10100111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b00101000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b01101011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b11000111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b10001100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b00001011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b00111011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b01010100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b01000100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b10100011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b10011110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b00011001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b11000000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b11100110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b00110010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b10111010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b11001000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b01111010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b11111100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b01010101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b10010011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b00101110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b10001000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b00110101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b10111110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b11000011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b00100110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b00011000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b10000001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b10111111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b11111101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b11100101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b00100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b01000010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b10101111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b01110111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b01100011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b11110001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b01110000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b00100001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b00111111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b00000101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b10000000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b01011101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b10100010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b01001011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b00100101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b01111000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b10100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b11111110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b00000100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b11101001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b10001010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b00010001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b01100110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b10011010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b10000110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b11101101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b01001111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b11000101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b10111011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b10000101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b10110000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b10011000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b10010100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b01110010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b01100111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b10001101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b11010100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b10110110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b01111001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b11100011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b01000000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b11000001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b00000000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b10111001 ;
      256'b????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b10100110 ;
      256'b???????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b00010011 ;
      256'b??????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b01011110 ;
      256'b?????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b11011101 ;
      256'b????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b01010010 ;
      256'b???????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b01111101 ;
      256'b??????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b10110111 ;
      256'b?????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b01110110 ;
      256'b????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b10100100 ;
      256'b???????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b01011011 ;
      256'b??????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b10110100 ;
      256'b?????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b11011100 ;
      256'b????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b00110110 ;
      256'b???????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b00110100 ;
      256'b??????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b01011000 ;
      256'b?????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b00011101 ;
      256'b????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b00010010 ;
      256'b???????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b11101010 ;
      256'b??????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b01111111 ;
      256'b?????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b01001110 ;
      256'b????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b11001101 ;
      256'b???????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b11011111 ;
      256'b??????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b00011011 ;
      256'b?????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b00100100 ;
      256'b????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b00001110 ;
      256'b???????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b00101111 ;
      256'b??????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b00001010 ;
      256'b?????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b00110111 ;
      256'b????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b00110000 ;
      256'b???????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b10011101 ;
      256'b??????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b01000110 ;
      256'b?????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b10010101 ;
      256'b????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b00001000 ;
      256'b???????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b00101010 ;
      256'b??????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b01100010 ;
      256'b?????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b10101011 ;
      256'b????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b11100010 ;
      256'b???????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b11111001 ;
      256'b??????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b11010001 ;
      256'b?????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b01010001 ;
      256'b????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b01101000 ;
      256'b???????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b10000011 ;
      256'b??????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b11110101 ;
      256'b?????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b01111110 ;
      256'b????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b01101100 ;
      256'b???????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b01001100 ;
      256'b??????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b00111101 ;
      256'b?????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b11100001 ;
      256'b????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b01110101 ;
      256'b???????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b10011011 ;
      256'b??????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b11100100 ;
      256'b?????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b01010011 ;
      256'b????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b00100011 ;
      256'b???????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b01000101 ;
      256'b??????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b01011111 ;
      256'b?????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b10110011 ;
      256'b????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b01000001 ;
      256'b???????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b11111011 ;
      256'b??????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b10001110 ;
      256'b?????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b10110010 ;
      256'b????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b11101111 ;
      256'b???????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b11111010 ;
      256'b??????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b10001001 ;
      256'b?????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b00011111 ;
      256'b????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b10001111 ;
      256'b???????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b11101100 ;
      256'b??????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b01001101 ;
      256'b?????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b10110101 ;
      256'b????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b11100111 ;
      256'b???????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b01010110 ;
      256'b??????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b11001110 ;
      256'b?????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b00000010 ;
      256'b????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b01100000 ;
      256'b???????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b10010001 ;
      256'b??????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b11011110 ;
      256'b?????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b11010110 ;
      256'b????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b11111111 ;
      256'b???1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b11110110 ;
      256'b??1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b11101110 ;
      256'b?1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b11111000 ;
      256'b1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b11000110 ;
      default:
        _2063_ = \t1.t3.s4.out ;
    endcase
  end
  assign p20[7:0] = \t2.t0.s0.out ^ \t2.t0.s4.out ;
  always @(posedge clk)
      \t2.t0.s0.out <= _2064_;
  wire [255:0] fangyuan17;
  assign fangyuan17 = { _2320_, _2319_, _2318_, _2317_, _2316_, _2315_, _2314_, _2313_, _2312_, _2311_, _2310_, _2309_, _2308_, _2307_, _2306_, _2305_, _2304_, _2303_, _2302_, _2301_, _2300_, _2299_, _2298_, _2297_, _2296_, _2295_, _2294_, _2293_, _2292_, _2291_, _2290_, _2289_, _2288_, _2287_, _2286_, _2285_, _2284_, _2283_, _2282_, _2281_, _2280_, _2279_, _2278_, _2277_, _2276_, _2275_, _2274_, _2273_, _2272_, _2271_, _2270_, _2269_, _2268_, _2267_, _2266_, _2265_, _2264_, _2263_, _2262_, _2261_, _2260_, _2259_, _2258_, _2257_, _2256_, _2255_, _2254_, _2253_, _2252_, _2251_, _2250_, _2249_, _2248_, _2247_, _2246_, _2245_, _2244_, _2243_, _2242_, _2241_, _2240_, _2239_, _2238_, _2237_, _2236_, _2235_, _2234_, _2233_, _2232_, _2231_, _2230_, _2229_, _2228_, _2227_, _2226_, _2225_, _2224_, _2223_, _2222_, _2221_, _2220_, _2219_, _2218_, _2217_, _2216_, _2215_, _2214_, _2213_, _2212_, _2211_, _2210_, _2209_, _2208_, _2207_, _2206_, _2205_, _2204_, _2203_, _2202_, _2201_, _2200_, _2199_, _2198_, _2197_, _2196_, _2195_, _2194_, _2193_, _2192_, _2191_, _2190_, _2189_, _2188_, _2187_, _2186_, _2185_, _2184_, _2183_, _2182_, _2181_, _2180_, _2179_, _2178_, _2177_, _2176_, _2175_, _2174_, _2173_, _2172_, _2171_, _2170_, _2169_, _2168_, _2167_, _2166_, _2165_, _2164_, _2163_, _2162_, _2161_, _2160_, _2159_, _2158_, _2157_, _2156_, _2155_, _2154_, _2153_, _2152_, _2151_, _2150_, _2149_, _2148_, _2147_, _2146_, _2145_, _2144_, _2143_, _2142_, _2141_, _2140_, _2139_, _2138_, _2137_, _2136_, _2135_, _2134_, _2133_, _2132_, _2131_, _2130_, _2129_, _2128_, _2127_, _2126_, _2125_, _2124_, _2123_, _2122_, _2121_, _2120_, _2119_, _2118_, _2117_, _2116_, _2115_, _2114_, _2113_, _2112_, _2111_, _2110_, _2109_, _2108_, _2107_, _2106_, _2105_, _2104_, _2103_, _2102_, _2101_, _2100_, _2099_, _2098_, _2097_, _2096_, _2095_, _2094_, _2093_, _2092_, _2091_, _2090_, _2089_, _2088_, _2087_, _2086_, _2085_, _2084_, _2083_, _2082_, _2081_, _2080_, _2079_, _2078_, _2077_, _2076_, _2075_, _2074_, _2073_, _2072_, _2071_, _2070_, _2069_, _2068_, _2067_, _2066_, _2065_ };

  always @(\t2.t0.s0.out or fangyuan17) begin
    casez (fangyuan17)
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1 :
        _2064_ = 8'b00010110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1? :
        _2064_ = 8'b10111011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?? :
        _2064_ = 8'b01010100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??? :
        _2064_ = 8'b10110000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???? :
        _2064_ = 8'b00001111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????? :
        _2064_ = 8'b00101101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????? :
        _2064_ = 8'b10011001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????? :
        _2064_ = 8'b01000001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????? :
        _2064_ = 8'b01101000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????? :
        _2064_ = 8'b01000010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????? :
        _2064_ = 8'b11100110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????? :
        _2064_ = 8'b10111111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????? :
        _2064_ = 8'b00001101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????? :
        _2064_ = 8'b10001001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????? :
        _2064_ = 8'b10100001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????? :
        _2064_ = 8'b10001100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????? :
        _2064_ = 8'b11011111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????? :
        _2064_ = 8'b00101000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????? :
        _2064_ = 8'b01010101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????? :
        _2064_ = 8'b11001110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????? :
        _2064_ = 8'b11101001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????? :
        _2064_ = 8'b10000111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????? :
        _2064_ = 8'b00011110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????? :
        _2064_ = 8'b10011011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????? :
        _2064_ = 8'b10010100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????? :
        _2064_ = 8'b10001110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????? :
        _2064_ = 8'b11011001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????? :
        _2064_ = 8'b01101001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????? :
        _2064_ = 8'b00010001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????? :
        _2064_ = 8'b10011000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????? :
        _2064_ = 8'b11111000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????? :
        _2064_ = 8'b11100001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????? :
        _2064_ = 8'b10011110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????? :
        _2064_ = 8'b00011101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????? :
        _2064_ = 8'b11000001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????? :
        _2064_ = 8'b10000110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????? :
        _2064_ = 8'b10111001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????? :
        _2064_ = 8'b01010111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????? :
        _2064_ = 8'b00110101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????? :
        _2064_ = 8'b01100001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????? :
        _2064_ = 8'b00001110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????? :
        _2064_ = 8'b11110110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????? :
        _2064_ = 8'b00000011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????? :
        _2064_ = 8'b01001000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????? :
        _2064_ = 8'b01100110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????? :
        _2064_ = 8'b10110101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????? :
        _2064_ = 8'b00111110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????? :
        _2064_ = 8'b01110000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????? :
        _2064_ = 8'b10001010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????? :
        _2064_ = 8'b10001011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????? :
        _2064_ = 8'b10111101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????? :
        _2064_ = 8'b01001011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????? :
        _2064_ = 8'b00011111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????? :
        _2064_ = 8'b01110100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????? :
        _2064_ = 8'b11011101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????? :
        _2064_ = 8'b11101000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????? :
        _2064_ = 8'b11000110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????? :
        _2064_ = 8'b10110100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????? :
        _2064_ = 8'b10100110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????? :
        _2064_ = 8'b00011100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????? :
        _2064_ = 8'b00101110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????? :
        _2064_ = 8'b00100101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????? :
        _2064_ = 8'b01111000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????? :
        _2064_ = 8'b10111010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????? :
        _2064_ = 8'b00001000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b10101110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b01111010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b01100101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b11101010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b11110100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b01010110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b01101100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b10101001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b01001110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b11010101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b10001101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b01101101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b00110111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b11001000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b11100111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b01111001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b11100100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b10010101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b10010001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b01100010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b10101100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b11010011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b11000010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b01011100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b00100100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b00000110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b01001001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b00001010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b00111010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b00110010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b11100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b11011011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b00001011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b01011110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b11011110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b00010100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b10111000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b11101110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b01000110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b10001000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b10010000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b00101010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b00100010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b11011100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b01001111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b10000001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b01100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b01110011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b00011001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b01011101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b01100100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b00111101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b01111110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b10100111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b11000100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b00010111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b01000100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b10010111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b01011111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b11101100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b00010011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b00001100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b11001101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b11010010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b11110011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b11111111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b00010000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b00100001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b11011010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b10110110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b10111100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b11110101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b00111000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b10011101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b10010010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b10001111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b01000000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b10100011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b01010001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b10101000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b10011111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b00111100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b01010000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b01111111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b00000010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b11111001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b01000101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b10000101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b00110011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b01001101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b01000011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b11111011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b10101010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b11101111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b11010000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b11001111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b01011000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b01001100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b01001010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b00111001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b10111110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b11001011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b01101010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b01011011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b10110001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b11111100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b00100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b11101101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b00000000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b11010001 ;
      256'b????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b01010011 ;
      256'b???????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b10000100 ;
      256'b??????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b00101111 ;
      256'b?????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b11100011 ;
      256'b????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b00101001 ;
      256'b???????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b10110011 ;
      256'b??????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b11010110 ;
      256'b?????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b00111011 ;
      256'b????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b01010010 ;
      256'b???????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b10100000 ;
      256'b??????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b01011010 ;
      256'b?????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b01101110 ;
      256'b????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b00011011 ;
      256'b???????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b00011010 ;
      256'b??????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b00101100 ;
      256'b?????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b10000011 ;
      256'b????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b00001001 ;
      256'b???????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b01110101 ;
      256'b??????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b10110010 ;
      256'b?????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b00100111 ;
      256'b????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b11101011 ;
      256'b???????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b11100010 ;
      256'b??????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b10000000 ;
      256'b?????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b00010010 ;
      256'b????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b00000111 ;
      256'b???????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b10011010 ;
      256'b??????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b00000101 ;
      256'b?????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b10010110 ;
      256'b????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b00011000 ;
      256'b???????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b11000011 ;
      256'b??????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b00100011 ;
      256'b?????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b11000111 ;
      256'b????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b00000100 ;
      256'b???????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b00010101 ;
      256'b??????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b00110001 ;
      256'b?????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b11011000 ;
      256'b????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b01110001 ;
      256'b???????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b11110001 ;
      256'b??????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b11100101 ;
      256'b?????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b10100101 ;
      256'b????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b00110100 ;
      256'b???????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b11001100 ;
      256'b??????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b11110111 ;
      256'b?????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b00111111 ;
      256'b????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b00110110 ;
      256'b???????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b00100110 ;
      256'b??????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b10010011 ;
      256'b?????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b11111101 ;
      256'b????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b10110111 ;
      256'b???????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b11000000 ;
      256'b??????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b01110010 ;
      256'b?????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b10100100 ;
      256'b????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b10011100 ;
      256'b???????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b10101111 ;
      256'b??????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b10100010 ;
      256'b?????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b11010100 ;
      256'b????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b10101101 ;
      256'b???????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b11110000 ;
      256'b??????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b01000111 ;
      256'b?????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b01011001 ;
      256'b????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b11111010 ;
      256'b???????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b01111101 ;
      256'b??????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b11001001 ;
      256'b?????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b10000010 ;
      256'b????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b11001010 ;
      256'b???????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b01110110 ;
      256'b??????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b10101011 ;
      256'b?????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b11010111 ;
      256'b????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b11111110 ;
      256'b???????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b00101011 ;
      256'b??????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b01100111 ;
      256'b?????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b00000001 ;
      256'b????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b00110000 ;
      256'b???????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b11000101 ;
      256'b??????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b01101111 ;
      256'b?????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b01101011 ;
      256'b????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b11110010 ;
      256'b???1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b01111011 ;
      256'b??1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b01110111 ;
      256'b?1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b01111100 ;
      256'b1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b01100011 ;
      default:
        _2064_ = \t2.t0.s0.out ;
    endcase
  end
  assign _2065_ = state_in[63:56] == 8'b11111111;
  assign _2066_ = state_in[63:56] == 8'b11111110;
  assign _2067_ = state_in[63:56] == 8'b11111101;
  assign _2068_ = state_in[63:56] == 8'b11111100;
  assign _2069_ = state_in[63:56] == 8'b11111011;
  assign _2070_ = state_in[63:56] == 8'b11111010;
  assign _2071_ = state_in[63:56] == 8'b11111001;
  assign _2072_ = state_in[63:56] == 8'b11111000;
  assign _2073_ = state_in[63:56] == 8'b11110111;
  assign _2074_ = state_in[63:56] == 8'b11110110;
  assign _2075_ = state_in[63:56] == 8'b11110101;
  assign _2076_ = state_in[63:56] == 8'b11110100;
  assign _2077_ = state_in[63:56] == 8'b11110011;
  assign _2078_ = state_in[63:56] == 8'b11110010;
  assign _2079_ = state_in[63:56] == 8'b11110001;
  assign _2080_ = state_in[63:56] == 8'b11110000;
  assign _2081_ = state_in[63:56] == 8'b11101111;
  assign _2082_ = state_in[63:56] == 8'b11101110;
  assign _2083_ = state_in[63:56] == 8'b11101101;
  assign _2084_ = state_in[63:56] == 8'b11101100;
  assign _2085_ = state_in[63:56] == 8'b11101011;
  assign _2086_ = state_in[63:56] == 8'b11101010;
  assign _2087_ = state_in[63:56] == 8'b11101001;
  assign _2088_ = state_in[63:56] == 8'b11101000;
  assign _2089_ = state_in[63:56] == 8'b11100111;
  assign _2090_ = state_in[63:56] == 8'b11100110;
  assign _2091_ = state_in[63:56] == 8'b11100101;
  assign _2092_ = state_in[63:56] == 8'b11100100;
  assign _2093_ = state_in[63:56] == 8'b11100011;
  assign _2094_ = state_in[63:56] == 8'b11100010;
  assign _2095_ = state_in[63:56] == 8'b11100001;
  assign _2096_ = state_in[63:56] == 8'b11100000;
  assign _2097_ = state_in[63:56] == 8'b11011111;
  assign _2098_ = state_in[63:56] == 8'b11011110;
  assign _2099_ = state_in[63:56] == 8'b11011101;
  assign _2100_ = state_in[63:56] == 8'b11011100;
  assign _2101_ = state_in[63:56] == 8'b11011011;
  assign _2102_ = state_in[63:56] == 8'b11011010;
  assign _2103_ = state_in[63:56] == 8'b11011001;
  assign _2104_ = state_in[63:56] == 8'b11011000;
  assign _2105_ = state_in[63:56] == 8'b11010111;
  assign _2106_ = state_in[63:56] == 8'b11010110;
  assign _2107_ = state_in[63:56] == 8'b11010101;
  assign _2108_ = state_in[63:56] == 8'b11010100;
  assign _2109_ = state_in[63:56] == 8'b11010011;
  assign _2110_ = state_in[63:56] == 8'b11010010;
  assign _2111_ = state_in[63:56] == 8'b11010001;
  assign _2112_ = state_in[63:56] == 8'b11010000;
  assign _2113_ = state_in[63:56] == 8'b11001111;
  assign _2114_ = state_in[63:56] == 8'b11001110;
  assign _2115_ = state_in[63:56] == 8'b11001101;
  assign _2116_ = state_in[63:56] == 8'b11001100;
  assign _2117_ = state_in[63:56] == 8'b11001011;
  assign _2118_ = state_in[63:56] == 8'b11001010;
  assign _2119_ = state_in[63:56] == 8'b11001001;
  assign _2120_ = state_in[63:56] == 8'b11001000;
  assign _2121_ = state_in[63:56] == 8'b11000111;
  assign _2122_ = state_in[63:56] == 8'b11000110;
  assign _2123_ = state_in[63:56] == 8'b11000101;
  assign _2124_ = state_in[63:56] == 8'b11000100;
  assign _2125_ = state_in[63:56] == 8'b11000011;
  assign _2126_ = state_in[63:56] == 8'b11000010;
  assign _2127_ = state_in[63:56] == 8'b11000001;
  assign _2128_ = state_in[63:56] == 8'b11000000;
  assign _2129_ = state_in[63:56] == 8'b10111111;
  assign _2130_ = state_in[63:56] == 8'b10111110;
  assign _2131_ = state_in[63:56] == 8'b10111101;
  assign _2132_ = state_in[63:56] == 8'b10111100;
  assign _2133_ = state_in[63:56] == 8'b10111011;
  assign _2134_ = state_in[63:56] == 8'b10111010;
  assign _2135_ = state_in[63:56] == 8'b10111001;
  assign _2136_ = state_in[63:56] == 8'b10111000;
  assign _2137_ = state_in[63:56] == 8'b10110111;
  assign _2138_ = state_in[63:56] == 8'b10110110;
  assign _2139_ = state_in[63:56] == 8'b10110101;
  assign _2140_ = state_in[63:56] == 8'b10110100;
  assign _2141_ = state_in[63:56] == 8'b10110011;
  assign _2142_ = state_in[63:56] == 8'b10110010;
  assign _2143_ = state_in[63:56] == 8'b10110001;
  assign _2144_ = state_in[63:56] == 8'b10110000;
  assign _2145_ = state_in[63:56] == 8'b10101111;
  assign _2146_ = state_in[63:56] == 8'b10101110;
  assign _2147_ = state_in[63:56] == 8'b10101101;
  assign _2148_ = state_in[63:56] == 8'b10101100;
  assign _2149_ = state_in[63:56] == 8'b10101011;
  assign _2150_ = state_in[63:56] == 8'b10101010;
  assign _2151_ = state_in[63:56] == 8'b10101001;
  assign _2152_ = state_in[63:56] == 8'b10101000;
  assign _2153_ = state_in[63:56] == 8'b10100111;
  assign _2154_ = state_in[63:56] == 8'b10100110;
  assign _2155_ = state_in[63:56] == 8'b10100101;
  assign _2156_ = state_in[63:56] == 8'b10100100;
  assign _2157_ = state_in[63:56] == 8'b10100011;
  assign _2158_ = state_in[63:56] == 8'b10100010;
  assign _2159_ = state_in[63:56] == 8'b10100001;
  assign _2160_ = state_in[63:56] == 8'b10100000;
  assign _2161_ = state_in[63:56] == 8'b10011111;
  assign _2162_ = state_in[63:56] == 8'b10011110;
  assign _2163_ = state_in[63:56] == 8'b10011101;
  assign _2164_ = state_in[63:56] == 8'b10011100;
  assign _2165_ = state_in[63:56] == 8'b10011011;
  assign _2166_ = state_in[63:56] == 8'b10011010;
  assign _2167_ = state_in[63:56] == 8'b10011001;
  assign _2168_ = state_in[63:56] == 8'b10011000;
  assign _2169_ = state_in[63:56] == 8'b10010111;
  assign _2170_ = state_in[63:56] == 8'b10010110;
  assign _2171_ = state_in[63:56] == 8'b10010101;
  assign _2172_ = state_in[63:56] == 8'b10010100;
  assign _2173_ = state_in[63:56] == 8'b10010011;
  assign _2174_ = state_in[63:56] == 8'b10010010;
  assign _2175_ = state_in[63:56] == 8'b10010001;
  assign _2176_ = state_in[63:56] == 8'b10010000;
  assign _2177_ = state_in[63:56] == 8'b10001111;
  assign _2178_ = state_in[63:56] == 8'b10001110;
  assign _2179_ = state_in[63:56] == 8'b10001101;
  assign _2180_ = state_in[63:56] == 8'b10001100;
  assign _2181_ = state_in[63:56] == 8'b10001011;
  assign _2182_ = state_in[63:56] == 8'b10001010;
  assign _2183_ = state_in[63:56] == 8'b10001001;
  assign _2184_ = state_in[63:56] == 8'b10001000;
  assign _2185_ = state_in[63:56] == 8'b10000111;
  assign _2186_ = state_in[63:56] == 8'b10000110;
  assign _2187_ = state_in[63:56] == 8'b10000101;
  assign _2188_ = state_in[63:56] == 8'b10000100;
  assign _2189_ = state_in[63:56] == 8'b10000011;
  assign _2190_ = state_in[63:56] == 8'b10000010;
  assign _2191_ = state_in[63:56] == 8'b10000001;
  assign _2192_ = state_in[63:56] == 8'b10000000;
  assign _2193_ = state_in[63:56] == 7'b1111111;
  assign _2194_ = state_in[63:56] == 7'b1111110;
  assign _2195_ = state_in[63:56] == 7'b1111101;
  assign _2196_ = state_in[63:56] == 7'b1111100;
  assign _2197_ = state_in[63:56] == 7'b1111011;
  assign _2198_ = state_in[63:56] == 7'b1111010;
  assign _2199_ = state_in[63:56] == 7'b1111001;
  assign _2200_ = state_in[63:56] == 7'b1111000;
  assign _2201_ = state_in[63:56] == 7'b1110111;
  assign _2202_ = state_in[63:56] == 7'b1110110;
  assign _2203_ = state_in[63:56] == 7'b1110101;
  assign _2204_ = state_in[63:56] == 7'b1110100;
  assign _2205_ = state_in[63:56] == 7'b1110011;
  assign _2206_ = state_in[63:56] == 7'b1110010;
  assign _2207_ = state_in[63:56] == 7'b1110001;
  assign _2208_ = state_in[63:56] == 7'b1110000;
  assign _2209_ = state_in[63:56] == 7'b1101111;
  assign _2210_ = state_in[63:56] == 7'b1101110;
  assign _2211_ = state_in[63:56] == 7'b1101101;
  assign _2212_ = state_in[63:56] == 7'b1101100;
  assign _2213_ = state_in[63:56] == 7'b1101011;
  assign _2214_ = state_in[63:56] == 7'b1101010;
  assign _2215_ = state_in[63:56] == 7'b1101001;
  assign _2216_ = state_in[63:56] == 7'b1101000;
  assign _2217_ = state_in[63:56] == 7'b1100111;
  assign _2218_ = state_in[63:56] == 7'b1100110;
  assign _2219_ = state_in[63:56] == 7'b1100101;
  assign _2220_ = state_in[63:56] == 7'b1100100;
  assign _2221_ = state_in[63:56] == 7'b1100011;
  assign _2222_ = state_in[63:56] == 7'b1100010;
  assign _2223_ = state_in[63:56] == 7'b1100001;
  assign _2224_ = state_in[63:56] == 7'b1100000;
  assign _2225_ = state_in[63:56] == 7'b1011111;
  assign _2226_ = state_in[63:56] == 7'b1011110;
  assign _2227_ = state_in[63:56] == 7'b1011101;
  assign _2228_ = state_in[63:56] == 7'b1011100;
  assign _2229_ = state_in[63:56] == 7'b1011011;
  assign _2230_ = state_in[63:56] == 7'b1011010;
  assign _2231_ = state_in[63:56] == 7'b1011001;
  assign _2232_ = state_in[63:56] == 7'b1011000;
  assign _2233_ = state_in[63:56] == 7'b1010111;
  assign _2234_ = state_in[63:56] == 7'b1010110;
  assign _2235_ = state_in[63:56] == 7'b1010101;
  assign _2236_ = state_in[63:56] == 7'b1010100;
  assign _2237_ = state_in[63:56] == 7'b1010011;
  assign _2238_ = state_in[63:56] == 7'b1010010;
  assign _2239_ = state_in[63:56] == 7'b1010001;
  assign _2240_ = state_in[63:56] == 7'b1010000;
  assign _2241_ = state_in[63:56] == 7'b1001111;
  assign _2242_ = state_in[63:56] == 7'b1001110;
  assign _2243_ = state_in[63:56] == 7'b1001101;
  assign _2244_ = state_in[63:56] == 7'b1001100;
  assign _2245_ = state_in[63:56] == 7'b1001011;
  assign _2246_ = state_in[63:56] == 7'b1001010;
  assign _2247_ = state_in[63:56] == 7'b1001001;
  assign _2248_ = state_in[63:56] == 7'b1001000;
  assign _2249_ = state_in[63:56] == 7'b1000111;
  assign _2250_ = state_in[63:56] == 7'b1000110;
  assign _2251_ = state_in[63:56] == 7'b1000101;
  assign _2252_ = state_in[63:56] == 7'b1000100;
  assign _2253_ = state_in[63:56] == 7'b1000011;
  assign _2254_ = state_in[63:56] == 7'b1000010;
  assign _2255_ = state_in[63:56] == 7'b1000001;
  assign _2256_ = state_in[63:56] == 7'b1000000;
  assign _2257_ = state_in[63:56] == 6'b111111;
  assign _2258_ = state_in[63:56] == 6'b111110;
  assign _2259_ = state_in[63:56] == 6'b111101;
  assign _2260_ = state_in[63:56] == 6'b111100;
  assign _2261_ = state_in[63:56] == 6'b111011;
  assign _2262_ = state_in[63:56] == 6'b111010;
  assign _2263_ = state_in[63:56] == 6'b111001;
  assign _2264_ = state_in[63:56] == 6'b111000;
  assign _2265_ = state_in[63:56] == 6'b110111;
  assign _2266_ = state_in[63:56] == 6'b110110;
  assign _2267_ = state_in[63:56] == 6'b110101;
  assign _2268_ = state_in[63:56] == 6'b110100;
  assign _2269_ = state_in[63:56] == 6'b110011;
  assign _2270_ = state_in[63:56] == 6'b110010;
  assign _2271_ = state_in[63:56] == 6'b110001;
  assign _2272_ = state_in[63:56] == 6'b110000;
  assign _2273_ = state_in[63:56] == 6'b101111;
  assign _2274_ = state_in[63:56] == 6'b101110;
  assign _2275_ = state_in[63:56] == 6'b101101;
  assign _2276_ = state_in[63:56] == 6'b101100;
  assign _2277_ = state_in[63:56] == 6'b101011;
  assign _2278_ = state_in[63:56] == 6'b101010;
  assign _2279_ = state_in[63:56] == 6'b101001;
  assign _2280_ = state_in[63:56] == 6'b101000;
  assign _2281_ = state_in[63:56] == 6'b100111;
  assign _2282_ = state_in[63:56] == 6'b100110;
  assign _2283_ = state_in[63:56] == 6'b100101;
  assign _2284_ = state_in[63:56] == 6'b100100;
  assign _2285_ = state_in[63:56] == 6'b100011;
  assign _2286_ = state_in[63:56] == 6'b100010;
  assign _2287_ = state_in[63:56] == 6'b100001;
  assign _2288_ = state_in[63:56] == 6'b100000;
  assign _2289_ = state_in[63:56] == 5'b11111;
  assign _2290_ = state_in[63:56] == 5'b11110;
  assign _2291_ = state_in[63:56] == 5'b11101;
  assign _2292_ = state_in[63:56] == 5'b11100;
  assign _2293_ = state_in[63:56] == 5'b11011;
  assign _2294_ = state_in[63:56] == 5'b11010;
  assign _2295_ = state_in[63:56] == 5'b11001;
  assign _2296_ = state_in[63:56] == 5'b11000;
  assign _2297_ = state_in[63:56] == 5'b10111;
  assign _2298_ = state_in[63:56] == 5'b10110;
  assign _2299_ = state_in[63:56] == 5'b10101;
  assign _2300_ = state_in[63:56] == 5'b10100;
  assign _2301_ = state_in[63:56] == 5'b10011;
  assign _2302_ = state_in[63:56] == 5'b10010;
  assign _2303_ = state_in[63:56] == 5'b10001;
  assign _2304_ = state_in[63:56] == 5'b10000;
  assign _2305_ = state_in[63:56] == 4'b1111;
  assign _2306_ = state_in[63:56] == 4'b1110;
  assign _2307_ = state_in[63:56] == 4'b1101;
  assign _2308_ = state_in[63:56] == 4'b1100;
  assign _2309_ = state_in[63:56] == 4'b1011;
  assign _2310_ = state_in[63:56] == 4'b1010;
  assign _2311_ = state_in[63:56] == 4'b1001;
  assign _2312_ = state_in[63:56] == 4'b1000;
  assign _2313_ = state_in[63:56] == 3'b111;
  assign _2314_ = state_in[63:56] == 3'b110;
  assign _2315_ = state_in[63:56] == 3'b101;
  assign _2316_ = state_in[63:56] == 3'b100;
  assign _2317_ = state_in[63:56] == 2'b11;
  assign _2318_ = state_in[63:56] == 2'b10;
  assign _2319_ = state_in[63:56] == 1'b1;
  assign _2320_ = ! state_in[63:56];
  always @(posedge clk)
      \t2.t0.s4.out <= _2321_;
  wire [255:0] fangyuan18;
  assign fangyuan18 = { _2320_, _2319_, _2318_, _2317_, _2316_, _2315_, _2314_, _2313_, _2312_, _2311_, _2310_, _2309_, _2308_, _2307_, _2306_, _2305_, _2304_, _2303_, _2302_, _2301_, _2300_, _2299_, _2298_, _2297_, _2296_, _2295_, _2294_, _2293_, _2292_, _2291_, _2290_, _2289_, _2288_, _2287_, _2286_, _2285_, _2284_, _2283_, _2282_, _2281_, _2280_, _2279_, _2278_, _2277_, _2276_, _2275_, _2274_, _2273_, _2272_, _2271_, _2270_, _2269_, _2268_, _2267_, _2266_, _2265_, _2264_, _2263_, _2262_, _2261_, _2260_, _2259_, _2258_, _2257_, _2256_, _2255_, _2254_, _2253_, _2252_, _2251_, _2250_, _2249_, _2248_, _2247_, _2246_, _2245_, _2244_, _2243_, _2242_, _2241_, _2240_, _2239_, _2238_, _2237_, _2236_, _2235_, _2234_, _2233_, _2232_, _2231_, _2230_, _2229_, _2228_, _2227_, _2226_, _2225_, _2224_, _2223_, _2222_, _2221_, _2220_, _2219_, _2218_, _2217_, _2216_, _2215_, _2214_, _2213_, _2212_, _2211_, _2210_, _2209_, _2208_, _2207_, _2206_, _2205_, _2204_, _2203_, _2202_, _2201_, _2200_, _2199_, _2198_, _2197_, _2196_, _2195_, _2194_, _2193_, _2192_, _2191_, _2190_, _2189_, _2188_, _2187_, _2186_, _2185_, _2184_, _2183_, _2182_, _2181_, _2180_, _2179_, _2178_, _2177_, _2176_, _2175_, _2174_, _2173_, _2172_, _2171_, _2170_, _2169_, _2168_, _2167_, _2166_, _2165_, _2164_, _2163_, _2162_, _2161_, _2160_, _2159_, _2158_, _2157_, _2156_, _2155_, _2154_, _2153_, _2152_, _2151_, _2150_, _2149_, _2148_, _2147_, _2146_, _2145_, _2144_, _2143_, _2142_, _2141_, _2140_, _2139_, _2138_, _2137_, _2136_, _2135_, _2134_, _2133_, _2132_, _2131_, _2130_, _2129_, _2128_, _2127_, _2126_, _2125_, _2124_, _2123_, _2122_, _2121_, _2120_, _2119_, _2118_, _2117_, _2116_, _2115_, _2114_, _2113_, _2112_, _2111_, _2110_, _2109_, _2108_, _2107_, _2106_, _2105_, _2104_, _2103_, _2102_, _2101_, _2100_, _2099_, _2098_, _2097_, _2096_, _2095_, _2094_, _2093_, _2092_, _2091_, _2090_, _2089_, _2088_, _2087_, _2086_, _2085_, _2084_, _2083_, _2082_, _2081_, _2080_, _2079_, _2078_, _2077_, _2076_, _2075_, _2074_, _2073_, _2072_, _2071_, _2070_, _2069_, _2068_, _2067_, _2066_, _2065_ };

  always @(\t2.t0.s4.out or fangyuan18) begin
    casez (fangyuan18)
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1 :
        _2321_ = 8'b00101100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1? :
        _2321_ = 8'b01101101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?? :
        _2321_ = 8'b10101000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??? :
        _2321_ = 8'b01111011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???? :
        _2321_ = 8'b00011110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????? :
        _2321_ = 8'b01011010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????? :
        _2321_ = 8'b00101001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????? :
        _2321_ = 8'b10000010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????? :
        _2321_ = 8'b11010000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????? :
        _2321_ = 8'b10000100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????? :
        _2321_ = 8'b11010111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????? :
        _2321_ = 8'b01100101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????? :
        _2321_ = 8'b00011010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????? :
        _2321_ = 8'b00001001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????? :
        _2321_ = 8'b01011001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????? :
        _2321_ = 8'b00000011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????? :
        _2321_ = 8'b10100101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????? :
        _2321_ = 8'b01010000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????? :
        _2321_ = 8'b10101010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????? :
        _2321_ = 8'b10000111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????? :
        _2321_ = 8'b11001001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????? :
        _2321_ = 8'b00010101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????? :
        _2321_ = 8'b00111100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????? :
        _2321_ = 8'b00101101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????? :
        _2321_ = 8'b00110011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????? :
        _2321_ = 8'b00000111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????? :
        _2321_ = 8'b10101001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????? :
        _2321_ = 8'b11010010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????? :
        _2321_ = 8'b00100010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????? :
        _2321_ = 8'b00101011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????? :
        _2321_ = 8'b11101011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????? :
        _2321_ = 8'b11011001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????? :
        _2321_ = 8'b00100111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????? :
        _2321_ = 8'b00111010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????? :
        _2321_ = 8'b10011001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????? :
        _2321_ = 8'b00010111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????? :
        _2321_ = 8'b01101001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????? :
        _2321_ = 8'b10101110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????? :
        _2321_ = 8'b01101010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????? :
        _2321_ = 8'b11000010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????? :
        _2321_ = 8'b00011100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????? :
        _2321_ = 8'b11110111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????? :
        _2321_ = 8'b00000110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????? :
        _2321_ = 8'b10010000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????? :
        _2321_ = 8'b11001100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????? :
        _2321_ = 8'b01110001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????? :
        _2321_ = 8'b01111100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????? :
        _2321_ = 8'b11100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????? :
        _2321_ = 8'b00001111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????? :
        _2321_ = 8'b00001101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????? :
        _2321_ = 8'b01100001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????? :
        _2321_ = 8'b10010110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????? :
        _2321_ = 8'b00111110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????? :
        _2321_ = 8'b11101000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????? :
        _2321_ = 8'b10100001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????? :
        _2321_ = 8'b11001011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????? :
        _2321_ = 8'b10010111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????? :
        _2321_ = 8'b01110011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????? :
        _2321_ = 8'b01010111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????? :
        _2321_ = 8'b00111000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????? :
        _2321_ = 8'b01011100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????? :
        _2321_ = 8'b01001010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????? :
        _2321_ = 8'b11110000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????? :
        _2321_ = 8'b01101111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????? :
        _2321_ = 8'b00010000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b01000111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b11110100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b11001010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b11001111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b11110011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b10101100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b11011000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b01001001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b10011100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b10110001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b00000001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b11011010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b01101110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b10001011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b11010101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b11110010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b11010011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b00110001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b00111001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b11000100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b01000011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b10111101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b10011111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b10111000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b01001000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b00001100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b10010010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b00010100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b01110100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b01100100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b11011011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b10101101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b00010110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b10111100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b10100111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b00101000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b01101011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b11000111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b10001100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b00001011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b00111011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b01010100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b01000100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b10100011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b10011110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b00011001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b11000000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b11100110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b00110010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b10111010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b11001000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b01111010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b11111100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b01010101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b10010011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b00101110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b10001000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b00110101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b10111110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b11000011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b00100110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b00011000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b10000001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b10111111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b11111101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b11100101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b00100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b01000010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b10101111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b01110111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b01100011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b11110001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b01110000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b00100001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b00111111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b00000101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b10000000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b01011101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b10100010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b01001011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b00100101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b01111000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b10100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b11111110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b00000100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b11101001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b10001010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b00010001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b01100110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b10011010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b10000110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b11101101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b01001111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b11000101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b10111011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b10000101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b10110000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b10011000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b10010100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b01110010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b01100111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b10001101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b11010100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b10110110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b01111001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b11100011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b01000000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b11000001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b00000000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b10111001 ;
      256'b????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b10100110 ;
      256'b???????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b00010011 ;
      256'b??????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b01011110 ;
      256'b?????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b11011101 ;
      256'b????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b01010010 ;
      256'b???????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b01111101 ;
      256'b??????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b10110111 ;
      256'b?????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b01110110 ;
      256'b????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b10100100 ;
      256'b???????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b01011011 ;
      256'b??????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b10110100 ;
      256'b?????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b11011100 ;
      256'b????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b00110110 ;
      256'b???????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b00110100 ;
      256'b??????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b01011000 ;
      256'b?????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b00011101 ;
      256'b????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b00010010 ;
      256'b???????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b11101010 ;
      256'b??????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b01111111 ;
      256'b?????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b01001110 ;
      256'b????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b11001101 ;
      256'b???????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b11011111 ;
      256'b??????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b00011011 ;
      256'b?????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b00100100 ;
      256'b????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b00001110 ;
      256'b???????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b00101111 ;
      256'b??????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b00001010 ;
      256'b?????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b00110111 ;
      256'b????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b00110000 ;
      256'b???????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b10011101 ;
      256'b??????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b01000110 ;
      256'b?????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b10010101 ;
      256'b????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b00001000 ;
      256'b???????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b00101010 ;
      256'b??????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b01100010 ;
      256'b?????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b10101011 ;
      256'b????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b11100010 ;
      256'b???????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b11111001 ;
      256'b??????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b11010001 ;
      256'b?????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b01010001 ;
      256'b????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b01101000 ;
      256'b???????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b10000011 ;
      256'b??????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b11110101 ;
      256'b?????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b01111110 ;
      256'b????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b01101100 ;
      256'b???????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b01001100 ;
      256'b??????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b00111101 ;
      256'b?????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b11100001 ;
      256'b????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b01110101 ;
      256'b???????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b10011011 ;
      256'b??????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b11100100 ;
      256'b?????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b01010011 ;
      256'b????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b00100011 ;
      256'b???????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b01000101 ;
      256'b??????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b01011111 ;
      256'b?????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b10110011 ;
      256'b????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b01000001 ;
      256'b???????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b11111011 ;
      256'b??????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b10001110 ;
      256'b?????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b10110010 ;
      256'b????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b11101111 ;
      256'b???????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b11111010 ;
      256'b??????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b10001001 ;
      256'b?????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b00011111 ;
      256'b????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b10001111 ;
      256'b???????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b11101100 ;
      256'b??????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b01001101 ;
      256'b?????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b10110101 ;
      256'b????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b11100111 ;
      256'b???????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b01010110 ;
      256'b??????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b11001110 ;
      256'b?????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b00000010 ;
      256'b????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b01100000 ;
      256'b???????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b10010001 ;
      256'b??????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b11011110 ;
      256'b?????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b11010110 ;
      256'b????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b11111111 ;
      256'b???1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b11110110 ;
      256'b??1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b11101110 ;
      256'b?1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b11111000 ;
      256'b1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b11000110 ;
      default:
        _2321_ = \t2.t0.s4.out ;
    endcase
  end
  assign p21[31:24] = \t2.t1.s0.out ^ \t2.t1.s4.out ;
  always @(posedge clk)
      \t2.t1.s0.out <= _2322_;
  wire [255:0] fangyuan19;
  assign fangyuan19 = { _2578_, _2577_, _2576_, _2575_, _2574_, _2573_, _2572_, _2571_, _2570_, _2569_, _2568_, _2567_, _2566_, _2565_, _2564_, _2563_, _2562_, _2561_, _2560_, _2559_, _2558_, _2557_, _2556_, _2555_, _2554_, _2553_, _2552_, _2551_, _2550_, _2549_, _2548_, _2547_, _2546_, _2545_, _2544_, _2543_, _2542_, _2541_, _2540_, _2539_, _2538_, _2537_, _2536_, _2535_, _2534_, _2533_, _2532_, _2531_, _2530_, _2529_, _2528_, _2527_, _2526_, _2525_, _2524_, _2523_, _2522_, _2521_, _2520_, _2519_, _2518_, _2517_, _2516_, _2515_, _2514_, _2513_, _2512_, _2511_, _2510_, _2509_, _2508_, _2507_, _2506_, _2505_, _2504_, _2503_, _2502_, _2501_, _2500_, _2499_, _2498_, _2497_, _2496_, _2495_, _2494_, _2493_, _2492_, _2491_, _2490_, _2489_, _2488_, _2487_, _2486_, _2485_, _2484_, _2483_, _2482_, _2481_, _2480_, _2479_, _2478_, _2477_, _2476_, _2475_, _2474_, _2473_, _2472_, _2471_, _2470_, _2469_, _2468_, _2467_, _2466_, _2465_, _2464_, _2463_, _2462_, _2461_, _2460_, _2459_, _2458_, _2457_, _2456_, _2455_, _2454_, _2453_, _2452_, _2451_, _2450_, _2449_, _2448_, _2447_, _2446_, _2445_, _2444_, _2443_, _2442_, _2441_, _2440_, _2439_, _2438_, _2437_, _2436_, _2435_, _2434_, _2433_, _2432_, _2431_, _2430_, _2429_, _2428_, _2427_, _2426_, _2425_, _2424_, _2423_, _2422_, _2421_, _2420_, _2419_, _2418_, _2417_, _2416_, _2415_, _2414_, _2413_, _2412_, _2411_, _2410_, _2409_, _2408_, _2407_, _2406_, _2405_, _2404_, _2403_, _2402_, _2401_, _2400_, _2399_, _2398_, _2397_, _2396_, _2395_, _2394_, _2393_, _2392_, _2391_, _2390_, _2389_, _2388_, _2387_, _2386_, _2385_, _2384_, _2383_, _2382_, _2381_, _2380_, _2379_, _2378_, _2377_, _2376_, _2375_, _2374_, _2373_, _2372_, _2371_, _2370_, _2369_, _2368_, _2367_, _2366_, _2365_, _2364_, _2363_, _2362_, _2361_, _2360_, _2359_, _2358_, _2357_, _2356_, _2355_, _2354_, _2353_, _2352_, _2351_, _2350_, _2349_, _2348_, _2347_, _2346_, _2345_, _2344_, _2343_, _2342_, _2341_, _2340_, _2339_, _2338_, _2337_, _2336_, _2335_, _2334_, _2333_, _2332_, _2331_, _2330_, _2329_, _2328_, _2327_, _2326_, _2325_, _2324_, _2323_ };

  always @(\t2.t1.s0.out or fangyuan19) begin
    casez (fangyuan19)
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1 :
        _2322_ = 8'b00010110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1? :
        _2322_ = 8'b10111011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?? :
        _2322_ = 8'b01010100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??? :
        _2322_ = 8'b10110000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???? :
        _2322_ = 8'b00001111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????? :
        _2322_ = 8'b00101101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????? :
        _2322_ = 8'b10011001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????? :
        _2322_ = 8'b01000001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????? :
        _2322_ = 8'b01101000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????? :
        _2322_ = 8'b01000010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????? :
        _2322_ = 8'b11100110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????? :
        _2322_ = 8'b10111111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????? :
        _2322_ = 8'b00001101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????? :
        _2322_ = 8'b10001001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????? :
        _2322_ = 8'b10100001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????? :
        _2322_ = 8'b10001100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????? :
        _2322_ = 8'b11011111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????? :
        _2322_ = 8'b00101000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????? :
        _2322_ = 8'b01010101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????? :
        _2322_ = 8'b11001110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????? :
        _2322_ = 8'b11101001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????? :
        _2322_ = 8'b10000111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????? :
        _2322_ = 8'b00011110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????? :
        _2322_ = 8'b10011011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????? :
        _2322_ = 8'b10010100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????? :
        _2322_ = 8'b10001110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????? :
        _2322_ = 8'b11011001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????? :
        _2322_ = 8'b01101001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????? :
        _2322_ = 8'b00010001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????? :
        _2322_ = 8'b10011000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????? :
        _2322_ = 8'b11111000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????? :
        _2322_ = 8'b11100001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????? :
        _2322_ = 8'b10011110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????? :
        _2322_ = 8'b00011101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????? :
        _2322_ = 8'b11000001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????? :
        _2322_ = 8'b10000110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????? :
        _2322_ = 8'b10111001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????? :
        _2322_ = 8'b01010111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????? :
        _2322_ = 8'b00110101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????? :
        _2322_ = 8'b01100001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????? :
        _2322_ = 8'b00001110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????? :
        _2322_ = 8'b11110110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????? :
        _2322_ = 8'b00000011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????? :
        _2322_ = 8'b01001000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????? :
        _2322_ = 8'b01100110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????? :
        _2322_ = 8'b10110101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????? :
        _2322_ = 8'b00111110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????? :
        _2322_ = 8'b01110000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????? :
        _2322_ = 8'b10001010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????? :
        _2322_ = 8'b10001011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????? :
        _2322_ = 8'b10111101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????? :
        _2322_ = 8'b01001011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????? :
        _2322_ = 8'b00011111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????? :
        _2322_ = 8'b01110100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????? :
        _2322_ = 8'b11011101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????? :
        _2322_ = 8'b11101000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????? :
        _2322_ = 8'b11000110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????? :
        _2322_ = 8'b10110100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????? :
        _2322_ = 8'b10100110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????? :
        _2322_ = 8'b00011100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????? :
        _2322_ = 8'b00101110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????? :
        _2322_ = 8'b00100101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????? :
        _2322_ = 8'b01111000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????? :
        _2322_ = 8'b10111010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????? :
        _2322_ = 8'b00001000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b10101110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b01111010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b01100101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b11101010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b11110100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b01010110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b01101100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b10101001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b01001110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b11010101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b10001101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b01101101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b00110111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b11001000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b11100111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b01111001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b11100100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b10010101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b10010001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b01100010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b10101100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b11010011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b11000010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b01011100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b00100100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b00000110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b01001001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b00001010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b00111010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b00110010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b11100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b11011011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b00001011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b01011110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b11011110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b00010100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b10111000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b11101110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b01000110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b10001000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b10010000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b00101010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b00100010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b11011100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b01001111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b10000001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b01100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b01110011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b00011001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b01011101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b01100100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b00111101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b01111110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b10100111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b11000100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b00010111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b01000100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b10010111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b01011111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b11101100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b00010011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b00001100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b11001101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b11010010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b11110011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b11111111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b00010000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b00100001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b11011010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b10110110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b10111100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b11110101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b00111000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b10011101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b10010010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b10001111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b01000000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b10100011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b01010001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b10101000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b10011111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b00111100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b01010000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b01111111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b00000010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b11111001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b01000101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b10000101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b00110011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b01001101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b01000011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b11111011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b10101010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b11101111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b11010000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b11001111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b01011000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b01001100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b01001010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b00111001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b10111110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b11001011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b01101010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b01011011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b10110001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b11111100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b00100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b11101101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b00000000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b11010001 ;
      256'b????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b01010011 ;
      256'b???????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b10000100 ;
      256'b??????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b00101111 ;
      256'b?????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b11100011 ;
      256'b????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b00101001 ;
      256'b???????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b10110011 ;
      256'b??????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b11010110 ;
      256'b?????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b00111011 ;
      256'b????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b01010010 ;
      256'b???????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b10100000 ;
      256'b??????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b01011010 ;
      256'b?????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b01101110 ;
      256'b????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b00011011 ;
      256'b???????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b00011010 ;
      256'b??????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b00101100 ;
      256'b?????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b10000011 ;
      256'b????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b00001001 ;
      256'b???????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b01110101 ;
      256'b??????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b10110010 ;
      256'b?????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b00100111 ;
      256'b????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b11101011 ;
      256'b???????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b11100010 ;
      256'b??????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b10000000 ;
      256'b?????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b00010010 ;
      256'b????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b00000111 ;
      256'b???????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b10011010 ;
      256'b??????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b00000101 ;
      256'b?????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b10010110 ;
      256'b????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b00011000 ;
      256'b???????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b11000011 ;
      256'b??????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b00100011 ;
      256'b?????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b11000111 ;
      256'b????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b00000100 ;
      256'b???????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b00010101 ;
      256'b??????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b00110001 ;
      256'b?????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b11011000 ;
      256'b????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b01110001 ;
      256'b???????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b11110001 ;
      256'b??????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b11100101 ;
      256'b?????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b10100101 ;
      256'b????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b00110100 ;
      256'b???????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b11001100 ;
      256'b??????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b11110111 ;
      256'b?????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b00111111 ;
      256'b????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b00110110 ;
      256'b???????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b00100110 ;
      256'b??????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b10010011 ;
      256'b?????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b11111101 ;
      256'b????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b10110111 ;
      256'b???????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b11000000 ;
      256'b??????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b01110010 ;
      256'b?????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b10100100 ;
      256'b????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b10011100 ;
      256'b???????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b10101111 ;
      256'b??????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b10100010 ;
      256'b?????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b11010100 ;
      256'b????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b10101101 ;
      256'b???????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b11110000 ;
      256'b??????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b01000111 ;
      256'b?????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b01011001 ;
      256'b????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b11111010 ;
      256'b???????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b01111101 ;
      256'b??????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b11001001 ;
      256'b?????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b10000010 ;
      256'b????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b11001010 ;
      256'b???????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b01110110 ;
      256'b??????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b10101011 ;
      256'b?????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b11010111 ;
      256'b????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b11111110 ;
      256'b???????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b00101011 ;
      256'b??????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b01100111 ;
      256'b?????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b00000001 ;
      256'b????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b00110000 ;
      256'b???????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b11000101 ;
      256'b??????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b01101111 ;
      256'b?????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b01101011 ;
      256'b????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b11110010 ;
      256'b???1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b01111011 ;
      256'b??1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b01110111 ;
      256'b?1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b01111100 ;
      256'b1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b01100011 ;
      default:
        _2322_ = \t2.t1.s0.out ;
    endcase
  end
  assign _2323_ = state_in[55:48] == 8'b11111111;
  assign _2324_ = state_in[55:48] == 8'b11111110;
  assign _2325_ = state_in[55:48] == 8'b11111101;
  assign _2326_ = state_in[55:48] == 8'b11111100;
  assign _2327_ = state_in[55:48] == 8'b11111011;
  assign _2328_ = state_in[55:48] == 8'b11111010;
  assign _2329_ = state_in[55:48] == 8'b11111001;
  assign _2330_ = state_in[55:48] == 8'b11111000;
  assign _2331_ = state_in[55:48] == 8'b11110111;
  assign _2332_ = state_in[55:48] == 8'b11110110;
  assign _2333_ = state_in[55:48] == 8'b11110101;
  assign _2334_ = state_in[55:48] == 8'b11110100;
  assign _2335_ = state_in[55:48] == 8'b11110011;
  assign _2336_ = state_in[55:48] == 8'b11110010;
  assign _2337_ = state_in[55:48] == 8'b11110001;
  assign _2338_ = state_in[55:48] == 8'b11110000;
  assign _2339_ = state_in[55:48] == 8'b11101111;
  assign _2340_ = state_in[55:48] == 8'b11101110;
  assign _2341_ = state_in[55:48] == 8'b11101101;
  assign _2342_ = state_in[55:48] == 8'b11101100;
  assign _2343_ = state_in[55:48] == 8'b11101011;
  assign _2344_ = state_in[55:48] == 8'b11101010;
  assign _2345_ = state_in[55:48] == 8'b11101001;
  assign _2346_ = state_in[55:48] == 8'b11101000;
  assign _2347_ = state_in[55:48] == 8'b11100111;
  assign _2348_ = state_in[55:48] == 8'b11100110;
  assign _2349_ = state_in[55:48] == 8'b11100101;
  assign _2350_ = state_in[55:48] == 8'b11100100;
  assign _2351_ = state_in[55:48] == 8'b11100011;
  assign _2352_ = state_in[55:48] == 8'b11100010;
  assign _2353_ = state_in[55:48] == 8'b11100001;
  assign _2354_ = state_in[55:48] == 8'b11100000;
  assign _2355_ = state_in[55:48] == 8'b11011111;
  assign _2356_ = state_in[55:48] == 8'b11011110;
  assign _2357_ = state_in[55:48] == 8'b11011101;
  assign _2358_ = state_in[55:48] == 8'b11011100;
  assign _2359_ = state_in[55:48] == 8'b11011011;
  assign _2360_ = state_in[55:48] == 8'b11011010;
  assign _2361_ = state_in[55:48] == 8'b11011001;
  assign _2362_ = state_in[55:48] == 8'b11011000;
  assign _2363_ = state_in[55:48] == 8'b11010111;
  assign _2364_ = state_in[55:48] == 8'b11010110;
  assign _2365_ = state_in[55:48] == 8'b11010101;
  assign _2366_ = state_in[55:48] == 8'b11010100;
  assign _2367_ = state_in[55:48] == 8'b11010011;
  assign _2368_ = state_in[55:48] == 8'b11010010;
  assign _2369_ = state_in[55:48] == 8'b11010001;
  assign _2370_ = state_in[55:48] == 8'b11010000;
  assign _2371_ = state_in[55:48] == 8'b11001111;
  assign _2372_ = state_in[55:48] == 8'b11001110;
  assign _2373_ = state_in[55:48] == 8'b11001101;
  assign _2374_ = state_in[55:48] == 8'b11001100;
  assign _2375_ = state_in[55:48] == 8'b11001011;
  assign _2376_ = state_in[55:48] == 8'b11001010;
  assign _2377_ = state_in[55:48] == 8'b11001001;
  assign _2378_ = state_in[55:48] == 8'b11001000;
  assign _2379_ = state_in[55:48] == 8'b11000111;
  assign _2380_ = state_in[55:48] == 8'b11000110;
  assign _2381_ = state_in[55:48] == 8'b11000101;
  assign _2382_ = state_in[55:48] == 8'b11000100;
  assign _2383_ = state_in[55:48] == 8'b11000011;
  assign _2384_ = state_in[55:48] == 8'b11000010;
  assign _2385_ = state_in[55:48] == 8'b11000001;
  assign _2386_ = state_in[55:48] == 8'b11000000;
  assign _2387_ = state_in[55:48] == 8'b10111111;
  assign _2388_ = state_in[55:48] == 8'b10111110;
  assign _2389_ = state_in[55:48] == 8'b10111101;
  assign _2390_ = state_in[55:48] == 8'b10111100;
  assign _2391_ = state_in[55:48] == 8'b10111011;
  assign _2392_ = state_in[55:48] == 8'b10111010;
  assign _2393_ = state_in[55:48] == 8'b10111001;
  assign _2394_ = state_in[55:48] == 8'b10111000;
  assign _2395_ = state_in[55:48] == 8'b10110111;
  assign _2396_ = state_in[55:48] == 8'b10110110;
  assign _2397_ = state_in[55:48] == 8'b10110101;
  assign _2398_ = state_in[55:48] == 8'b10110100;
  assign _2399_ = state_in[55:48] == 8'b10110011;
  assign _2400_ = state_in[55:48] == 8'b10110010;
  assign _2401_ = state_in[55:48] == 8'b10110001;
  assign _2402_ = state_in[55:48] == 8'b10110000;
  assign _2403_ = state_in[55:48] == 8'b10101111;
  assign _2404_ = state_in[55:48] == 8'b10101110;
  assign _2405_ = state_in[55:48] == 8'b10101101;
  assign _2406_ = state_in[55:48] == 8'b10101100;
  assign _2407_ = state_in[55:48] == 8'b10101011;
  assign _2408_ = state_in[55:48] == 8'b10101010;
  assign _2409_ = state_in[55:48] == 8'b10101001;
  assign _2410_ = state_in[55:48] == 8'b10101000;
  assign _2411_ = state_in[55:48] == 8'b10100111;
  assign _2412_ = state_in[55:48] == 8'b10100110;
  assign _2413_ = state_in[55:48] == 8'b10100101;
  assign _2414_ = state_in[55:48] == 8'b10100100;
  assign _2415_ = state_in[55:48] == 8'b10100011;
  assign _2416_ = state_in[55:48] == 8'b10100010;
  assign _2417_ = state_in[55:48] == 8'b10100001;
  assign _2418_ = state_in[55:48] == 8'b10100000;
  assign _2419_ = state_in[55:48] == 8'b10011111;
  assign _2420_ = state_in[55:48] == 8'b10011110;
  assign _2421_ = state_in[55:48] == 8'b10011101;
  assign _2422_ = state_in[55:48] == 8'b10011100;
  assign _2423_ = state_in[55:48] == 8'b10011011;
  assign _2424_ = state_in[55:48] == 8'b10011010;
  assign _2425_ = state_in[55:48] == 8'b10011001;
  assign _2426_ = state_in[55:48] == 8'b10011000;
  assign _2427_ = state_in[55:48] == 8'b10010111;
  assign _2428_ = state_in[55:48] == 8'b10010110;
  assign _2429_ = state_in[55:48] == 8'b10010101;
  assign _2430_ = state_in[55:48] == 8'b10010100;
  assign _2431_ = state_in[55:48] == 8'b10010011;
  assign _2432_ = state_in[55:48] == 8'b10010010;
  assign _2433_ = state_in[55:48] == 8'b10010001;
  assign _2434_ = state_in[55:48] == 8'b10010000;
  assign _2435_ = state_in[55:48] == 8'b10001111;
  assign _2436_ = state_in[55:48] == 8'b10001110;
  assign _2437_ = state_in[55:48] == 8'b10001101;
  assign _2438_ = state_in[55:48] == 8'b10001100;
  assign _2439_ = state_in[55:48] == 8'b10001011;
  assign _2440_ = state_in[55:48] == 8'b10001010;
  assign _2441_ = state_in[55:48] == 8'b10001001;
  assign _2442_ = state_in[55:48] == 8'b10001000;
  assign _2443_ = state_in[55:48] == 8'b10000111;
  assign _2444_ = state_in[55:48] == 8'b10000110;
  assign _2445_ = state_in[55:48] == 8'b10000101;
  assign _2446_ = state_in[55:48] == 8'b10000100;
  assign _2447_ = state_in[55:48] == 8'b10000011;
  assign _2448_ = state_in[55:48] == 8'b10000010;
  assign _2449_ = state_in[55:48] == 8'b10000001;
  assign _2450_ = state_in[55:48] == 8'b10000000;
  assign _2451_ = state_in[55:48] == 7'b1111111;
  assign _2452_ = state_in[55:48] == 7'b1111110;
  assign _2453_ = state_in[55:48] == 7'b1111101;
  assign _2454_ = state_in[55:48] == 7'b1111100;
  assign _2455_ = state_in[55:48] == 7'b1111011;
  assign _2456_ = state_in[55:48] == 7'b1111010;
  assign _2457_ = state_in[55:48] == 7'b1111001;
  assign _2458_ = state_in[55:48] == 7'b1111000;
  assign _2459_ = state_in[55:48] == 7'b1110111;
  assign _2460_ = state_in[55:48] == 7'b1110110;
  assign _2461_ = state_in[55:48] == 7'b1110101;
  assign _2462_ = state_in[55:48] == 7'b1110100;
  assign _2463_ = state_in[55:48] == 7'b1110011;
  assign _2464_ = state_in[55:48] == 7'b1110010;
  assign _2465_ = state_in[55:48] == 7'b1110001;
  assign _2466_ = state_in[55:48] == 7'b1110000;
  assign _2467_ = state_in[55:48] == 7'b1101111;
  assign _2468_ = state_in[55:48] == 7'b1101110;
  assign _2469_ = state_in[55:48] == 7'b1101101;
  assign _2470_ = state_in[55:48] == 7'b1101100;
  assign _2471_ = state_in[55:48] == 7'b1101011;
  assign _2472_ = state_in[55:48] == 7'b1101010;
  assign _2473_ = state_in[55:48] == 7'b1101001;
  assign _2474_ = state_in[55:48] == 7'b1101000;
  assign _2475_ = state_in[55:48] == 7'b1100111;
  assign _2476_ = state_in[55:48] == 7'b1100110;
  assign _2477_ = state_in[55:48] == 7'b1100101;
  assign _2478_ = state_in[55:48] == 7'b1100100;
  assign _2479_ = state_in[55:48] == 7'b1100011;
  assign _2480_ = state_in[55:48] == 7'b1100010;
  assign _2481_ = state_in[55:48] == 7'b1100001;
  assign _2482_ = state_in[55:48] == 7'b1100000;
  assign _2483_ = state_in[55:48] == 7'b1011111;
  assign _2484_ = state_in[55:48] == 7'b1011110;
  assign _2485_ = state_in[55:48] == 7'b1011101;
  assign _2486_ = state_in[55:48] == 7'b1011100;
  assign _2487_ = state_in[55:48] == 7'b1011011;
  assign _2488_ = state_in[55:48] == 7'b1011010;
  assign _2489_ = state_in[55:48] == 7'b1011001;
  assign _2490_ = state_in[55:48] == 7'b1011000;
  assign _2491_ = state_in[55:48] == 7'b1010111;
  assign _2492_ = state_in[55:48] == 7'b1010110;
  assign _2493_ = state_in[55:48] == 7'b1010101;
  assign _2494_ = state_in[55:48] == 7'b1010100;
  assign _2495_ = state_in[55:48] == 7'b1010011;
  assign _2496_ = state_in[55:48] == 7'b1010010;
  assign _2497_ = state_in[55:48] == 7'b1010001;
  assign _2498_ = state_in[55:48] == 7'b1010000;
  assign _2499_ = state_in[55:48] == 7'b1001111;
  assign _2500_ = state_in[55:48] == 7'b1001110;
  assign _2501_ = state_in[55:48] == 7'b1001101;
  assign _2502_ = state_in[55:48] == 7'b1001100;
  assign _2503_ = state_in[55:48] == 7'b1001011;
  assign _2504_ = state_in[55:48] == 7'b1001010;
  assign _2505_ = state_in[55:48] == 7'b1001001;
  assign _2506_ = state_in[55:48] == 7'b1001000;
  assign _2507_ = state_in[55:48] == 7'b1000111;
  assign _2508_ = state_in[55:48] == 7'b1000110;
  assign _2509_ = state_in[55:48] == 7'b1000101;
  assign _2510_ = state_in[55:48] == 7'b1000100;
  assign _2511_ = state_in[55:48] == 7'b1000011;
  assign _2512_ = state_in[55:48] == 7'b1000010;
  assign _2513_ = state_in[55:48] == 7'b1000001;
  assign _2514_ = state_in[55:48] == 7'b1000000;
  assign _2515_ = state_in[55:48] == 6'b111111;
  assign _2516_ = state_in[55:48] == 6'b111110;
  assign _2517_ = state_in[55:48] == 6'b111101;
  assign _2518_ = state_in[55:48] == 6'b111100;
  assign _2519_ = state_in[55:48] == 6'b111011;
  assign _2520_ = state_in[55:48] == 6'b111010;
  assign _2521_ = state_in[55:48] == 6'b111001;
  assign _2522_ = state_in[55:48] == 6'b111000;
  assign _2523_ = state_in[55:48] == 6'b110111;
  assign _2524_ = state_in[55:48] == 6'b110110;
  assign _2525_ = state_in[55:48] == 6'b110101;
  assign _2526_ = state_in[55:48] == 6'b110100;
  assign _2527_ = state_in[55:48] == 6'b110011;
  assign _2528_ = state_in[55:48] == 6'b110010;
  assign _2529_ = state_in[55:48] == 6'b110001;
  assign _2530_ = state_in[55:48] == 6'b110000;
  assign _2531_ = state_in[55:48] == 6'b101111;
  assign _2532_ = state_in[55:48] == 6'b101110;
  assign _2533_ = state_in[55:48] == 6'b101101;
  assign _2534_ = state_in[55:48] == 6'b101100;
  assign _2535_ = state_in[55:48] == 6'b101011;
  assign _2536_ = state_in[55:48] == 6'b101010;
  assign _2537_ = state_in[55:48] == 6'b101001;
  assign _2538_ = state_in[55:48] == 6'b101000;
  assign _2539_ = state_in[55:48] == 6'b100111;
  assign _2540_ = state_in[55:48] == 6'b100110;
  assign _2541_ = state_in[55:48] == 6'b100101;
  assign _2542_ = state_in[55:48] == 6'b100100;
  assign _2543_ = state_in[55:48] == 6'b100011;
  assign _2544_ = state_in[55:48] == 6'b100010;
  assign _2545_ = state_in[55:48] == 6'b100001;
  assign _2546_ = state_in[55:48] == 6'b100000;
  assign _2547_ = state_in[55:48] == 5'b11111;
  assign _2548_ = state_in[55:48] == 5'b11110;
  assign _2549_ = state_in[55:48] == 5'b11101;
  assign _2550_ = state_in[55:48] == 5'b11100;
  assign _2551_ = state_in[55:48] == 5'b11011;
  assign _2552_ = state_in[55:48] == 5'b11010;
  assign _2553_ = state_in[55:48] == 5'b11001;
  assign _2554_ = state_in[55:48] == 5'b11000;
  assign _2555_ = state_in[55:48] == 5'b10111;
  assign _2556_ = state_in[55:48] == 5'b10110;
  assign _2557_ = state_in[55:48] == 5'b10101;
  assign _2558_ = state_in[55:48] == 5'b10100;
  assign _2559_ = state_in[55:48] == 5'b10011;
  assign _2560_ = state_in[55:48] == 5'b10010;
  assign _2561_ = state_in[55:48] == 5'b10001;
  assign _2562_ = state_in[55:48] == 5'b10000;
  assign _2563_ = state_in[55:48] == 4'b1111;
  assign _2564_ = state_in[55:48] == 4'b1110;
  assign _2565_ = state_in[55:48] == 4'b1101;
  assign _2566_ = state_in[55:48] == 4'b1100;
  assign _2567_ = state_in[55:48] == 4'b1011;
  assign _2568_ = state_in[55:48] == 4'b1010;
  assign _2569_ = state_in[55:48] == 4'b1001;
  assign _2570_ = state_in[55:48] == 4'b1000;
  assign _2571_ = state_in[55:48] == 3'b111;
  assign _2572_ = state_in[55:48] == 3'b110;
  assign _2573_ = state_in[55:48] == 3'b101;
  assign _2574_ = state_in[55:48] == 3'b100;
  assign _2575_ = state_in[55:48] == 2'b11;
  assign _2576_ = state_in[55:48] == 2'b10;
  assign _2577_ = state_in[55:48] == 1'b1;
  assign _2578_ = ! state_in[55:48];
  always @(posedge clk)
      \t2.t1.s4.out <= _2579_;
  wire [255:0] fangyuan20;
  assign fangyuan20 = { _2578_, _2577_, _2576_, _2575_, _2574_, _2573_, _2572_, _2571_, _2570_, _2569_, _2568_, _2567_, _2566_, _2565_, _2564_, _2563_, _2562_, _2561_, _2560_, _2559_, _2558_, _2557_, _2556_, _2555_, _2554_, _2553_, _2552_, _2551_, _2550_, _2549_, _2548_, _2547_, _2546_, _2545_, _2544_, _2543_, _2542_, _2541_, _2540_, _2539_, _2538_, _2537_, _2536_, _2535_, _2534_, _2533_, _2532_, _2531_, _2530_, _2529_, _2528_, _2527_, _2526_, _2525_, _2524_, _2523_, _2522_, _2521_, _2520_, _2519_, _2518_, _2517_, _2516_, _2515_, _2514_, _2513_, _2512_, _2511_, _2510_, _2509_, _2508_, _2507_, _2506_, _2505_, _2504_, _2503_, _2502_, _2501_, _2500_, _2499_, _2498_, _2497_, _2496_, _2495_, _2494_, _2493_, _2492_, _2491_, _2490_, _2489_, _2488_, _2487_, _2486_, _2485_, _2484_, _2483_, _2482_, _2481_, _2480_, _2479_, _2478_, _2477_, _2476_, _2475_, _2474_, _2473_, _2472_, _2471_, _2470_, _2469_, _2468_, _2467_, _2466_, _2465_, _2464_, _2463_, _2462_, _2461_, _2460_, _2459_, _2458_, _2457_, _2456_, _2455_, _2454_, _2453_, _2452_, _2451_, _2450_, _2449_, _2448_, _2447_, _2446_, _2445_, _2444_, _2443_, _2442_, _2441_, _2440_, _2439_, _2438_, _2437_, _2436_, _2435_, _2434_, _2433_, _2432_, _2431_, _2430_, _2429_, _2428_, _2427_, _2426_, _2425_, _2424_, _2423_, _2422_, _2421_, _2420_, _2419_, _2418_, _2417_, _2416_, _2415_, _2414_, _2413_, _2412_, _2411_, _2410_, _2409_, _2408_, _2407_, _2406_, _2405_, _2404_, _2403_, _2402_, _2401_, _2400_, _2399_, _2398_, _2397_, _2396_, _2395_, _2394_, _2393_, _2392_, _2391_, _2390_, _2389_, _2388_, _2387_, _2386_, _2385_, _2384_, _2383_, _2382_, _2381_, _2380_, _2379_, _2378_, _2377_, _2376_, _2375_, _2374_, _2373_, _2372_, _2371_, _2370_, _2369_, _2368_, _2367_, _2366_, _2365_, _2364_, _2363_, _2362_, _2361_, _2360_, _2359_, _2358_, _2357_, _2356_, _2355_, _2354_, _2353_, _2352_, _2351_, _2350_, _2349_, _2348_, _2347_, _2346_, _2345_, _2344_, _2343_, _2342_, _2341_, _2340_, _2339_, _2338_, _2337_, _2336_, _2335_, _2334_, _2333_, _2332_, _2331_, _2330_, _2329_, _2328_, _2327_, _2326_, _2325_, _2324_, _2323_ };

  always @(\t2.t1.s4.out or fangyuan20) begin
    casez (fangyuan20)
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1 :
        _2579_ = 8'b00101100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1? :
        _2579_ = 8'b01101101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?? :
        _2579_ = 8'b10101000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??? :
        _2579_ = 8'b01111011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???? :
        _2579_ = 8'b00011110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????? :
        _2579_ = 8'b01011010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????? :
        _2579_ = 8'b00101001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????? :
        _2579_ = 8'b10000010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????? :
        _2579_ = 8'b11010000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????? :
        _2579_ = 8'b10000100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????? :
        _2579_ = 8'b11010111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????? :
        _2579_ = 8'b01100101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????? :
        _2579_ = 8'b00011010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????? :
        _2579_ = 8'b00001001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????? :
        _2579_ = 8'b01011001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????? :
        _2579_ = 8'b00000011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????? :
        _2579_ = 8'b10100101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????? :
        _2579_ = 8'b01010000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????? :
        _2579_ = 8'b10101010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????? :
        _2579_ = 8'b10000111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????? :
        _2579_ = 8'b11001001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????? :
        _2579_ = 8'b00010101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????? :
        _2579_ = 8'b00111100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????? :
        _2579_ = 8'b00101101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????? :
        _2579_ = 8'b00110011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????? :
        _2579_ = 8'b00000111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????? :
        _2579_ = 8'b10101001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????? :
        _2579_ = 8'b11010010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????? :
        _2579_ = 8'b00100010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????? :
        _2579_ = 8'b00101011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????? :
        _2579_ = 8'b11101011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????? :
        _2579_ = 8'b11011001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????? :
        _2579_ = 8'b00100111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????? :
        _2579_ = 8'b00111010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????? :
        _2579_ = 8'b10011001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????? :
        _2579_ = 8'b00010111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????? :
        _2579_ = 8'b01101001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????? :
        _2579_ = 8'b10101110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????? :
        _2579_ = 8'b01101010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????? :
        _2579_ = 8'b11000010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????? :
        _2579_ = 8'b00011100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????? :
        _2579_ = 8'b11110111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????? :
        _2579_ = 8'b00000110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????? :
        _2579_ = 8'b10010000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????? :
        _2579_ = 8'b11001100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????? :
        _2579_ = 8'b01110001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????? :
        _2579_ = 8'b01111100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????? :
        _2579_ = 8'b11100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????? :
        _2579_ = 8'b00001111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????? :
        _2579_ = 8'b00001101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????? :
        _2579_ = 8'b01100001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????? :
        _2579_ = 8'b10010110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????? :
        _2579_ = 8'b00111110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????? :
        _2579_ = 8'b11101000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????? :
        _2579_ = 8'b10100001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????? :
        _2579_ = 8'b11001011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????? :
        _2579_ = 8'b10010111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????? :
        _2579_ = 8'b01110011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????? :
        _2579_ = 8'b01010111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????? :
        _2579_ = 8'b00111000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????? :
        _2579_ = 8'b01011100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????? :
        _2579_ = 8'b01001010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????? :
        _2579_ = 8'b11110000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????? :
        _2579_ = 8'b01101111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????? :
        _2579_ = 8'b00010000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b01000111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b11110100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b11001010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b11001111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b11110011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b10101100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b11011000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b01001001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b10011100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b10110001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b00000001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b11011010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b01101110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b10001011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b11010101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b11110010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b11010011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b00110001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b00111001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b11000100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b01000011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b10111101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b10011111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b10111000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b01001000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b00001100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b10010010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b00010100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b01110100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b01100100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b11011011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b10101101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b00010110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b10111100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b10100111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b00101000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b01101011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b11000111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b10001100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b00001011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b00111011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b01010100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b01000100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b10100011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b10011110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b00011001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b11000000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b11100110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b00110010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b10111010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b11001000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b01111010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b11111100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b01010101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b10010011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b00101110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b10001000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b00110101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b10111110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b11000011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b00100110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b00011000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b10000001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b10111111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b11111101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b11100101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b00100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b01000010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b10101111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b01110111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b01100011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b11110001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b01110000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b00100001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b00111111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b00000101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b10000000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b01011101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b10100010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b01001011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b00100101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b01111000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b10100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b11111110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b00000100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b11101001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b10001010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b00010001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b01100110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b10011010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b10000110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b11101101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b01001111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b11000101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b10111011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b10000101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b10110000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b10011000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b10010100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b01110010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b01100111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b10001101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b11010100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b10110110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b01111001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b11100011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b01000000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b11000001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b00000000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b10111001 ;
      256'b????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b10100110 ;
      256'b???????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b00010011 ;
      256'b??????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b01011110 ;
      256'b?????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b11011101 ;
      256'b????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b01010010 ;
      256'b???????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b01111101 ;
      256'b??????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b10110111 ;
      256'b?????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b01110110 ;
      256'b????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b10100100 ;
      256'b???????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b01011011 ;
      256'b??????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b10110100 ;
      256'b?????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b11011100 ;
      256'b????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b00110110 ;
      256'b???????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b00110100 ;
      256'b??????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b01011000 ;
      256'b?????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b00011101 ;
      256'b????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b00010010 ;
      256'b???????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b11101010 ;
      256'b??????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b01111111 ;
      256'b?????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b01001110 ;
      256'b????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b11001101 ;
      256'b???????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b11011111 ;
      256'b??????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b00011011 ;
      256'b?????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b00100100 ;
      256'b????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b00001110 ;
      256'b???????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b00101111 ;
      256'b??????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b00001010 ;
      256'b?????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b00110111 ;
      256'b????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b00110000 ;
      256'b???????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b10011101 ;
      256'b??????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b01000110 ;
      256'b?????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b10010101 ;
      256'b????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b00001000 ;
      256'b???????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b00101010 ;
      256'b??????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b01100010 ;
      256'b?????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b10101011 ;
      256'b????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b11100010 ;
      256'b???????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b11111001 ;
      256'b??????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b11010001 ;
      256'b?????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b01010001 ;
      256'b????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b01101000 ;
      256'b???????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b10000011 ;
      256'b??????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b11110101 ;
      256'b?????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b01111110 ;
      256'b????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b01101100 ;
      256'b???????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b01001100 ;
      256'b??????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b00111101 ;
      256'b?????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b11100001 ;
      256'b????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b01110101 ;
      256'b???????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b10011011 ;
      256'b??????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b11100100 ;
      256'b?????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b01010011 ;
      256'b????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b00100011 ;
      256'b???????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b01000101 ;
      256'b??????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b01011111 ;
      256'b?????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b10110011 ;
      256'b????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b01000001 ;
      256'b???????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b11111011 ;
      256'b??????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b10001110 ;
      256'b?????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b10110010 ;
      256'b????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b11101111 ;
      256'b???????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b11111010 ;
      256'b??????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b10001001 ;
      256'b?????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b00011111 ;
      256'b????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b10001111 ;
      256'b???????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b11101100 ;
      256'b??????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b01001101 ;
      256'b?????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b10110101 ;
      256'b????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b11100111 ;
      256'b???????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b01010110 ;
      256'b??????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b11001110 ;
      256'b?????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b00000010 ;
      256'b????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b01100000 ;
      256'b???????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b10010001 ;
      256'b??????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b11011110 ;
      256'b?????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b11010110 ;
      256'b????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b11111111 ;
      256'b???1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b11110110 ;
      256'b??1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b11101110 ;
      256'b?1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b11111000 ;
      256'b1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b11000110 ;
      default:
        _2579_ = \t2.t1.s4.out ;
    endcase
  end
  assign p22[23:16] = \t2.t2.s0.out ^ \t2.t2.s4.out ;
  always @(posedge clk)
      \t2.t2.s0.out <= _2580_;
  wire [255:0] fangyuan21;
  assign fangyuan21 = { _2836_, _2835_, _2834_, _2833_, _2832_, _2831_, _2830_, _2829_, _2828_, _2827_, _2826_, _2825_, _2824_, _2823_, _2822_, _2821_, _2820_, _2819_, _2818_, _2817_, _2816_, _2815_, _2814_, _2813_, _2812_, _2811_, _2810_, _2809_, _2808_, _2807_, _2806_, _2805_, _2804_, _2803_, _2802_, _2801_, _2800_, _2799_, _2798_, _2797_, _2796_, _2795_, _2794_, _2793_, _2792_, _2791_, _2790_, _2789_, _2788_, _2787_, _2786_, _2785_, _2784_, _2783_, _2782_, _2781_, _2780_, _2779_, _2778_, _2777_, _2776_, _2775_, _2774_, _2773_, _2772_, _2771_, _2770_, _2769_, _2768_, _2767_, _2766_, _2765_, _2764_, _2763_, _2762_, _2761_, _2760_, _2759_, _2758_, _2757_, _2756_, _2755_, _2754_, _2753_, _2752_, _2751_, _2750_, _2749_, _2748_, _2747_, _2746_, _2745_, _2744_, _2743_, _2742_, _2741_, _2740_, _2739_, _2738_, _2737_, _2736_, _2735_, _2734_, _2733_, _2732_, _2731_, _2730_, _2729_, _2728_, _2727_, _2726_, _2725_, _2724_, _2723_, _2722_, _2721_, _2720_, _2719_, _2718_, _2717_, _2716_, _2715_, _2714_, _2713_, _2712_, _2711_, _2710_, _2709_, _2708_, _2707_, _2706_, _2705_, _2704_, _2703_, _2702_, _2701_, _2700_, _2699_, _2698_, _2697_, _2696_, _2695_, _2694_, _2693_, _2692_, _2691_, _2690_, _2689_, _2688_, _2687_, _2686_, _2685_, _2684_, _2683_, _2682_, _2681_, _2680_, _2679_, _2678_, _2677_, _2676_, _2675_, _2674_, _2673_, _2672_, _2671_, _2670_, _2669_, _2668_, _2667_, _2666_, _2665_, _2664_, _2663_, _2662_, _2661_, _2660_, _2659_, _2658_, _2657_, _2656_, _2655_, _2654_, _2653_, _2652_, _2651_, _2650_, _2649_, _2648_, _2647_, _2646_, _2645_, _2644_, _2643_, _2642_, _2641_, _2640_, _2639_, _2638_, _2637_, _2636_, _2635_, _2634_, _2633_, _2632_, _2631_, _2630_, _2629_, _2628_, _2627_, _2626_, _2625_, _2624_, _2623_, _2622_, _2621_, _2620_, _2619_, _2618_, _2617_, _2616_, _2615_, _2614_, _2613_, _2612_, _2611_, _2610_, _2609_, _2608_, _2607_, _2606_, _2605_, _2604_, _2603_, _2602_, _2601_, _2600_, _2599_, _2598_, _2597_, _2596_, _2595_, _2594_, _2593_, _2592_, _2591_, _2590_, _2589_, _2588_, _2587_, _2586_, _2585_, _2584_, _2583_, _2582_, _2581_ };

  always @(\t2.t2.s0.out or fangyuan21) begin
    casez (fangyuan21)
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1 :
        _2580_ = 8'b00010110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1? :
        _2580_ = 8'b10111011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?? :
        _2580_ = 8'b01010100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??? :
        _2580_ = 8'b10110000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???? :
        _2580_ = 8'b00001111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????? :
        _2580_ = 8'b00101101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????? :
        _2580_ = 8'b10011001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????? :
        _2580_ = 8'b01000001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????? :
        _2580_ = 8'b01101000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????? :
        _2580_ = 8'b01000010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????? :
        _2580_ = 8'b11100110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????? :
        _2580_ = 8'b10111111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????? :
        _2580_ = 8'b00001101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????? :
        _2580_ = 8'b10001001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????? :
        _2580_ = 8'b10100001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????? :
        _2580_ = 8'b10001100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????? :
        _2580_ = 8'b11011111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????? :
        _2580_ = 8'b00101000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????? :
        _2580_ = 8'b01010101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????? :
        _2580_ = 8'b11001110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????? :
        _2580_ = 8'b11101001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????? :
        _2580_ = 8'b10000111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????? :
        _2580_ = 8'b00011110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????? :
        _2580_ = 8'b10011011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????? :
        _2580_ = 8'b10010100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????? :
        _2580_ = 8'b10001110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????? :
        _2580_ = 8'b11011001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????? :
        _2580_ = 8'b01101001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????? :
        _2580_ = 8'b00010001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????? :
        _2580_ = 8'b10011000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????? :
        _2580_ = 8'b11111000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????? :
        _2580_ = 8'b11100001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????? :
        _2580_ = 8'b10011110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????? :
        _2580_ = 8'b00011101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????? :
        _2580_ = 8'b11000001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????? :
        _2580_ = 8'b10000110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????? :
        _2580_ = 8'b10111001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????? :
        _2580_ = 8'b01010111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????? :
        _2580_ = 8'b00110101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????? :
        _2580_ = 8'b01100001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????? :
        _2580_ = 8'b00001110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????? :
        _2580_ = 8'b11110110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????? :
        _2580_ = 8'b00000011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????? :
        _2580_ = 8'b01001000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????? :
        _2580_ = 8'b01100110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????? :
        _2580_ = 8'b10110101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????? :
        _2580_ = 8'b00111110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????? :
        _2580_ = 8'b01110000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????? :
        _2580_ = 8'b10001010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????? :
        _2580_ = 8'b10001011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????? :
        _2580_ = 8'b10111101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????? :
        _2580_ = 8'b01001011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????? :
        _2580_ = 8'b00011111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????? :
        _2580_ = 8'b01110100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????? :
        _2580_ = 8'b11011101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????? :
        _2580_ = 8'b11101000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????? :
        _2580_ = 8'b11000110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????? :
        _2580_ = 8'b10110100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????? :
        _2580_ = 8'b10100110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????? :
        _2580_ = 8'b00011100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????? :
        _2580_ = 8'b00101110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????? :
        _2580_ = 8'b00100101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????? :
        _2580_ = 8'b01111000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????? :
        _2580_ = 8'b10111010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????? :
        _2580_ = 8'b00001000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b10101110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b01111010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b01100101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b11101010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b11110100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b01010110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b01101100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b10101001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b01001110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b11010101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b10001101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b01101101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b00110111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b11001000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b11100111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b01111001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b11100100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b10010101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b10010001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b01100010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b10101100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b11010011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b11000010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b01011100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b00100100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b00000110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b01001001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b00001010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b00111010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b00110010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b11100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b11011011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b00001011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b01011110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b11011110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b00010100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b10111000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b11101110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b01000110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b10001000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b10010000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b00101010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b00100010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b11011100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b01001111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b10000001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b01100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b01110011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b00011001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b01011101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b01100100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b00111101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b01111110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b10100111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b11000100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b00010111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b01000100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b10010111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b01011111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b11101100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b00010011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b00001100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b11001101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b11010010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b11110011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b11111111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b00010000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b00100001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b11011010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b10110110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b10111100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b11110101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b00111000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b10011101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b10010010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b10001111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b01000000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b10100011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b01010001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b10101000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b10011111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b00111100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b01010000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b01111111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b00000010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b11111001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b01000101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b10000101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b00110011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b01001101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b01000011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b11111011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b10101010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b11101111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b11010000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b11001111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b01011000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b01001100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b01001010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b00111001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b10111110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b11001011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b01101010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b01011011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b10110001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b11111100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b00100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b11101101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b00000000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b11010001 ;
      256'b????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b01010011 ;
      256'b???????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b10000100 ;
      256'b??????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b00101111 ;
      256'b?????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b11100011 ;
      256'b????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b00101001 ;
      256'b???????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b10110011 ;
      256'b??????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b11010110 ;
      256'b?????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b00111011 ;
      256'b????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b01010010 ;
      256'b???????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b10100000 ;
      256'b??????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b01011010 ;
      256'b?????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b01101110 ;
      256'b????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b00011011 ;
      256'b???????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b00011010 ;
      256'b??????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b00101100 ;
      256'b?????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b10000011 ;
      256'b????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b00001001 ;
      256'b???????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b01110101 ;
      256'b??????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b10110010 ;
      256'b?????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b00100111 ;
      256'b????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b11101011 ;
      256'b???????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b11100010 ;
      256'b??????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b10000000 ;
      256'b?????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b00010010 ;
      256'b????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b00000111 ;
      256'b???????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b10011010 ;
      256'b??????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b00000101 ;
      256'b?????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b10010110 ;
      256'b????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b00011000 ;
      256'b???????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b11000011 ;
      256'b??????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b00100011 ;
      256'b?????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b11000111 ;
      256'b????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b00000100 ;
      256'b???????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b00010101 ;
      256'b??????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b00110001 ;
      256'b?????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b11011000 ;
      256'b????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b01110001 ;
      256'b???????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b11110001 ;
      256'b??????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b11100101 ;
      256'b?????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b10100101 ;
      256'b????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b00110100 ;
      256'b???????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b11001100 ;
      256'b??????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b11110111 ;
      256'b?????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b00111111 ;
      256'b????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b00110110 ;
      256'b???????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b00100110 ;
      256'b??????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b10010011 ;
      256'b?????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b11111101 ;
      256'b????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b10110111 ;
      256'b???????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b11000000 ;
      256'b??????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b01110010 ;
      256'b?????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b10100100 ;
      256'b????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b10011100 ;
      256'b???????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b10101111 ;
      256'b??????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b10100010 ;
      256'b?????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b11010100 ;
      256'b????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b10101101 ;
      256'b???????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b11110000 ;
      256'b??????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b01000111 ;
      256'b?????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b01011001 ;
      256'b????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b11111010 ;
      256'b???????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b01111101 ;
      256'b??????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b11001001 ;
      256'b?????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b10000010 ;
      256'b????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b11001010 ;
      256'b???????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b01110110 ;
      256'b??????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b10101011 ;
      256'b?????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b11010111 ;
      256'b????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b11111110 ;
      256'b???????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b00101011 ;
      256'b??????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b01100111 ;
      256'b?????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b00000001 ;
      256'b????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b00110000 ;
      256'b???????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b11000101 ;
      256'b??????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b01101111 ;
      256'b?????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b01101011 ;
      256'b????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b11110010 ;
      256'b???1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b01111011 ;
      256'b??1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b01110111 ;
      256'b?1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b01111100 ;
      256'b1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b01100011 ;
      default:
        _2580_ = \t2.t2.s0.out ;
    endcase
  end
  assign _2581_ = state_in[47:40] == 8'b11111111;
  assign _2582_ = state_in[47:40] == 8'b11111110;
  assign _2583_ = state_in[47:40] == 8'b11111101;
  assign _2584_ = state_in[47:40] == 8'b11111100;
  assign _2585_ = state_in[47:40] == 8'b11111011;
  assign _2586_ = state_in[47:40] == 8'b11111010;
  assign _2587_ = state_in[47:40] == 8'b11111001;
  assign _2588_ = state_in[47:40] == 8'b11111000;
  assign _2589_ = state_in[47:40] == 8'b11110111;
  assign _2590_ = state_in[47:40] == 8'b11110110;
  assign _2591_ = state_in[47:40] == 8'b11110101;
  assign _2592_ = state_in[47:40] == 8'b11110100;
  assign _2593_ = state_in[47:40] == 8'b11110011;
  assign _2594_ = state_in[47:40] == 8'b11110010;
  assign _2595_ = state_in[47:40] == 8'b11110001;
  assign _2596_ = state_in[47:40] == 8'b11110000;
  assign _2597_ = state_in[47:40] == 8'b11101111;
  assign _2598_ = state_in[47:40] == 8'b11101110;
  assign _2599_ = state_in[47:40] == 8'b11101101;
  assign _2600_ = state_in[47:40] == 8'b11101100;
  assign _2601_ = state_in[47:40] == 8'b11101011;
  assign _2602_ = state_in[47:40] == 8'b11101010;
  assign _2603_ = state_in[47:40] == 8'b11101001;
  assign _2604_ = state_in[47:40] == 8'b11101000;
  assign _2605_ = state_in[47:40] == 8'b11100111;
  assign _2606_ = state_in[47:40] == 8'b11100110;
  assign _2607_ = state_in[47:40] == 8'b11100101;
  assign _2608_ = state_in[47:40] == 8'b11100100;
  assign _2609_ = state_in[47:40] == 8'b11100011;
  assign _2610_ = state_in[47:40] == 8'b11100010;
  assign _2611_ = state_in[47:40] == 8'b11100001;
  assign _2612_ = state_in[47:40] == 8'b11100000;
  assign _2613_ = state_in[47:40] == 8'b11011111;
  assign _2614_ = state_in[47:40] == 8'b11011110;
  assign _2615_ = state_in[47:40] == 8'b11011101;
  assign _2616_ = state_in[47:40] == 8'b11011100;
  assign _2617_ = state_in[47:40] == 8'b11011011;
  assign _2618_ = state_in[47:40] == 8'b11011010;
  assign _2619_ = state_in[47:40] == 8'b11011001;
  assign _2620_ = state_in[47:40] == 8'b11011000;
  assign _2621_ = state_in[47:40] == 8'b11010111;
  assign _2622_ = state_in[47:40] == 8'b11010110;
  assign _2623_ = state_in[47:40] == 8'b11010101;
  assign _2624_ = state_in[47:40] == 8'b11010100;
  assign _2625_ = state_in[47:40] == 8'b11010011;
  assign _2626_ = state_in[47:40] == 8'b11010010;
  assign _2627_ = state_in[47:40] == 8'b11010001;
  assign _2628_ = state_in[47:40] == 8'b11010000;
  assign _2629_ = state_in[47:40] == 8'b11001111;
  assign _2630_ = state_in[47:40] == 8'b11001110;
  assign _2631_ = state_in[47:40] == 8'b11001101;
  assign _2632_ = state_in[47:40] == 8'b11001100;
  assign _2633_ = state_in[47:40] == 8'b11001011;
  assign _2634_ = state_in[47:40] == 8'b11001010;
  assign _2635_ = state_in[47:40] == 8'b11001001;
  assign _2636_ = state_in[47:40] == 8'b11001000;
  assign _2637_ = state_in[47:40] == 8'b11000111;
  assign _2638_ = state_in[47:40] == 8'b11000110;
  assign _2639_ = state_in[47:40] == 8'b11000101;
  assign _2640_ = state_in[47:40] == 8'b11000100;
  assign _2641_ = state_in[47:40] == 8'b11000011;
  assign _2642_ = state_in[47:40] == 8'b11000010;
  assign _2643_ = state_in[47:40] == 8'b11000001;
  assign _2644_ = state_in[47:40] == 8'b11000000;
  assign _2645_ = state_in[47:40] == 8'b10111111;
  assign _2646_ = state_in[47:40] == 8'b10111110;
  assign _2647_ = state_in[47:40] == 8'b10111101;
  assign _2648_ = state_in[47:40] == 8'b10111100;
  assign _2649_ = state_in[47:40] == 8'b10111011;
  assign _2650_ = state_in[47:40] == 8'b10111010;
  assign _2651_ = state_in[47:40] == 8'b10111001;
  assign _2652_ = state_in[47:40] == 8'b10111000;
  assign _2653_ = state_in[47:40] == 8'b10110111;
  assign _2654_ = state_in[47:40] == 8'b10110110;
  assign _2655_ = state_in[47:40] == 8'b10110101;
  assign _2656_ = state_in[47:40] == 8'b10110100;
  assign _2657_ = state_in[47:40] == 8'b10110011;
  assign _2658_ = state_in[47:40] == 8'b10110010;
  assign _2659_ = state_in[47:40] == 8'b10110001;
  assign _2660_ = state_in[47:40] == 8'b10110000;
  assign _2661_ = state_in[47:40] == 8'b10101111;
  assign _2662_ = state_in[47:40] == 8'b10101110;
  assign _2663_ = state_in[47:40] == 8'b10101101;
  assign _2664_ = state_in[47:40] == 8'b10101100;
  assign _2665_ = state_in[47:40] == 8'b10101011;
  assign _2666_ = state_in[47:40] == 8'b10101010;
  assign _2667_ = state_in[47:40] == 8'b10101001;
  assign _2668_ = state_in[47:40] == 8'b10101000;
  assign _2669_ = state_in[47:40] == 8'b10100111;
  assign _2670_ = state_in[47:40] == 8'b10100110;
  assign _2671_ = state_in[47:40] == 8'b10100101;
  assign _2672_ = state_in[47:40] == 8'b10100100;
  assign _2673_ = state_in[47:40] == 8'b10100011;
  assign _2674_ = state_in[47:40] == 8'b10100010;
  assign _2675_ = state_in[47:40] == 8'b10100001;
  assign _2676_ = state_in[47:40] == 8'b10100000;
  assign _2677_ = state_in[47:40] == 8'b10011111;
  assign _2678_ = state_in[47:40] == 8'b10011110;
  assign _2679_ = state_in[47:40] == 8'b10011101;
  assign _2680_ = state_in[47:40] == 8'b10011100;
  assign _2681_ = state_in[47:40] == 8'b10011011;
  assign _2682_ = state_in[47:40] == 8'b10011010;
  assign _2683_ = state_in[47:40] == 8'b10011001;
  assign _2684_ = state_in[47:40] == 8'b10011000;
  assign _2685_ = state_in[47:40] == 8'b10010111;
  assign _2686_ = state_in[47:40] == 8'b10010110;
  assign _2687_ = state_in[47:40] == 8'b10010101;
  assign _2688_ = state_in[47:40] == 8'b10010100;
  assign _2689_ = state_in[47:40] == 8'b10010011;
  assign _2690_ = state_in[47:40] == 8'b10010010;
  assign _2691_ = state_in[47:40] == 8'b10010001;
  assign _2692_ = state_in[47:40] == 8'b10010000;
  assign _2693_ = state_in[47:40] == 8'b10001111;
  assign _2694_ = state_in[47:40] == 8'b10001110;
  assign _2695_ = state_in[47:40] == 8'b10001101;
  assign _2696_ = state_in[47:40] == 8'b10001100;
  assign _2697_ = state_in[47:40] == 8'b10001011;
  assign _2698_ = state_in[47:40] == 8'b10001010;
  assign _2699_ = state_in[47:40] == 8'b10001001;
  assign _2700_ = state_in[47:40] == 8'b10001000;
  assign _2701_ = state_in[47:40] == 8'b10000111;
  assign _2702_ = state_in[47:40] == 8'b10000110;
  assign _2703_ = state_in[47:40] == 8'b10000101;
  assign _2704_ = state_in[47:40] == 8'b10000100;
  assign _2705_ = state_in[47:40] == 8'b10000011;
  assign _2706_ = state_in[47:40] == 8'b10000010;
  assign _2707_ = state_in[47:40] == 8'b10000001;
  assign _2708_ = state_in[47:40] == 8'b10000000;
  assign _2709_ = state_in[47:40] == 7'b1111111;
  assign _2710_ = state_in[47:40] == 7'b1111110;
  assign _2711_ = state_in[47:40] == 7'b1111101;
  assign _2712_ = state_in[47:40] == 7'b1111100;
  assign _2713_ = state_in[47:40] == 7'b1111011;
  assign _2714_ = state_in[47:40] == 7'b1111010;
  assign _2715_ = state_in[47:40] == 7'b1111001;
  assign _2716_ = state_in[47:40] == 7'b1111000;
  assign _2717_ = state_in[47:40] == 7'b1110111;
  assign _2718_ = state_in[47:40] == 7'b1110110;
  assign _2719_ = state_in[47:40] == 7'b1110101;
  assign _2720_ = state_in[47:40] == 7'b1110100;
  assign _2721_ = state_in[47:40] == 7'b1110011;
  assign _2722_ = state_in[47:40] == 7'b1110010;
  assign _2723_ = state_in[47:40] == 7'b1110001;
  assign _2724_ = state_in[47:40] == 7'b1110000;
  assign _2725_ = state_in[47:40] == 7'b1101111;
  assign _2726_ = state_in[47:40] == 7'b1101110;
  assign _2727_ = state_in[47:40] == 7'b1101101;
  assign _2728_ = state_in[47:40] == 7'b1101100;
  assign _2729_ = state_in[47:40] == 7'b1101011;
  assign _2730_ = state_in[47:40] == 7'b1101010;
  assign _2731_ = state_in[47:40] == 7'b1101001;
  assign _2732_ = state_in[47:40] == 7'b1101000;
  assign _2733_ = state_in[47:40] == 7'b1100111;
  assign _2734_ = state_in[47:40] == 7'b1100110;
  assign _2735_ = state_in[47:40] == 7'b1100101;
  assign _2736_ = state_in[47:40] == 7'b1100100;
  assign _2737_ = state_in[47:40] == 7'b1100011;
  assign _2738_ = state_in[47:40] == 7'b1100010;
  assign _2739_ = state_in[47:40] == 7'b1100001;
  assign _2740_ = state_in[47:40] == 7'b1100000;
  assign _2741_ = state_in[47:40] == 7'b1011111;
  assign _2742_ = state_in[47:40] == 7'b1011110;
  assign _2743_ = state_in[47:40] == 7'b1011101;
  assign _2744_ = state_in[47:40] == 7'b1011100;
  assign _2745_ = state_in[47:40] == 7'b1011011;
  assign _2746_ = state_in[47:40] == 7'b1011010;
  assign _2747_ = state_in[47:40] == 7'b1011001;
  assign _2748_ = state_in[47:40] == 7'b1011000;
  assign _2749_ = state_in[47:40] == 7'b1010111;
  assign _2750_ = state_in[47:40] == 7'b1010110;
  assign _2751_ = state_in[47:40] == 7'b1010101;
  assign _2752_ = state_in[47:40] == 7'b1010100;
  assign _2753_ = state_in[47:40] == 7'b1010011;
  assign _2754_ = state_in[47:40] == 7'b1010010;
  assign _2755_ = state_in[47:40] == 7'b1010001;
  assign _2756_ = state_in[47:40] == 7'b1010000;
  assign _2757_ = state_in[47:40] == 7'b1001111;
  assign _2758_ = state_in[47:40] == 7'b1001110;
  assign _2759_ = state_in[47:40] == 7'b1001101;
  assign _2760_ = state_in[47:40] == 7'b1001100;
  assign _2761_ = state_in[47:40] == 7'b1001011;
  assign _2762_ = state_in[47:40] == 7'b1001010;
  assign _2763_ = state_in[47:40] == 7'b1001001;
  assign _2764_ = state_in[47:40] == 7'b1001000;
  assign _2765_ = state_in[47:40] == 7'b1000111;
  assign _2766_ = state_in[47:40] == 7'b1000110;
  assign _2767_ = state_in[47:40] == 7'b1000101;
  assign _2768_ = state_in[47:40] == 7'b1000100;
  assign _2769_ = state_in[47:40] == 7'b1000011;
  assign _2770_ = state_in[47:40] == 7'b1000010;
  assign _2771_ = state_in[47:40] == 7'b1000001;
  assign _2772_ = state_in[47:40] == 7'b1000000;
  assign _2773_ = state_in[47:40] == 6'b111111;
  assign _2774_ = state_in[47:40] == 6'b111110;
  assign _2775_ = state_in[47:40] == 6'b111101;
  assign _2776_ = state_in[47:40] == 6'b111100;
  assign _2777_ = state_in[47:40] == 6'b111011;
  assign _2778_ = state_in[47:40] == 6'b111010;
  assign _2779_ = state_in[47:40] == 6'b111001;
  assign _2780_ = state_in[47:40] == 6'b111000;
  assign _2781_ = state_in[47:40] == 6'b110111;
  assign _2782_ = state_in[47:40] == 6'b110110;
  assign _2783_ = state_in[47:40] == 6'b110101;
  assign _2784_ = state_in[47:40] == 6'b110100;
  assign _2785_ = state_in[47:40] == 6'b110011;
  assign _2786_ = state_in[47:40] == 6'b110010;
  assign _2787_ = state_in[47:40] == 6'b110001;
  assign _2788_ = state_in[47:40] == 6'b110000;
  assign _2789_ = state_in[47:40] == 6'b101111;
  assign _2790_ = state_in[47:40] == 6'b101110;
  assign _2791_ = state_in[47:40] == 6'b101101;
  assign _2792_ = state_in[47:40] == 6'b101100;
  assign _2793_ = state_in[47:40] == 6'b101011;
  assign _2794_ = state_in[47:40] == 6'b101010;
  assign _2795_ = state_in[47:40] == 6'b101001;
  assign _2796_ = state_in[47:40] == 6'b101000;
  assign _2797_ = state_in[47:40] == 6'b100111;
  assign _2798_ = state_in[47:40] == 6'b100110;
  assign _2799_ = state_in[47:40] == 6'b100101;
  assign _2800_ = state_in[47:40] == 6'b100100;
  assign _2801_ = state_in[47:40] == 6'b100011;
  assign _2802_ = state_in[47:40] == 6'b100010;
  assign _2803_ = state_in[47:40] == 6'b100001;
  assign _2804_ = state_in[47:40] == 6'b100000;
  assign _2805_ = state_in[47:40] == 5'b11111;
  assign _2806_ = state_in[47:40] == 5'b11110;
  assign _2807_ = state_in[47:40] == 5'b11101;
  assign _2808_ = state_in[47:40] == 5'b11100;
  assign _2809_ = state_in[47:40] == 5'b11011;
  assign _2810_ = state_in[47:40] == 5'b11010;
  assign _2811_ = state_in[47:40] == 5'b11001;
  assign _2812_ = state_in[47:40] == 5'b11000;
  assign _2813_ = state_in[47:40] == 5'b10111;
  assign _2814_ = state_in[47:40] == 5'b10110;
  assign _2815_ = state_in[47:40] == 5'b10101;
  assign _2816_ = state_in[47:40] == 5'b10100;
  assign _2817_ = state_in[47:40] == 5'b10011;
  assign _2818_ = state_in[47:40] == 5'b10010;
  assign _2819_ = state_in[47:40] == 5'b10001;
  assign _2820_ = state_in[47:40] == 5'b10000;
  assign _2821_ = state_in[47:40] == 4'b1111;
  assign _2822_ = state_in[47:40] == 4'b1110;
  assign _2823_ = state_in[47:40] == 4'b1101;
  assign _2824_ = state_in[47:40] == 4'b1100;
  assign _2825_ = state_in[47:40] == 4'b1011;
  assign _2826_ = state_in[47:40] == 4'b1010;
  assign _2827_ = state_in[47:40] == 4'b1001;
  assign _2828_ = state_in[47:40] == 4'b1000;
  assign _2829_ = state_in[47:40] == 3'b111;
  assign _2830_ = state_in[47:40] == 3'b110;
  assign _2831_ = state_in[47:40] == 3'b101;
  assign _2832_ = state_in[47:40] == 3'b100;
  assign _2833_ = state_in[47:40] == 2'b11;
  assign _2834_ = state_in[47:40] == 2'b10;
  assign _2835_ = state_in[47:40] == 1'b1;
  assign _2836_ = ! state_in[47:40];
  always @(posedge clk)
      \t2.t2.s4.out <= _2837_;
  wire [255:0] fangyuan22;
  assign fangyuan22 = { _2836_, _2835_, _2834_, _2833_, _2832_, _2831_, _2830_, _2829_, _2828_, _2827_, _2826_, _2825_, _2824_, _2823_, _2822_, _2821_, _2820_, _2819_, _2818_, _2817_, _2816_, _2815_, _2814_, _2813_, _2812_, _2811_, _2810_, _2809_, _2808_, _2807_, _2806_, _2805_, _2804_, _2803_, _2802_, _2801_, _2800_, _2799_, _2798_, _2797_, _2796_, _2795_, _2794_, _2793_, _2792_, _2791_, _2790_, _2789_, _2788_, _2787_, _2786_, _2785_, _2784_, _2783_, _2782_, _2781_, _2780_, _2779_, _2778_, _2777_, _2776_, _2775_, _2774_, _2773_, _2772_, _2771_, _2770_, _2769_, _2768_, _2767_, _2766_, _2765_, _2764_, _2763_, _2762_, _2761_, _2760_, _2759_, _2758_, _2757_, _2756_, _2755_, _2754_, _2753_, _2752_, _2751_, _2750_, _2749_, _2748_, _2747_, _2746_, _2745_, _2744_, _2743_, _2742_, _2741_, _2740_, _2739_, _2738_, _2737_, _2736_, _2735_, _2734_, _2733_, _2732_, _2731_, _2730_, _2729_, _2728_, _2727_, _2726_, _2725_, _2724_, _2723_, _2722_, _2721_, _2720_, _2719_, _2718_, _2717_, _2716_, _2715_, _2714_, _2713_, _2712_, _2711_, _2710_, _2709_, _2708_, _2707_, _2706_, _2705_, _2704_, _2703_, _2702_, _2701_, _2700_, _2699_, _2698_, _2697_, _2696_, _2695_, _2694_, _2693_, _2692_, _2691_, _2690_, _2689_, _2688_, _2687_, _2686_, _2685_, _2684_, _2683_, _2682_, _2681_, _2680_, _2679_, _2678_, _2677_, _2676_, _2675_, _2674_, _2673_, _2672_, _2671_, _2670_, _2669_, _2668_, _2667_, _2666_, _2665_, _2664_, _2663_, _2662_, _2661_, _2660_, _2659_, _2658_, _2657_, _2656_, _2655_, _2654_, _2653_, _2652_, _2651_, _2650_, _2649_, _2648_, _2647_, _2646_, _2645_, _2644_, _2643_, _2642_, _2641_, _2640_, _2639_, _2638_, _2637_, _2636_, _2635_, _2634_, _2633_, _2632_, _2631_, _2630_, _2629_, _2628_, _2627_, _2626_, _2625_, _2624_, _2623_, _2622_, _2621_, _2620_, _2619_, _2618_, _2617_, _2616_, _2615_, _2614_, _2613_, _2612_, _2611_, _2610_, _2609_, _2608_, _2607_, _2606_, _2605_, _2604_, _2603_, _2602_, _2601_, _2600_, _2599_, _2598_, _2597_, _2596_, _2595_, _2594_, _2593_, _2592_, _2591_, _2590_, _2589_, _2588_, _2587_, _2586_, _2585_, _2584_, _2583_, _2582_, _2581_ };

  always @(\t2.t2.s4.out or fangyuan22) begin
    casez (fangyuan22)
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1 :
        _2837_ = 8'b00101100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1? :
        _2837_ = 8'b01101101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?? :
        _2837_ = 8'b10101000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??? :
        _2837_ = 8'b01111011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???? :
        _2837_ = 8'b00011110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????? :
        _2837_ = 8'b01011010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????? :
        _2837_ = 8'b00101001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????? :
        _2837_ = 8'b10000010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????? :
        _2837_ = 8'b11010000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????? :
        _2837_ = 8'b10000100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????? :
        _2837_ = 8'b11010111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????? :
        _2837_ = 8'b01100101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????? :
        _2837_ = 8'b00011010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????? :
        _2837_ = 8'b00001001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????? :
        _2837_ = 8'b01011001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????? :
        _2837_ = 8'b00000011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????? :
        _2837_ = 8'b10100101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????? :
        _2837_ = 8'b01010000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????? :
        _2837_ = 8'b10101010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????? :
        _2837_ = 8'b10000111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????? :
        _2837_ = 8'b11001001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????? :
        _2837_ = 8'b00010101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????? :
        _2837_ = 8'b00111100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????? :
        _2837_ = 8'b00101101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????? :
        _2837_ = 8'b00110011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????? :
        _2837_ = 8'b00000111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????? :
        _2837_ = 8'b10101001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????? :
        _2837_ = 8'b11010010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????? :
        _2837_ = 8'b00100010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????? :
        _2837_ = 8'b00101011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????? :
        _2837_ = 8'b11101011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????? :
        _2837_ = 8'b11011001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????? :
        _2837_ = 8'b00100111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????? :
        _2837_ = 8'b00111010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????? :
        _2837_ = 8'b10011001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????? :
        _2837_ = 8'b00010111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????? :
        _2837_ = 8'b01101001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????? :
        _2837_ = 8'b10101110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????? :
        _2837_ = 8'b01101010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????? :
        _2837_ = 8'b11000010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????? :
        _2837_ = 8'b00011100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????? :
        _2837_ = 8'b11110111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????? :
        _2837_ = 8'b00000110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????? :
        _2837_ = 8'b10010000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????? :
        _2837_ = 8'b11001100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????? :
        _2837_ = 8'b01110001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????? :
        _2837_ = 8'b01111100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????? :
        _2837_ = 8'b11100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????? :
        _2837_ = 8'b00001111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????? :
        _2837_ = 8'b00001101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????? :
        _2837_ = 8'b01100001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????? :
        _2837_ = 8'b10010110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????? :
        _2837_ = 8'b00111110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????? :
        _2837_ = 8'b11101000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????? :
        _2837_ = 8'b10100001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????? :
        _2837_ = 8'b11001011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????? :
        _2837_ = 8'b10010111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????? :
        _2837_ = 8'b01110011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????? :
        _2837_ = 8'b01010111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????? :
        _2837_ = 8'b00111000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????? :
        _2837_ = 8'b01011100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????? :
        _2837_ = 8'b01001010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????? :
        _2837_ = 8'b11110000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????? :
        _2837_ = 8'b01101111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????? :
        _2837_ = 8'b00010000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b01000111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b11110100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b11001010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b11001111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b11110011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b10101100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b11011000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b01001001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b10011100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b10110001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b00000001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b11011010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b01101110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b10001011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b11010101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b11110010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b11010011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b00110001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b00111001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b11000100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b01000011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b10111101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b10011111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b10111000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b01001000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b00001100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b10010010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b00010100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b01110100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b01100100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b11011011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b10101101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b00010110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b10111100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b10100111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b00101000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b01101011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b11000111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b10001100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b00001011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b00111011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b01010100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b01000100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b10100011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b10011110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b00011001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b11000000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b11100110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b00110010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b10111010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b11001000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b01111010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b11111100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b01010101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b10010011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b00101110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b10001000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b00110101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b10111110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b11000011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b00100110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b00011000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b10000001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b10111111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b11111101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b11100101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b00100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b01000010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b10101111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b01110111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b01100011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b11110001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b01110000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b00100001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b00111111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b00000101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b10000000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b01011101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b10100010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b01001011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b00100101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b01111000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b10100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b11111110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b00000100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b11101001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b10001010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b00010001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b01100110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b10011010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b10000110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b11101101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b01001111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b11000101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b10111011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b10000101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b10110000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b10011000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b10010100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b01110010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b01100111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b10001101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b11010100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b10110110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b01111001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b11100011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b01000000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b11000001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b00000000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b10111001 ;
      256'b????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b10100110 ;
      256'b???????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b00010011 ;
      256'b??????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b01011110 ;
      256'b?????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b11011101 ;
      256'b????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b01010010 ;
      256'b???????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b01111101 ;
      256'b??????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b10110111 ;
      256'b?????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b01110110 ;
      256'b????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b10100100 ;
      256'b???????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b01011011 ;
      256'b??????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b10110100 ;
      256'b?????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b11011100 ;
      256'b????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b00110110 ;
      256'b???????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b00110100 ;
      256'b??????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b01011000 ;
      256'b?????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b00011101 ;
      256'b????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b00010010 ;
      256'b???????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b11101010 ;
      256'b??????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b01111111 ;
      256'b?????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b01001110 ;
      256'b????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b11001101 ;
      256'b???????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b11011111 ;
      256'b??????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b00011011 ;
      256'b?????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b00100100 ;
      256'b????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b00001110 ;
      256'b???????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b00101111 ;
      256'b??????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b00001010 ;
      256'b?????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b00110111 ;
      256'b????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b00110000 ;
      256'b???????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b10011101 ;
      256'b??????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b01000110 ;
      256'b?????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b10010101 ;
      256'b????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b00001000 ;
      256'b???????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b00101010 ;
      256'b??????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b01100010 ;
      256'b?????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b10101011 ;
      256'b????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b11100010 ;
      256'b???????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b11111001 ;
      256'b??????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b11010001 ;
      256'b?????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b01010001 ;
      256'b????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b01101000 ;
      256'b???????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b10000011 ;
      256'b??????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b11110101 ;
      256'b?????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b01111110 ;
      256'b????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b01101100 ;
      256'b???????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b01001100 ;
      256'b??????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b00111101 ;
      256'b?????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b11100001 ;
      256'b????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b01110101 ;
      256'b???????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b10011011 ;
      256'b??????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b11100100 ;
      256'b?????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b01010011 ;
      256'b????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b00100011 ;
      256'b???????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b01000101 ;
      256'b??????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b01011111 ;
      256'b?????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b10110011 ;
      256'b????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b01000001 ;
      256'b???????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b11111011 ;
      256'b??????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b10001110 ;
      256'b?????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b10110010 ;
      256'b????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b11101111 ;
      256'b???????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b11111010 ;
      256'b??????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b10001001 ;
      256'b?????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b00011111 ;
      256'b????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b10001111 ;
      256'b???????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b11101100 ;
      256'b??????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b01001101 ;
      256'b?????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b10110101 ;
      256'b????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b11100111 ;
      256'b???????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b01010110 ;
      256'b??????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b11001110 ;
      256'b?????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b00000010 ;
      256'b????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b01100000 ;
      256'b???????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b10010001 ;
      256'b??????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b11011110 ;
      256'b?????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b11010110 ;
      256'b????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b11111111 ;
      256'b???1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b11110110 ;
      256'b??1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b11101110 ;
      256'b?1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b11111000 ;
      256'b1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b11000110 ;
      default:
        _2837_ = \t2.t2.s4.out ;
    endcase
  end
  assign p23[15:8] = \t2.t3.s0.out ^ \t2.t3.s4.out ;
  always @(posedge clk)
      \t2.t3.s0.out <= _2838_;
  wire [255:0] fangyuan23;
  assign fangyuan23 = { _3094_, _3093_, _3092_, _3091_, _3090_, _3089_, _3088_, _3087_, _3086_, _3085_, _3084_, _3083_, _3082_, _3081_, _3080_, _3079_, _3078_, _3077_, _3076_, _3075_, _3074_, _3073_, _3072_, _3071_, _3070_, _3069_, _3068_, _3067_, _3066_, _3065_, _3064_, _3063_, _3062_, _3061_, _3060_, _3059_, _3058_, _3057_, _3056_, _3055_, _3054_, _3053_, _3052_, _3051_, _3050_, _3049_, _3048_, _3047_, _3046_, _3045_, _3044_, _3043_, _3042_, _3041_, _3040_, _3039_, _3038_, _3037_, _3036_, _3035_, _3034_, _3033_, _3032_, _3031_, _3030_, _3029_, _3028_, _3027_, _3026_, _3025_, _3024_, _3023_, _3022_, _3021_, _3020_, _3019_, _3018_, _3017_, _3016_, _3015_, _3014_, _3013_, _3012_, _3011_, _3010_, _3009_, _3008_, _3007_, _3006_, _3005_, _3004_, _3003_, _3002_, _3001_, _3000_, _2999_, _2998_, _2997_, _2996_, _2995_, _2994_, _2993_, _2992_, _2991_, _2990_, _2989_, _2988_, _2987_, _2986_, _2985_, _2984_, _2983_, _2982_, _2981_, _2980_, _2979_, _2978_, _2977_, _2976_, _2975_, _2974_, _2973_, _2972_, _2971_, _2970_, _2969_, _2968_, _2967_, _2966_, _2965_, _2964_, _2963_, _2962_, _2961_, _2960_, _2959_, _2958_, _2957_, _2956_, _2955_, _2954_, _2953_, _2952_, _2951_, _2950_, _2949_, _2948_, _2947_, _2946_, _2945_, _2944_, _2943_, _2942_, _2941_, _2940_, _2939_, _2938_, _2937_, _2936_, _2935_, _2934_, _2933_, _2932_, _2931_, _2930_, _2929_, _2928_, _2927_, _2926_, _2925_, _2924_, _2923_, _2922_, _2921_, _2920_, _2919_, _2918_, _2917_, _2916_, _2915_, _2914_, _2913_, _2912_, _2911_, _2910_, _2909_, _2908_, _2907_, _2906_, _2905_, _2904_, _2903_, _2902_, _2901_, _2900_, _2899_, _2898_, _2897_, _2896_, _2895_, _2894_, _2893_, _2892_, _2891_, _2890_, _2889_, _2888_, _2887_, _2886_, _2885_, _2884_, _2883_, _2882_, _2881_, _2880_, _2879_, _2878_, _2877_, _2876_, _2875_, _2874_, _2873_, _2872_, _2871_, _2870_, _2869_, _2868_, _2867_, _2866_, _2865_, _2864_, _2863_, _2862_, _2861_, _2860_, _2859_, _2858_, _2857_, _2856_, _2855_, _2854_, _2853_, _2852_, _2851_, _2850_, _2849_, _2848_, _2847_, _2846_, _2845_, _2844_, _2843_, _2842_, _2841_, _2840_, _2839_ };

  always @(\t2.t3.s0.out or fangyuan23) begin
    casez (fangyuan23)
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1 :
        _2838_ = 8'b00010110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1? :
        _2838_ = 8'b10111011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?? :
        _2838_ = 8'b01010100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??? :
        _2838_ = 8'b10110000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???? :
        _2838_ = 8'b00001111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????? :
        _2838_ = 8'b00101101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????? :
        _2838_ = 8'b10011001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????? :
        _2838_ = 8'b01000001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????? :
        _2838_ = 8'b01101000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????? :
        _2838_ = 8'b01000010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????? :
        _2838_ = 8'b11100110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????? :
        _2838_ = 8'b10111111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????? :
        _2838_ = 8'b00001101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????? :
        _2838_ = 8'b10001001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????? :
        _2838_ = 8'b10100001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????? :
        _2838_ = 8'b10001100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????? :
        _2838_ = 8'b11011111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????? :
        _2838_ = 8'b00101000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????? :
        _2838_ = 8'b01010101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????? :
        _2838_ = 8'b11001110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????? :
        _2838_ = 8'b11101001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????? :
        _2838_ = 8'b10000111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????? :
        _2838_ = 8'b00011110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????? :
        _2838_ = 8'b10011011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????? :
        _2838_ = 8'b10010100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????? :
        _2838_ = 8'b10001110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????? :
        _2838_ = 8'b11011001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????? :
        _2838_ = 8'b01101001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????? :
        _2838_ = 8'b00010001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????? :
        _2838_ = 8'b10011000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????? :
        _2838_ = 8'b11111000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????? :
        _2838_ = 8'b11100001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????? :
        _2838_ = 8'b10011110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????? :
        _2838_ = 8'b00011101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????? :
        _2838_ = 8'b11000001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????? :
        _2838_ = 8'b10000110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????? :
        _2838_ = 8'b10111001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????? :
        _2838_ = 8'b01010111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????? :
        _2838_ = 8'b00110101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????? :
        _2838_ = 8'b01100001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????? :
        _2838_ = 8'b00001110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????? :
        _2838_ = 8'b11110110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????? :
        _2838_ = 8'b00000011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????? :
        _2838_ = 8'b01001000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????? :
        _2838_ = 8'b01100110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????? :
        _2838_ = 8'b10110101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????? :
        _2838_ = 8'b00111110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????? :
        _2838_ = 8'b01110000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????? :
        _2838_ = 8'b10001010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????? :
        _2838_ = 8'b10001011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????? :
        _2838_ = 8'b10111101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????? :
        _2838_ = 8'b01001011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????? :
        _2838_ = 8'b00011111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????? :
        _2838_ = 8'b01110100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????? :
        _2838_ = 8'b11011101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????? :
        _2838_ = 8'b11101000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????? :
        _2838_ = 8'b11000110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????? :
        _2838_ = 8'b10110100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????? :
        _2838_ = 8'b10100110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????? :
        _2838_ = 8'b00011100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????? :
        _2838_ = 8'b00101110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????? :
        _2838_ = 8'b00100101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????? :
        _2838_ = 8'b01111000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????? :
        _2838_ = 8'b10111010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????? :
        _2838_ = 8'b00001000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b10101110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b01111010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b01100101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b11101010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b11110100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b01010110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b01101100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b10101001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b01001110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b11010101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b10001101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b01101101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b00110111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b11001000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b11100111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b01111001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b11100100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b10010101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b10010001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b01100010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b10101100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b11010011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b11000010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b01011100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b00100100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b00000110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b01001001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b00001010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b00111010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b00110010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b11100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b11011011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b00001011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b01011110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b11011110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b00010100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b10111000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b11101110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b01000110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b10001000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b10010000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b00101010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b00100010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b11011100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b01001111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b10000001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b01100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b01110011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b00011001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b01011101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b01100100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b00111101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b01111110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b10100111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b11000100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b00010111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b01000100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b10010111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b01011111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b11101100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b00010011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b00001100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b11001101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b11010010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b11110011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b11111111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b00010000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b00100001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b11011010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b10110110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b10111100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b11110101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b00111000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b10011101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b10010010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b10001111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b01000000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b10100011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b01010001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b10101000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b10011111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b00111100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b01010000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b01111111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b00000010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b11111001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b01000101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b10000101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b00110011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b01001101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b01000011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b11111011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b10101010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b11101111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b11010000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b11001111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b01011000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b01001100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b01001010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b00111001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b10111110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b11001011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b01101010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b01011011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b10110001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b11111100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b00100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b11101101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b00000000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b11010001 ;
      256'b????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b01010011 ;
      256'b???????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b10000100 ;
      256'b??????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b00101111 ;
      256'b?????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b11100011 ;
      256'b????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b00101001 ;
      256'b???????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b10110011 ;
      256'b??????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b11010110 ;
      256'b?????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b00111011 ;
      256'b????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b01010010 ;
      256'b???????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b10100000 ;
      256'b??????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b01011010 ;
      256'b?????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b01101110 ;
      256'b????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b00011011 ;
      256'b???????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b00011010 ;
      256'b??????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b00101100 ;
      256'b?????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b10000011 ;
      256'b????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b00001001 ;
      256'b???????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b01110101 ;
      256'b??????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b10110010 ;
      256'b?????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b00100111 ;
      256'b????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b11101011 ;
      256'b???????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b11100010 ;
      256'b??????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b10000000 ;
      256'b?????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b00010010 ;
      256'b????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b00000111 ;
      256'b???????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b10011010 ;
      256'b??????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b00000101 ;
      256'b?????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b10010110 ;
      256'b????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b00011000 ;
      256'b???????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b11000011 ;
      256'b??????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b00100011 ;
      256'b?????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b11000111 ;
      256'b????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b00000100 ;
      256'b???????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b00010101 ;
      256'b??????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b00110001 ;
      256'b?????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b11011000 ;
      256'b????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b01110001 ;
      256'b???????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b11110001 ;
      256'b??????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b11100101 ;
      256'b?????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b10100101 ;
      256'b????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b00110100 ;
      256'b???????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b11001100 ;
      256'b??????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b11110111 ;
      256'b?????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b00111111 ;
      256'b????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b00110110 ;
      256'b???????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b00100110 ;
      256'b??????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b10010011 ;
      256'b?????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b11111101 ;
      256'b????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b10110111 ;
      256'b???????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b11000000 ;
      256'b??????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b01110010 ;
      256'b?????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b10100100 ;
      256'b????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b10011100 ;
      256'b???????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b10101111 ;
      256'b??????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b10100010 ;
      256'b?????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b11010100 ;
      256'b????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b10101101 ;
      256'b???????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b11110000 ;
      256'b??????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b01000111 ;
      256'b?????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b01011001 ;
      256'b????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b11111010 ;
      256'b???????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b01111101 ;
      256'b??????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b11001001 ;
      256'b?????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b10000010 ;
      256'b????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b11001010 ;
      256'b???????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b01110110 ;
      256'b??????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b10101011 ;
      256'b?????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b11010111 ;
      256'b????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b11111110 ;
      256'b???????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b00101011 ;
      256'b??????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b01100111 ;
      256'b?????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b00000001 ;
      256'b????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b00110000 ;
      256'b???????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b11000101 ;
      256'b??????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b01101111 ;
      256'b?????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b01101011 ;
      256'b????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b11110010 ;
      256'b???1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b01111011 ;
      256'b??1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b01110111 ;
      256'b?1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b01111100 ;
      256'b1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b01100011 ;
      default:
        _2838_ = \t2.t3.s0.out ;
    endcase
  end
  assign _2839_ = state_in[39:32] == 8'b11111111;
  assign _2840_ = state_in[39:32] == 8'b11111110;
  assign _2841_ = state_in[39:32] == 8'b11111101;
  assign _2842_ = state_in[39:32] == 8'b11111100;
  assign _2843_ = state_in[39:32] == 8'b11111011;
  assign _2844_ = state_in[39:32] == 8'b11111010;
  assign _2845_ = state_in[39:32] == 8'b11111001;
  assign _2846_ = state_in[39:32] == 8'b11111000;
  assign _2847_ = state_in[39:32] == 8'b11110111;
  assign _2848_ = state_in[39:32] == 8'b11110110;
  assign _2849_ = state_in[39:32] == 8'b11110101;
  assign _2850_ = state_in[39:32] == 8'b11110100;
  assign _2851_ = state_in[39:32] == 8'b11110011;
  assign _2852_ = state_in[39:32] == 8'b11110010;
  assign _2853_ = state_in[39:32] == 8'b11110001;
  assign _2854_ = state_in[39:32] == 8'b11110000;
  assign _2855_ = state_in[39:32] == 8'b11101111;
  assign _2856_ = state_in[39:32] == 8'b11101110;
  assign _2857_ = state_in[39:32] == 8'b11101101;
  assign _2858_ = state_in[39:32] == 8'b11101100;
  assign _2859_ = state_in[39:32] == 8'b11101011;
  assign _2860_ = state_in[39:32] == 8'b11101010;
  assign _2861_ = state_in[39:32] == 8'b11101001;
  assign _2862_ = state_in[39:32] == 8'b11101000;
  assign _2863_ = state_in[39:32] == 8'b11100111;
  assign _2864_ = state_in[39:32] == 8'b11100110;
  assign _2865_ = state_in[39:32] == 8'b11100101;
  assign _2866_ = state_in[39:32] == 8'b11100100;
  assign _2867_ = state_in[39:32] == 8'b11100011;
  assign _2868_ = state_in[39:32] == 8'b11100010;
  assign _2869_ = state_in[39:32] == 8'b11100001;
  assign _2870_ = state_in[39:32] == 8'b11100000;
  assign _2871_ = state_in[39:32] == 8'b11011111;
  assign _2872_ = state_in[39:32] == 8'b11011110;
  assign _2873_ = state_in[39:32] == 8'b11011101;
  assign _2874_ = state_in[39:32] == 8'b11011100;
  assign _2875_ = state_in[39:32] == 8'b11011011;
  assign _2876_ = state_in[39:32] == 8'b11011010;
  assign _2877_ = state_in[39:32] == 8'b11011001;
  assign _2878_ = state_in[39:32] == 8'b11011000;
  assign _2879_ = state_in[39:32] == 8'b11010111;
  assign _2880_ = state_in[39:32] == 8'b11010110;
  assign _2881_ = state_in[39:32] == 8'b11010101;
  assign _2882_ = state_in[39:32] == 8'b11010100;
  assign _2883_ = state_in[39:32] == 8'b11010011;
  assign _2884_ = state_in[39:32] == 8'b11010010;
  assign _2885_ = state_in[39:32] == 8'b11010001;
  assign _2886_ = state_in[39:32] == 8'b11010000;
  assign _2887_ = state_in[39:32] == 8'b11001111;
  assign _2888_ = state_in[39:32] == 8'b11001110;
  assign _2889_ = state_in[39:32] == 8'b11001101;
  assign _2890_ = state_in[39:32] == 8'b11001100;
  assign _2891_ = state_in[39:32] == 8'b11001011;
  assign _2892_ = state_in[39:32] == 8'b11001010;
  assign _2893_ = state_in[39:32] == 8'b11001001;
  assign _2894_ = state_in[39:32] == 8'b11001000;
  assign _2895_ = state_in[39:32] == 8'b11000111;
  assign _2896_ = state_in[39:32] == 8'b11000110;
  assign _2897_ = state_in[39:32] == 8'b11000101;
  assign _2898_ = state_in[39:32] == 8'b11000100;
  assign _2899_ = state_in[39:32] == 8'b11000011;
  assign _2900_ = state_in[39:32] == 8'b11000010;
  assign _2901_ = state_in[39:32] == 8'b11000001;
  assign _2902_ = state_in[39:32] == 8'b11000000;
  assign _2903_ = state_in[39:32] == 8'b10111111;
  assign _2904_ = state_in[39:32] == 8'b10111110;
  assign _2905_ = state_in[39:32] == 8'b10111101;
  assign _2906_ = state_in[39:32] == 8'b10111100;
  assign _2907_ = state_in[39:32] == 8'b10111011;
  assign _2908_ = state_in[39:32] == 8'b10111010;
  assign _2909_ = state_in[39:32] == 8'b10111001;
  assign _2910_ = state_in[39:32] == 8'b10111000;
  assign _2911_ = state_in[39:32] == 8'b10110111;
  assign _2912_ = state_in[39:32] == 8'b10110110;
  assign _2913_ = state_in[39:32] == 8'b10110101;
  assign _2914_ = state_in[39:32] == 8'b10110100;
  assign _2915_ = state_in[39:32] == 8'b10110011;
  assign _2916_ = state_in[39:32] == 8'b10110010;
  assign _2917_ = state_in[39:32] == 8'b10110001;
  assign _2918_ = state_in[39:32] == 8'b10110000;
  assign _2919_ = state_in[39:32] == 8'b10101111;
  assign _2920_ = state_in[39:32] == 8'b10101110;
  assign _2921_ = state_in[39:32] == 8'b10101101;
  assign _2922_ = state_in[39:32] == 8'b10101100;
  assign _2923_ = state_in[39:32] == 8'b10101011;
  assign _2924_ = state_in[39:32] == 8'b10101010;
  assign _2925_ = state_in[39:32] == 8'b10101001;
  assign _2926_ = state_in[39:32] == 8'b10101000;
  assign _2927_ = state_in[39:32] == 8'b10100111;
  assign _2928_ = state_in[39:32] == 8'b10100110;
  assign _2929_ = state_in[39:32] == 8'b10100101;
  assign _2930_ = state_in[39:32] == 8'b10100100;
  assign _2931_ = state_in[39:32] == 8'b10100011;
  assign _2932_ = state_in[39:32] == 8'b10100010;
  assign _2933_ = state_in[39:32] == 8'b10100001;
  assign _2934_ = state_in[39:32] == 8'b10100000;
  assign _2935_ = state_in[39:32] == 8'b10011111;
  assign _2936_ = state_in[39:32] == 8'b10011110;
  assign _2937_ = state_in[39:32] == 8'b10011101;
  assign _2938_ = state_in[39:32] == 8'b10011100;
  assign _2939_ = state_in[39:32] == 8'b10011011;
  assign _2940_ = state_in[39:32] == 8'b10011010;
  assign _2941_ = state_in[39:32] == 8'b10011001;
  assign _2942_ = state_in[39:32] == 8'b10011000;
  assign _2943_ = state_in[39:32] == 8'b10010111;
  assign _2944_ = state_in[39:32] == 8'b10010110;
  assign _2945_ = state_in[39:32] == 8'b10010101;
  assign _2946_ = state_in[39:32] == 8'b10010100;
  assign _2947_ = state_in[39:32] == 8'b10010011;
  assign _2948_ = state_in[39:32] == 8'b10010010;
  assign _2949_ = state_in[39:32] == 8'b10010001;
  assign _2950_ = state_in[39:32] == 8'b10010000;
  assign _2951_ = state_in[39:32] == 8'b10001111;
  assign _2952_ = state_in[39:32] == 8'b10001110;
  assign _2953_ = state_in[39:32] == 8'b10001101;
  assign _2954_ = state_in[39:32] == 8'b10001100;
  assign _2955_ = state_in[39:32] == 8'b10001011;
  assign _2956_ = state_in[39:32] == 8'b10001010;
  assign _2957_ = state_in[39:32] == 8'b10001001;
  assign _2958_ = state_in[39:32] == 8'b10001000;
  assign _2959_ = state_in[39:32] == 8'b10000111;
  assign _2960_ = state_in[39:32] == 8'b10000110;
  assign _2961_ = state_in[39:32] == 8'b10000101;
  assign _2962_ = state_in[39:32] == 8'b10000100;
  assign _2963_ = state_in[39:32] == 8'b10000011;
  assign _2964_ = state_in[39:32] == 8'b10000010;
  assign _2965_ = state_in[39:32] == 8'b10000001;
  assign _2966_ = state_in[39:32] == 8'b10000000;
  assign _2967_ = state_in[39:32] == 7'b1111111;
  assign _2968_ = state_in[39:32] == 7'b1111110;
  assign _2969_ = state_in[39:32] == 7'b1111101;
  assign _2970_ = state_in[39:32] == 7'b1111100;
  assign _2971_ = state_in[39:32] == 7'b1111011;
  assign _2972_ = state_in[39:32] == 7'b1111010;
  assign _2973_ = state_in[39:32] == 7'b1111001;
  assign _2974_ = state_in[39:32] == 7'b1111000;
  assign _2975_ = state_in[39:32] == 7'b1110111;
  assign _2976_ = state_in[39:32] == 7'b1110110;
  assign _2977_ = state_in[39:32] == 7'b1110101;
  assign _2978_ = state_in[39:32] == 7'b1110100;
  assign _2979_ = state_in[39:32] == 7'b1110011;
  assign _2980_ = state_in[39:32] == 7'b1110010;
  assign _2981_ = state_in[39:32] == 7'b1110001;
  assign _2982_ = state_in[39:32] == 7'b1110000;
  assign _2983_ = state_in[39:32] == 7'b1101111;
  assign _2984_ = state_in[39:32] == 7'b1101110;
  assign _2985_ = state_in[39:32] == 7'b1101101;
  assign _2986_ = state_in[39:32] == 7'b1101100;
  assign _2987_ = state_in[39:32] == 7'b1101011;
  assign _2988_ = state_in[39:32] == 7'b1101010;
  assign _2989_ = state_in[39:32] == 7'b1101001;
  assign _2990_ = state_in[39:32] == 7'b1101000;
  assign _2991_ = state_in[39:32] == 7'b1100111;
  assign _2992_ = state_in[39:32] == 7'b1100110;
  assign _2993_ = state_in[39:32] == 7'b1100101;
  assign _2994_ = state_in[39:32] == 7'b1100100;
  assign _2995_ = state_in[39:32] == 7'b1100011;
  assign _2996_ = state_in[39:32] == 7'b1100010;
  assign _2997_ = state_in[39:32] == 7'b1100001;
  assign _2998_ = state_in[39:32] == 7'b1100000;
  assign _2999_ = state_in[39:32] == 7'b1011111;
  assign _3000_ = state_in[39:32] == 7'b1011110;
  assign _3001_ = state_in[39:32] == 7'b1011101;
  assign _3002_ = state_in[39:32] == 7'b1011100;
  assign _3003_ = state_in[39:32] == 7'b1011011;
  assign _3004_ = state_in[39:32] == 7'b1011010;
  assign _3005_ = state_in[39:32] == 7'b1011001;
  assign _3006_ = state_in[39:32] == 7'b1011000;
  assign _3007_ = state_in[39:32] == 7'b1010111;
  assign _3008_ = state_in[39:32] == 7'b1010110;
  assign _3009_ = state_in[39:32] == 7'b1010101;
  assign _3010_ = state_in[39:32] == 7'b1010100;
  assign _3011_ = state_in[39:32] == 7'b1010011;
  assign _3012_ = state_in[39:32] == 7'b1010010;
  assign _3013_ = state_in[39:32] == 7'b1010001;
  assign _3014_ = state_in[39:32] == 7'b1010000;
  assign _3015_ = state_in[39:32] == 7'b1001111;
  assign _3016_ = state_in[39:32] == 7'b1001110;
  assign _3017_ = state_in[39:32] == 7'b1001101;
  assign _3018_ = state_in[39:32] == 7'b1001100;
  assign _3019_ = state_in[39:32] == 7'b1001011;
  assign _3020_ = state_in[39:32] == 7'b1001010;
  assign _3021_ = state_in[39:32] == 7'b1001001;
  assign _3022_ = state_in[39:32] == 7'b1001000;
  assign _3023_ = state_in[39:32] == 7'b1000111;
  assign _3024_ = state_in[39:32] == 7'b1000110;
  assign _3025_ = state_in[39:32] == 7'b1000101;
  assign _3026_ = state_in[39:32] == 7'b1000100;
  assign _3027_ = state_in[39:32] == 7'b1000011;
  assign _3028_ = state_in[39:32] == 7'b1000010;
  assign _3029_ = state_in[39:32] == 7'b1000001;
  assign _3030_ = state_in[39:32] == 7'b1000000;
  assign _3031_ = state_in[39:32] == 6'b111111;
  assign _3032_ = state_in[39:32] == 6'b111110;
  assign _3033_ = state_in[39:32] == 6'b111101;
  assign _3034_ = state_in[39:32] == 6'b111100;
  assign _3035_ = state_in[39:32] == 6'b111011;
  assign _3036_ = state_in[39:32] == 6'b111010;
  assign _3037_ = state_in[39:32] == 6'b111001;
  assign _3038_ = state_in[39:32] == 6'b111000;
  assign _3039_ = state_in[39:32] == 6'b110111;
  assign _3040_ = state_in[39:32] == 6'b110110;
  assign _3041_ = state_in[39:32] == 6'b110101;
  assign _3042_ = state_in[39:32] == 6'b110100;
  assign _3043_ = state_in[39:32] == 6'b110011;
  assign _3044_ = state_in[39:32] == 6'b110010;
  assign _3045_ = state_in[39:32] == 6'b110001;
  assign _3046_ = state_in[39:32] == 6'b110000;
  assign _3047_ = state_in[39:32] == 6'b101111;
  assign _3048_ = state_in[39:32] == 6'b101110;
  assign _3049_ = state_in[39:32] == 6'b101101;
  assign _3050_ = state_in[39:32] == 6'b101100;
  assign _3051_ = state_in[39:32] == 6'b101011;
  assign _3052_ = state_in[39:32] == 6'b101010;
  assign _3053_ = state_in[39:32] == 6'b101001;
  assign _3054_ = state_in[39:32] == 6'b101000;
  assign _3055_ = state_in[39:32] == 6'b100111;
  assign _3056_ = state_in[39:32] == 6'b100110;
  assign _3057_ = state_in[39:32] == 6'b100101;
  assign _3058_ = state_in[39:32] == 6'b100100;
  assign _3059_ = state_in[39:32] == 6'b100011;
  assign _3060_ = state_in[39:32] == 6'b100010;
  assign _3061_ = state_in[39:32] == 6'b100001;
  assign _3062_ = state_in[39:32] == 6'b100000;
  assign _3063_ = state_in[39:32] == 5'b11111;
  assign _3064_ = state_in[39:32] == 5'b11110;
  assign _3065_ = state_in[39:32] == 5'b11101;
  assign _3066_ = state_in[39:32] == 5'b11100;
  assign _3067_ = state_in[39:32] == 5'b11011;
  assign _3068_ = state_in[39:32] == 5'b11010;
  assign _3069_ = state_in[39:32] == 5'b11001;
  assign _3070_ = state_in[39:32] == 5'b11000;
  assign _3071_ = state_in[39:32] == 5'b10111;
  assign _3072_ = state_in[39:32] == 5'b10110;
  assign _3073_ = state_in[39:32] == 5'b10101;
  assign _3074_ = state_in[39:32] == 5'b10100;
  assign _3075_ = state_in[39:32] == 5'b10011;
  assign _3076_ = state_in[39:32] == 5'b10010;
  assign _3077_ = state_in[39:32] == 5'b10001;
  assign _3078_ = state_in[39:32] == 5'b10000;
  assign _3079_ = state_in[39:32] == 4'b1111;
  assign _3080_ = state_in[39:32] == 4'b1110;
  assign _3081_ = state_in[39:32] == 4'b1101;
  assign _3082_ = state_in[39:32] == 4'b1100;
  assign _3083_ = state_in[39:32] == 4'b1011;
  assign _3084_ = state_in[39:32] == 4'b1010;
  assign _3085_ = state_in[39:32] == 4'b1001;
  assign _3086_ = state_in[39:32] == 4'b1000;
  assign _3087_ = state_in[39:32] == 3'b111;
  assign _3088_ = state_in[39:32] == 3'b110;
  assign _3089_ = state_in[39:32] == 3'b101;
  assign _3090_ = state_in[39:32] == 3'b100;
  assign _3091_ = state_in[39:32] == 2'b11;
  assign _3092_ = state_in[39:32] == 2'b10;
  assign _3093_ = state_in[39:32] == 1'b1;
  assign _3094_ = ! state_in[39:32];
  always @(posedge clk)
      \t2.t3.s4.out <= _3095_;
  wire [255:0] fangyuan24;
  assign fangyuan24 = { _3094_, _3093_, _3092_, _3091_, _3090_, _3089_, _3088_, _3087_, _3086_, _3085_, _3084_, _3083_, _3082_, _3081_, _3080_, _3079_, _3078_, _3077_, _3076_, _3075_, _3074_, _3073_, _3072_, _3071_, _3070_, _3069_, _3068_, _3067_, _3066_, _3065_, _3064_, _3063_, _3062_, _3061_, _3060_, _3059_, _3058_, _3057_, _3056_, _3055_, _3054_, _3053_, _3052_, _3051_, _3050_, _3049_, _3048_, _3047_, _3046_, _3045_, _3044_, _3043_, _3042_, _3041_, _3040_, _3039_, _3038_, _3037_, _3036_, _3035_, _3034_, _3033_, _3032_, _3031_, _3030_, _3029_, _3028_, _3027_, _3026_, _3025_, _3024_, _3023_, _3022_, _3021_, _3020_, _3019_, _3018_, _3017_, _3016_, _3015_, _3014_, _3013_, _3012_, _3011_, _3010_, _3009_, _3008_, _3007_, _3006_, _3005_, _3004_, _3003_, _3002_, _3001_, _3000_, _2999_, _2998_, _2997_, _2996_, _2995_, _2994_, _2993_, _2992_, _2991_, _2990_, _2989_, _2988_, _2987_, _2986_, _2985_, _2984_, _2983_, _2982_, _2981_, _2980_, _2979_, _2978_, _2977_, _2976_, _2975_, _2974_, _2973_, _2972_, _2971_, _2970_, _2969_, _2968_, _2967_, _2966_, _2965_, _2964_, _2963_, _2962_, _2961_, _2960_, _2959_, _2958_, _2957_, _2956_, _2955_, _2954_, _2953_, _2952_, _2951_, _2950_, _2949_, _2948_, _2947_, _2946_, _2945_, _2944_, _2943_, _2942_, _2941_, _2940_, _2939_, _2938_, _2937_, _2936_, _2935_, _2934_, _2933_, _2932_, _2931_, _2930_, _2929_, _2928_, _2927_, _2926_, _2925_, _2924_, _2923_, _2922_, _2921_, _2920_, _2919_, _2918_, _2917_, _2916_, _2915_, _2914_, _2913_, _2912_, _2911_, _2910_, _2909_, _2908_, _2907_, _2906_, _2905_, _2904_, _2903_, _2902_, _2901_, _2900_, _2899_, _2898_, _2897_, _2896_, _2895_, _2894_, _2893_, _2892_, _2891_, _2890_, _2889_, _2888_, _2887_, _2886_, _2885_, _2884_, _2883_, _2882_, _2881_, _2880_, _2879_, _2878_, _2877_, _2876_, _2875_, _2874_, _2873_, _2872_, _2871_, _2870_, _2869_, _2868_, _2867_, _2866_, _2865_, _2864_, _2863_, _2862_, _2861_, _2860_, _2859_, _2858_, _2857_, _2856_, _2855_, _2854_, _2853_, _2852_, _2851_, _2850_, _2849_, _2848_, _2847_, _2846_, _2845_, _2844_, _2843_, _2842_, _2841_, _2840_, _2839_ };

  always @(\t2.t3.s4.out or fangyuan24) begin
    casez (fangyuan24)
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1 :
        _3095_ = 8'b00101100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1? :
        _3095_ = 8'b01101101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?? :
        _3095_ = 8'b10101000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??? :
        _3095_ = 8'b01111011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???? :
        _3095_ = 8'b00011110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????? :
        _3095_ = 8'b01011010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????? :
        _3095_ = 8'b00101001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????? :
        _3095_ = 8'b10000010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????? :
        _3095_ = 8'b11010000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????? :
        _3095_ = 8'b10000100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????? :
        _3095_ = 8'b11010111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????? :
        _3095_ = 8'b01100101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????? :
        _3095_ = 8'b00011010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????? :
        _3095_ = 8'b00001001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????? :
        _3095_ = 8'b01011001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????? :
        _3095_ = 8'b00000011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????? :
        _3095_ = 8'b10100101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????? :
        _3095_ = 8'b01010000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????? :
        _3095_ = 8'b10101010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????? :
        _3095_ = 8'b10000111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????? :
        _3095_ = 8'b11001001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????? :
        _3095_ = 8'b00010101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????? :
        _3095_ = 8'b00111100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????? :
        _3095_ = 8'b00101101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????? :
        _3095_ = 8'b00110011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????? :
        _3095_ = 8'b00000111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????? :
        _3095_ = 8'b10101001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????? :
        _3095_ = 8'b11010010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????? :
        _3095_ = 8'b00100010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????? :
        _3095_ = 8'b00101011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????? :
        _3095_ = 8'b11101011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????? :
        _3095_ = 8'b11011001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????? :
        _3095_ = 8'b00100111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????? :
        _3095_ = 8'b00111010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????? :
        _3095_ = 8'b10011001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????? :
        _3095_ = 8'b00010111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????? :
        _3095_ = 8'b01101001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????? :
        _3095_ = 8'b10101110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????? :
        _3095_ = 8'b01101010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????? :
        _3095_ = 8'b11000010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????? :
        _3095_ = 8'b00011100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????? :
        _3095_ = 8'b11110111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????? :
        _3095_ = 8'b00000110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????? :
        _3095_ = 8'b10010000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????? :
        _3095_ = 8'b11001100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????? :
        _3095_ = 8'b01110001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????? :
        _3095_ = 8'b01111100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????? :
        _3095_ = 8'b11100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????? :
        _3095_ = 8'b00001111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????? :
        _3095_ = 8'b00001101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????? :
        _3095_ = 8'b01100001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????? :
        _3095_ = 8'b10010110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????? :
        _3095_ = 8'b00111110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????? :
        _3095_ = 8'b11101000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????? :
        _3095_ = 8'b10100001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????? :
        _3095_ = 8'b11001011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????? :
        _3095_ = 8'b10010111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????? :
        _3095_ = 8'b01110011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????? :
        _3095_ = 8'b01010111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????? :
        _3095_ = 8'b00111000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????? :
        _3095_ = 8'b01011100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????? :
        _3095_ = 8'b01001010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????? :
        _3095_ = 8'b11110000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????? :
        _3095_ = 8'b01101111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????? :
        _3095_ = 8'b00010000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b01000111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b11110100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b11001010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b11001111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b11110011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b10101100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b11011000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b01001001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b10011100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b10110001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b00000001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b11011010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b01101110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b10001011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b11010101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b11110010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b11010011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b00110001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b00111001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b11000100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b01000011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b10111101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b10011111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b10111000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b01001000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b00001100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b10010010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b00010100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b01110100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b01100100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b11011011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b10101101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b00010110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b10111100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b10100111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b00101000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b01101011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b11000111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b10001100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b00001011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b00111011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b01010100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b01000100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b10100011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b10011110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b00011001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b11000000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b11100110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b00110010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b10111010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b11001000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b01111010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b11111100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b01010101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b10010011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b00101110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b10001000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b00110101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b10111110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b11000011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b00100110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b00011000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b10000001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b10111111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b11111101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b11100101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b00100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b01000010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b10101111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b01110111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b01100011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b11110001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b01110000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b00100001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b00111111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b00000101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b10000000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b01011101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b10100010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b01001011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b00100101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b01111000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b10100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b11111110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b00000100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b11101001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b10001010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b00010001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b01100110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b10011010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b10000110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b11101101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b01001111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b11000101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b10111011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b10000101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b10110000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b10011000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b10010100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b01110010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b01100111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b10001101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b11010100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b10110110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b01111001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b11100011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b01000000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b11000001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b00000000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b10111001 ;
      256'b????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b10100110 ;
      256'b???????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b00010011 ;
      256'b??????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b01011110 ;
      256'b?????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b11011101 ;
      256'b????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b01010010 ;
      256'b???????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b01111101 ;
      256'b??????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b10110111 ;
      256'b?????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b01110110 ;
      256'b????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b10100100 ;
      256'b???????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b01011011 ;
      256'b??????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b10110100 ;
      256'b?????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b11011100 ;
      256'b????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b00110110 ;
      256'b???????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b00110100 ;
      256'b??????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b01011000 ;
      256'b?????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b00011101 ;
      256'b????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b00010010 ;
      256'b???????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b11101010 ;
      256'b??????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b01111111 ;
      256'b?????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b01001110 ;
      256'b????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b11001101 ;
      256'b???????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b11011111 ;
      256'b??????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b00011011 ;
      256'b?????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b00100100 ;
      256'b????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b00001110 ;
      256'b???????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b00101111 ;
      256'b??????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b00001010 ;
      256'b?????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b00110111 ;
      256'b????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b00110000 ;
      256'b???????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b10011101 ;
      256'b??????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b01000110 ;
      256'b?????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b10010101 ;
      256'b????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b00001000 ;
      256'b???????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b00101010 ;
      256'b??????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b01100010 ;
      256'b?????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b10101011 ;
      256'b????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b11100010 ;
      256'b???????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b11111001 ;
      256'b??????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b11010001 ;
      256'b?????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b01010001 ;
      256'b????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b01101000 ;
      256'b???????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b10000011 ;
      256'b??????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b11110101 ;
      256'b?????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b01111110 ;
      256'b????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b01101100 ;
      256'b???????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b01001100 ;
      256'b??????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b00111101 ;
      256'b?????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b11100001 ;
      256'b????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b01110101 ;
      256'b???????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b10011011 ;
      256'b??????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b11100100 ;
      256'b?????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b01010011 ;
      256'b????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b00100011 ;
      256'b???????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b01000101 ;
      256'b??????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b01011111 ;
      256'b?????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b10110011 ;
      256'b????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b01000001 ;
      256'b???????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b11111011 ;
      256'b??????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b10001110 ;
      256'b?????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b10110010 ;
      256'b????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b11101111 ;
      256'b???????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b11111010 ;
      256'b??????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b10001001 ;
      256'b?????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b00011111 ;
      256'b????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b10001111 ;
      256'b???????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b11101100 ;
      256'b??????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b01001101 ;
      256'b?????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b10110101 ;
      256'b????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b11100111 ;
      256'b???????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b01010110 ;
      256'b??????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b11001110 ;
      256'b?????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b00000010 ;
      256'b????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b01100000 ;
      256'b???????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b10010001 ;
      256'b??????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b11011110 ;
      256'b?????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b11010110 ;
      256'b????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b11111111 ;
      256'b???1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b11110110 ;
      256'b??1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b11101110 ;
      256'b?1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b11111000 ;
      256'b1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b11000110 ;
      default:
        _3095_ = \t2.t3.s4.out ;
    endcase
  end
  assign p30[7:0] = \t3.t0.s0.out ^ \t3.t0.s4.out ;
  always @(posedge clk)
      \t3.t0.s0.out <= _3096_;
  wire [255:0] fangyuan25;
  assign fangyuan25 = { _3352_, _3351_, _3350_, _3349_, _3348_, _3347_, _3346_, _3345_, _3344_, _3343_, _3342_, _3341_, _3340_, _3339_, _3338_, _3337_, _3336_, _3335_, _3334_, _3333_, _3332_, _3331_, _3330_, _3329_, _3328_, _3327_, _3326_, _3325_, _3324_, _3323_, _3322_, _3321_, _3320_, _3319_, _3318_, _3317_, _3316_, _3315_, _3314_, _3313_, _3312_, _3311_, _3310_, _3309_, _3308_, _3307_, _3306_, _3305_, _3304_, _3303_, _3302_, _3301_, _3300_, _3299_, _3298_, _3297_, _3296_, _3295_, _3294_, _3293_, _3292_, _3291_, _3290_, _3289_, _3288_, _3287_, _3286_, _3285_, _3284_, _3283_, _3282_, _3281_, _3280_, _3279_, _3278_, _3277_, _3276_, _3275_, _3274_, _3273_, _3272_, _3271_, _3270_, _3269_, _3268_, _3267_, _3266_, _3265_, _3264_, _3263_, _3262_, _3261_, _3260_, _3259_, _3258_, _3257_, _3256_, _3255_, _3254_, _3253_, _3252_, _3251_, _3250_, _3249_, _3248_, _3247_, _3246_, _3245_, _3244_, _3243_, _3242_, _3241_, _3240_, _3239_, _3238_, _3237_, _3236_, _3235_, _3234_, _3233_, _3232_, _3231_, _3230_, _3229_, _3228_, _3227_, _3226_, _3225_, _3224_, _3223_, _3222_, _3221_, _3220_, _3219_, _3218_, _3217_, _3216_, _3215_, _3214_, _3213_, _3212_, _3211_, _3210_, _3209_, _3208_, _3207_, _3206_, _3205_, _3204_, _3203_, _3202_, _3201_, _3200_, _3199_, _3198_, _3197_, _3196_, _3195_, _3194_, _3193_, _3192_, _3191_, _3190_, _3189_, _3188_, _3187_, _3186_, _3185_, _3184_, _3183_, _3182_, _3181_, _3180_, _3179_, _3178_, _3177_, _3176_, _3175_, _3174_, _3173_, _3172_, _3171_, _3170_, _3169_, _3168_, _3167_, _3166_, _3165_, _3164_, _3163_, _3162_, _3161_, _3160_, _3159_, _3158_, _3157_, _3156_, _3155_, _3154_, _3153_, _3152_, _3151_, _3150_, _3149_, _3148_, _3147_, _3146_, _3145_, _3144_, _3143_, _3142_, _3141_, _3140_, _3139_, _3138_, _3137_, _3136_, _3135_, _3134_, _3133_, _3132_, _3131_, _3130_, _3129_, _3128_, _3127_, _3126_, _3125_, _3124_, _3123_, _3122_, _3121_, _3120_, _3119_, _3118_, _3117_, _3116_, _3115_, _3114_, _3113_, _3112_, _3111_, _3110_, _3109_, _3108_, _3107_, _3106_, _3105_, _3104_, _3103_, _3102_, _3101_, _3100_, _3099_, _3098_, _3097_ };

  always @(\t3.t0.s0.out or fangyuan25) begin
    casez (fangyuan25)
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1 :
        _3096_ = 8'b00010110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1? :
        _3096_ = 8'b10111011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?? :
        _3096_ = 8'b01010100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??? :
        _3096_ = 8'b10110000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???? :
        _3096_ = 8'b00001111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????? :
        _3096_ = 8'b00101101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????? :
        _3096_ = 8'b10011001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????? :
        _3096_ = 8'b01000001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????? :
        _3096_ = 8'b01101000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????? :
        _3096_ = 8'b01000010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????? :
        _3096_ = 8'b11100110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????? :
        _3096_ = 8'b10111111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????? :
        _3096_ = 8'b00001101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????? :
        _3096_ = 8'b10001001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????? :
        _3096_ = 8'b10100001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????? :
        _3096_ = 8'b10001100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????? :
        _3096_ = 8'b11011111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????? :
        _3096_ = 8'b00101000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????? :
        _3096_ = 8'b01010101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????? :
        _3096_ = 8'b11001110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????? :
        _3096_ = 8'b11101001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????? :
        _3096_ = 8'b10000111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????? :
        _3096_ = 8'b00011110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????? :
        _3096_ = 8'b10011011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????? :
        _3096_ = 8'b10010100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????? :
        _3096_ = 8'b10001110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????? :
        _3096_ = 8'b11011001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????? :
        _3096_ = 8'b01101001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????? :
        _3096_ = 8'b00010001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????? :
        _3096_ = 8'b10011000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????? :
        _3096_ = 8'b11111000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????? :
        _3096_ = 8'b11100001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????? :
        _3096_ = 8'b10011110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????? :
        _3096_ = 8'b00011101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????? :
        _3096_ = 8'b11000001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????? :
        _3096_ = 8'b10000110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????? :
        _3096_ = 8'b10111001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????? :
        _3096_ = 8'b01010111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????? :
        _3096_ = 8'b00110101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????? :
        _3096_ = 8'b01100001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????? :
        _3096_ = 8'b00001110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????? :
        _3096_ = 8'b11110110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????? :
        _3096_ = 8'b00000011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????? :
        _3096_ = 8'b01001000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????? :
        _3096_ = 8'b01100110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????? :
        _3096_ = 8'b10110101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????? :
        _3096_ = 8'b00111110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????? :
        _3096_ = 8'b01110000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????? :
        _3096_ = 8'b10001010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????? :
        _3096_ = 8'b10001011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????? :
        _3096_ = 8'b10111101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????? :
        _3096_ = 8'b01001011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????? :
        _3096_ = 8'b00011111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????? :
        _3096_ = 8'b01110100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????? :
        _3096_ = 8'b11011101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????? :
        _3096_ = 8'b11101000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????? :
        _3096_ = 8'b11000110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????? :
        _3096_ = 8'b10110100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????? :
        _3096_ = 8'b10100110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????? :
        _3096_ = 8'b00011100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????? :
        _3096_ = 8'b00101110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????? :
        _3096_ = 8'b00100101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????? :
        _3096_ = 8'b01111000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????? :
        _3096_ = 8'b10111010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????? :
        _3096_ = 8'b00001000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b10101110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b01111010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b01100101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b11101010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b11110100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b01010110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b01101100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b10101001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b01001110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b11010101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b10001101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b01101101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b00110111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b11001000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b11100111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b01111001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b11100100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b10010101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b10010001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b01100010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b10101100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b11010011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b11000010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b01011100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b00100100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b00000110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b01001001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b00001010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b00111010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b00110010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b11100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b11011011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b00001011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b01011110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b11011110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b00010100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b10111000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b11101110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b01000110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b10001000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b10010000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b00101010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b00100010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b11011100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b01001111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b10000001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b01100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b01110011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b00011001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b01011101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b01100100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b00111101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b01111110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b10100111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b11000100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b00010111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b01000100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b10010111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b01011111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b11101100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b00010011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b00001100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b11001101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b11010010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b11110011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b11111111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b00010000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b00100001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b11011010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b10110110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b10111100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b11110101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b00111000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b10011101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b10010010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b10001111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b01000000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b10100011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b01010001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b10101000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b10011111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b00111100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b01010000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b01111111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b00000010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b11111001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b01000101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b10000101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b00110011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b01001101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b01000011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b11111011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b10101010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b11101111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b11010000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b11001111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b01011000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b01001100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b01001010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b00111001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b10111110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b11001011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b01101010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b01011011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b10110001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b11111100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b00100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b11101101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b00000000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b11010001 ;
      256'b????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b01010011 ;
      256'b???????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b10000100 ;
      256'b??????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b00101111 ;
      256'b?????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b11100011 ;
      256'b????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b00101001 ;
      256'b???????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b10110011 ;
      256'b??????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b11010110 ;
      256'b?????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b00111011 ;
      256'b????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b01010010 ;
      256'b???????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b10100000 ;
      256'b??????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b01011010 ;
      256'b?????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b01101110 ;
      256'b????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b00011011 ;
      256'b???????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b00011010 ;
      256'b??????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b00101100 ;
      256'b?????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b10000011 ;
      256'b????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b00001001 ;
      256'b???????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b01110101 ;
      256'b??????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b10110010 ;
      256'b?????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b00100111 ;
      256'b????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b11101011 ;
      256'b???????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b11100010 ;
      256'b??????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b10000000 ;
      256'b?????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b00010010 ;
      256'b????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b00000111 ;
      256'b???????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b10011010 ;
      256'b??????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b00000101 ;
      256'b?????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b10010110 ;
      256'b????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b00011000 ;
      256'b???????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b11000011 ;
      256'b??????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b00100011 ;
      256'b?????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b11000111 ;
      256'b????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b00000100 ;
      256'b???????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b00010101 ;
      256'b??????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b00110001 ;
      256'b?????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b11011000 ;
      256'b????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b01110001 ;
      256'b???????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b11110001 ;
      256'b??????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b11100101 ;
      256'b?????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b10100101 ;
      256'b????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b00110100 ;
      256'b???????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b11001100 ;
      256'b??????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b11110111 ;
      256'b?????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b00111111 ;
      256'b????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b00110110 ;
      256'b???????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b00100110 ;
      256'b??????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b10010011 ;
      256'b?????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b11111101 ;
      256'b????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b10110111 ;
      256'b???????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b11000000 ;
      256'b??????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b01110010 ;
      256'b?????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b10100100 ;
      256'b????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b10011100 ;
      256'b???????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b10101111 ;
      256'b??????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b10100010 ;
      256'b?????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b11010100 ;
      256'b????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b10101101 ;
      256'b???????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b11110000 ;
      256'b??????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b01000111 ;
      256'b?????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b01011001 ;
      256'b????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b11111010 ;
      256'b???????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b01111101 ;
      256'b??????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b11001001 ;
      256'b?????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b10000010 ;
      256'b????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b11001010 ;
      256'b???????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b01110110 ;
      256'b??????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b10101011 ;
      256'b?????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b11010111 ;
      256'b????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b11111110 ;
      256'b???????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b00101011 ;
      256'b??????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b01100111 ;
      256'b?????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b00000001 ;
      256'b????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b00110000 ;
      256'b???????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b11000101 ;
      256'b??????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b01101111 ;
      256'b?????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b01101011 ;
      256'b????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b11110010 ;
      256'b???1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b01111011 ;
      256'b??1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b01110111 ;
      256'b?1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b01111100 ;
      256'b1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b01100011 ;
      default:
        _3096_ = \t3.t0.s0.out ;
    endcase
  end
  assign _3097_ = state_in[31:24] == 8'b11111111;
  assign _3098_ = state_in[31:24] == 8'b11111110;
  assign _3099_ = state_in[31:24] == 8'b11111101;
  assign _3100_ = state_in[31:24] == 8'b11111100;
  assign _3101_ = state_in[31:24] == 8'b11111011;
  assign _3102_ = state_in[31:24] == 8'b11111010;
  assign _3103_ = state_in[31:24] == 8'b11111001;
  assign _3104_ = state_in[31:24] == 8'b11111000;
  assign _3105_ = state_in[31:24] == 8'b11110111;
  assign _3106_ = state_in[31:24] == 8'b11110110;
  assign _3107_ = state_in[31:24] == 8'b11110101;
  assign _3108_ = state_in[31:24] == 8'b11110100;
  assign _3109_ = state_in[31:24] == 8'b11110011;
  assign _3110_ = state_in[31:24] == 8'b11110010;
  assign _3111_ = state_in[31:24] == 8'b11110001;
  assign _3112_ = state_in[31:24] == 8'b11110000;
  assign _3113_ = state_in[31:24] == 8'b11101111;
  assign _3114_ = state_in[31:24] == 8'b11101110;
  assign _3115_ = state_in[31:24] == 8'b11101101;
  assign _3116_ = state_in[31:24] == 8'b11101100;
  assign _3117_ = state_in[31:24] == 8'b11101011;
  assign _3118_ = state_in[31:24] == 8'b11101010;
  assign _3119_ = state_in[31:24] == 8'b11101001;
  assign _3120_ = state_in[31:24] == 8'b11101000;
  assign _3121_ = state_in[31:24] == 8'b11100111;
  assign _3122_ = state_in[31:24] == 8'b11100110;
  assign _3123_ = state_in[31:24] == 8'b11100101;
  assign _3124_ = state_in[31:24] == 8'b11100100;
  assign _3125_ = state_in[31:24] == 8'b11100011;
  assign _3126_ = state_in[31:24] == 8'b11100010;
  assign _3127_ = state_in[31:24] == 8'b11100001;
  assign _3128_ = state_in[31:24] == 8'b11100000;
  assign _3129_ = state_in[31:24] == 8'b11011111;
  assign _3130_ = state_in[31:24] == 8'b11011110;
  assign _3131_ = state_in[31:24] == 8'b11011101;
  assign _3132_ = state_in[31:24] == 8'b11011100;
  assign _3133_ = state_in[31:24] == 8'b11011011;
  assign _3134_ = state_in[31:24] == 8'b11011010;
  assign _3135_ = state_in[31:24] == 8'b11011001;
  assign _3136_ = state_in[31:24] == 8'b11011000;
  assign _3137_ = state_in[31:24] == 8'b11010111;
  assign _3138_ = state_in[31:24] == 8'b11010110;
  assign _3139_ = state_in[31:24] == 8'b11010101;
  assign _3140_ = state_in[31:24] == 8'b11010100;
  assign _3141_ = state_in[31:24] == 8'b11010011;
  assign _3142_ = state_in[31:24] == 8'b11010010;
  assign _3143_ = state_in[31:24] == 8'b11010001;
  assign _3144_ = state_in[31:24] == 8'b11010000;
  assign _3145_ = state_in[31:24] == 8'b11001111;
  assign _3146_ = state_in[31:24] == 8'b11001110;
  assign _3147_ = state_in[31:24] == 8'b11001101;
  assign _3148_ = state_in[31:24] == 8'b11001100;
  assign _3149_ = state_in[31:24] == 8'b11001011;
  assign _3150_ = state_in[31:24] == 8'b11001010;
  assign _3151_ = state_in[31:24] == 8'b11001001;
  assign _3152_ = state_in[31:24] == 8'b11001000;
  assign _3153_ = state_in[31:24] == 8'b11000111;
  assign _3154_ = state_in[31:24] == 8'b11000110;
  assign _3155_ = state_in[31:24] == 8'b11000101;
  assign _3156_ = state_in[31:24] == 8'b11000100;
  assign _3157_ = state_in[31:24] == 8'b11000011;
  assign _3158_ = state_in[31:24] == 8'b11000010;
  assign _3159_ = state_in[31:24] == 8'b11000001;
  assign _3160_ = state_in[31:24] == 8'b11000000;
  assign _3161_ = state_in[31:24] == 8'b10111111;
  assign _3162_ = state_in[31:24] == 8'b10111110;
  assign _3163_ = state_in[31:24] == 8'b10111101;
  assign _3164_ = state_in[31:24] == 8'b10111100;
  assign _3165_ = state_in[31:24] == 8'b10111011;
  assign _3166_ = state_in[31:24] == 8'b10111010;
  assign _3167_ = state_in[31:24] == 8'b10111001;
  assign _3168_ = state_in[31:24] == 8'b10111000;
  assign _3169_ = state_in[31:24] == 8'b10110111;
  assign _3170_ = state_in[31:24] == 8'b10110110;
  assign _3171_ = state_in[31:24] == 8'b10110101;
  assign _3172_ = state_in[31:24] == 8'b10110100;
  assign _3173_ = state_in[31:24] == 8'b10110011;
  assign _3174_ = state_in[31:24] == 8'b10110010;
  assign _3175_ = state_in[31:24] == 8'b10110001;
  assign _3176_ = state_in[31:24] == 8'b10110000;
  assign _3177_ = state_in[31:24] == 8'b10101111;
  assign _3178_ = state_in[31:24] == 8'b10101110;
  assign _3179_ = state_in[31:24] == 8'b10101101;
  assign _3180_ = state_in[31:24] == 8'b10101100;
  assign _3181_ = state_in[31:24] == 8'b10101011;
  assign _3182_ = state_in[31:24] == 8'b10101010;
  assign _3183_ = state_in[31:24] == 8'b10101001;
  assign _3184_ = state_in[31:24] == 8'b10101000;
  assign _3185_ = state_in[31:24] == 8'b10100111;
  assign _3186_ = state_in[31:24] == 8'b10100110;
  assign _3187_ = state_in[31:24] == 8'b10100101;
  assign _3188_ = state_in[31:24] == 8'b10100100;
  assign _3189_ = state_in[31:24] == 8'b10100011;
  assign _3190_ = state_in[31:24] == 8'b10100010;
  assign _3191_ = state_in[31:24] == 8'b10100001;
  assign _3192_ = state_in[31:24] == 8'b10100000;
  assign _3193_ = state_in[31:24] == 8'b10011111;
  assign _3194_ = state_in[31:24] == 8'b10011110;
  assign _3195_ = state_in[31:24] == 8'b10011101;
  assign _3196_ = state_in[31:24] == 8'b10011100;
  assign _3197_ = state_in[31:24] == 8'b10011011;
  assign _3198_ = state_in[31:24] == 8'b10011010;
  assign _3199_ = state_in[31:24] == 8'b10011001;
  assign _3200_ = state_in[31:24] == 8'b10011000;
  assign _3201_ = state_in[31:24] == 8'b10010111;
  assign _3202_ = state_in[31:24] == 8'b10010110;
  assign _3203_ = state_in[31:24] == 8'b10010101;
  assign _3204_ = state_in[31:24] == 8'b10010100;
  assign _3205_ = state_in[31:24] == 8'b10010011;
  assign _3206_ = state_in[31:24] == 8'b10010010;
  assign _3207_ = state_in[31:24] == 8'b10010001;
  assign _3208_ = state_in[31:24] == 8'b10010000;
  assign _3209_ = state_in[31:24] == 8'b10001111;
  assign _3210_ = state_in[31:24] == 8'b10001110;
  assign _3211_ = state_in[31:24] == 8'b10001101;
  assign _3212_ = state_in[31:24] == 8'b10001100;
  assign _3213_ = state_in[31:24] == 8'b10001011;
  assign _3214_ = state_in[31:24] == 8'b10001010;
  assign _3215_ = state_in[31:24] == 8'b10001001;
  assign _3216_ = state_in[31:24] == 8'b10001000;
  assign _3217_ = state_in[31:24] == 8'b10000111;
  assign _3218_ = state_in[31:24] == 8'b10000110;
  assign _3219_ = state_in[31:24] == 8'b10000101;
  assign _3220_ = state_in[31:24] == 8'b10000100;
  assign _3221_ = state_in[31:24] == 8'b10000011;
  assign _3222_ = state_in[31:24] == 8'b10000010;
  assign _3223_ = state_in[31:24] == 8'b10000001;
  assign _3224_ = state_in[31:24] == 8'b10000000;
  assign _3225_ = state_in[31:24] == 7'b1111111;
  assign _3226_ = state_in[31:24] == 7'b1111110;
  assign _3227_ = state_in[31:24] == 7'b1111101;
  assign _3228_ = state_in[31:24] == 7'b1111100;
  assign _3229_ = state_in[31:24] == 7'b1111011;
  assign _3230_ = state_in[31:24] == 7'b1111010;
  assign _3231_ = state_in[31:24] == 7'b1111001;
  assign _3232_ = state_in[31:24] == 7'b1111000;
  assign _3233_ = state_in[31:24] == 7'b1110111;
  assign _3234_ = state_in[31:24] == 7'b1110110;
  assign _3235_ = state_in[31:24] == 7'b1110101;
  assign _3236_ = state_in[31:24] == 7'b1110100;
  assign _3237_ = state_in[31:24] == 7'b1110011;
  assign _3238_ = state_in[31:24] == 7'b1110010;
  assign _3239_ = state_in[31:24] == 7'b1110001;
  assign _3240_ = state_in[31:24] == 7'b1110000;
  assign _3241_ = state_in[31:24] == 7'b1101111;
  assign _3242_ = state_in[31:24] == 7'b1101110;
  assign _3243_ = state_in[31:24] == 7'b1101101;
  assign _3244_ = state_in[31:24] == 7'b1101100;
  assign _3245_ = state_in[31:24] == 7'b1101011;
  assign _3246_ = state_in[31:24] == 7'b1101010;
  assign _3247_ = state_in[31:24] == 7'b1101001;
  assign _3248_ = state_in[31:24] == 7'b1101000;
  assign _3249_ = state_in[31:24] == 7'b1100111;
  assign _3250_ = state_in[31:24] == 7'b1100110;
  assign _3251_ = state_in[31:24] == 7'b1100101;
  assign _3252_ = state_in[31:24] == 7'b1100100;
  assign _3253_ = state_in[31:24] == 7'b1100011;
  assign _3254_ = state_in[31:24] == 7'b1100010;
  assign _3255_ = state_in[31:24] == 7'b1100001;
  assign _3256_ = state_in[31:24] == 7'b1100000;
  assign _3257_ = state_in[31:24] == 7'b1011111;
  assign _3258_ = state_in[31:24] == 7'b1011110;
  assign _3259_ = state_in[31:24] == 7'b1011101;
  assign _3260_ = state_in[31:24] == 7'b1011100;
  assign _3261_ = state_in[31:24] == 7'b1011011;
  assign _3262_ = state_in[31:24] == 7'b1011010;
  assign _3263_ = state_in[31:24] == 7'b1011001;
  assign _3264_ = state_in[31:24] == 7'b1011000;
  assign _3265_ = state_in[31:24] == 7'b1010111;
  assign _3266_ = state_in[31:24] == 7'b1010110;
  assign _3267_ = state_in[31:24] == 7'b1010101;
  assign _3268_ = state_in[31:24] == 7'b1010100;
  assign _3269_ = state_in[31:24] == 7'b1010011;
  assign _3270_ = state_in[31:24] == 7'b1010010;
  assign _3271_ = state_in[31:24] == 7'b1010001;
  assign _3272_ = state_in[31:24] == 7'b1010000;
  assign _3273_ = state_in[31:24] == 7'b1001111;
  assign _3274_ = state_in[31:24] == 7'b1001110;
  assign _3275_ = state_in[31:24] == 7'b1001101;
  assign _3276_ = state_in[31:24] == 7'b1001100;
  assign _3277_ = state_in[31:24] == 7'b1001011;
  assign _3278_ = state_in[31:24] == 7'b1001010;
  assign _3279_ = state_in[31:24] == 7'b1001001;
  assign _3280_ = state_in[31:24] == 7'b1001000;
  assign _3281_ = state_in[31:24] == 7'b1000111;
  assign _3282_ = state_in[31:24] == 7'b1000110;
  assign _3283_ = state_in[31:24] == 7'b1000101;
  assign _3284_ = state_in[31:24] == 7'b1000100;
  assign _3285_ = state_in[31:24] == 7'b1000011;
  assign _3286_ = state_in[31:24] == 7'b1000010;
  assign _3287_ = state_in[31:24] == 7'b1000001;
  assign _3288_ = state_in[31:24] == 7'b1000000;
  assign _3289_ = state_in[31:24] == 6'b111111;
  assign _3290_ = state_in[31:24] == 6'b111110;
  assign _3291_ = state_in[31:24] == 6'b111101;
  assign _3292_ = state_in[31:24] == 6'b111100;
  assign _3293_ = state_in[31:24] == 6'b111011;
  assign _3294_ = state_in[31:24] == 6'b111010;
  assign _3295_ = state_in[31:24] == 6'b111001;
  assign _3296_ = state_in[31:24] == 6'b111000;
  assign _3297_ = state_in[31:24] == 6'b110111;
  assign _3298_ = state_in[31:24] == 6'b110110;
  assign _3299_ = state_in[31:24] == 6'b110101;
  assign _3300_ = state_in[31:24] == 6'b110100;
  assign _3301_ = state_in[31:24] == 6'b110011;
  assign _3302_ = state_in[31:24] == 6'b110010;
  assign _3303_ = state_in[31:24] == 6'b110001;
  assign _3304_ = state_in[31:24] == 6'b110000;
  assign _3305_ = state_in[31:24] == 6'b101111;
  assign _3306_ = state_in[31:24] == 6'b101110;
  assign _3307_ = state_in[31:24] == 6'b101101;
  assign _3308_ = state_in[31:24] == 6'b101100;
  assign _3309_ = state_in[31:24] == 6'b101011;
  assign _3310_ = state_in[31:24] == 6'b101010;
  assign _3311_ = state_in[31:24] == 6'b101001;
  assign _3312_ = state_in[31:24] == 6'b101000;
  assign _3313_ = state_in[31:24] == 6'b100111;
  assign _3314_ = state_in[31:24] == 6'b100110;
  assign _3315_ = state_in[31:24] == 6'b100101;
  assign _3316_ = state_in[31:24] == 6'b100100;
  assign _3317_ = state_in[31:24] == 6'b100011;
  assign _3318_ = state_in[31:24] == 6'b100010;
  assign _3319_ = state_in[31:24] == 6'b100001;
  assign _3320_ = state_in[31:24] == 6'b100000;
  assign _3321_ = state_in[31:24] == 5'b11111;
  assign _3322_ = state_in[31:24] == 5'b11110;
  assign _3323_ = state_in[31:24] == 5'b11101;
  assign _3324_ = state_in[31:24] == 5'b11100;
  assign _3325_ = state_in[31:24] == 5'b11011;
  assign _3326_ = state_in[31:24] == 5'b11010;
  assign _3327_ = state_in[31:24] == 5'b11001;
  assign _3328_ = state_in[31:24] == 5'b11000;
  assign _3329_ = state_in[31:24] == 5'b10111;
  assign _3330_ = state_in[31:24] == 5'b10110;
  assign _3331_ = state_in[31:24] == 5'b10101;
  assign _3332_ = state_in[31:24] == 5'b10100;
  assign _3333_ = state_in[31:24] == 5'b10011;
  assign _3334_ = state_in[31:24] == 5'b10010;
  assign _3335_ = state_in[31:24] == 5'b10001;
  assign _3336_ = state_in[31:24] == 5'b10000;
  assign _3337_ = state_in[31:24] == 4'b1111;
  assign _3338_ = state_in[31:24] == 4'b1110;
  assign _3339_ = state_in[31:24] == 4'b1101;
  assign _3340_ = state_in[31:24] == 4'b1100;
  assign _3341_ = state_in[31:24] == 4'b1011;
  assign _3342_ = state_in[31:24] == 4'b1010;
  assign _3343_ = state_in[31:24] == 4'b1001;
  assign _3344_ = state_in[31:24] == 4'b1000;
  assign _3345_ = state_in[31:24] == 3'b111;
  assign _3346_ = state_in[31:24] == 3'b110;
  assign _3347_ = state_in[31:24] == 3'b101;
  assign _3348_ = state_in[31:24] == 3'b100;
  assign _3349_ = state_in[31:24] == 2'b11;
  assign _3350_ = state_in[31:24] == 2'b10;
  assign _3351_ = state_in[31:24] == 1'b1;
  assign _3352_ = ! state_in[31:24];
  always @(posedge clk)
      \t3.t0.s4.out <= _3353_;
  wire [255:0] fangyuan26;
  assign fangyuan26 = { _3352_, _3351_, _3350_, _3349_, _3348_, _3347_, _3346_, _3345_, _3344_, _3343_, _3342_, _3341_, _3340_, _3339_, _3338_, _3337_, _3336_, _3335_, _3334_, _3333_, _3332_, _3331_, _3330_, _3329_, _3328_, _3327_, _3326_, _3325_, _3324_, _3323_, _3322_, _3321_, _3320_, _3319_, _3318_, _3317_, _3316_, _3315_, _3314_, _3313_, _3312_, _3311_, _3310_, _3309_, _3308_, _3307_, _3306_, _3305_, _3304_, _3303_, _3302_, _3301_, _3300_, _3299_, _3298_, _3297_, _3296_, _3295_, _3294_, _3293_, _3292_, _3291_, _3290_, _3289_, _3288_, _3287_, _3286_, _3285_, _3284_, _3283_, _3282_, _3281_, _3280_, _3279_, _3278_, _3277_, _3276_, _3275_, _3274_, _3273_, _3272_, _3271_, _3270_, _3269_, _3268_, _3267_, _3266_, _3265_, _3264_, _3263_, _3262_, _3261_, _3260_, _3259_, _3258_, _3257_, _3256_, _3255_, _3254_, _3253_, _3252_, _3251_, _3250_, _3249_, _3248_, _3247_, _3246_, _3245_, _3244_, _3243_, _3242_, _3241_, _3240_, _3239_, _3238_, _3237_, _3236_, _3235_, _3234_, _3233_, _3232_, _3231_, _3230_, _3229_, _3228_, _3227_, _3226_, _3225_, _3224_, _3223_, _3222_, _3221_, _3220_, _3219_, _3218_, _3217_, _3216_, _3215_, _3214_, _3213_, _3212_, _3211_, _3210_, _3209_, _3208_, _3207_, _3206_, _3205_, _3204_, _3203_, _3202_, _3201_, _3200_, _3199_, _3198_, _3197_, _3196_, _3195_, _3194_, _3193_, _3192_, _3191_, _3190_, _3189_, _3188_, _3187_, _3186_, _3185_, _3184_, _3183_, _3182_, _3181_, _3180_, _3179_, _3178_, _3177_, _3176_, _3175_, _3174_, _3173_, _3172_, _3171_, _3170_, _3169_, _3168_, _3167_, _3166_, _3165_, _3164_, _3163_, _3162_, _3161_, _3160_, _3159_, _3158_, _3157_, _3156_, _3155_, _3154_, _3153_, _3152_, _3151_, _3150_, _3149_, _3148_, _3147_, _3146_, _3145_, _3144_, _3143_, _3142_, _3141_, _3140_, _3139_, _3138_, _3137_, _3136_, _3135_, _3134_, _3133_, _3132_, _3131_, _3130_, _3129_, _3128_, _3127_, _3126_, _3125_, _3124_, _3123_, _3122_, _3121_, _3120_, _3119_, _3118_, _3117_, _3116_, _3115_, _3114_, _3113_, _3112_, _3111_, _3110_, _3109_, _3108_, _3107_, _3106_, _3105_, _3104_, _3103_, _3102_, _3101_, _3100_, _3099_, _3098_, _3097_ };

  always @(\t3.t0.s4.out or fangyuan26) begin
    casez (fangyuan26)
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1 :
        _3353_ = 8'b00101100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1? :
        _3353_ = 8'b01101101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?? :
        _3353_ = 8'b10101000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??? :
        _3353_ = 8'b01111011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???? :
        _3353_ = 8'b00011110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????? :
        _3353_ = 8'b01011010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????? :
        _3353_ = 8'b00101001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????? :
        _3353_ = 8'b10000010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????? :
        _3353_ = 8'b11010000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????? :
        _3353_ = 8'b10000100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????? :
        _3353_ = 8'b11010111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????? :
        _3353_ = 8'b01100101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????? :
        _3353_ = 8'b00011010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????? :
        _3353_ = 8'b00001001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????? :
        _3353_ = 8'b01011001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????? :
        _3353_ = 8'b00000011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????? :
        _3353_ = 8'b10100101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????? :
        _3353_ = 8'b01010000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????? :
        _3353_ = 8'b10101010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????? :
        _3353_ = 8'b10000111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????? :
        _3353_ = 8'b11001001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????? :
        _3353_ = 8'b00010101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????? :
        _3353_ = 8'b00111100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????? :
        _3353_ = 8'b00101101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????? :
        _3353_ = 8'b00110011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????? :
        _3353_ = 8'b00000111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????? :
        _3353_ = 8'b10101001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????? :
        _3353_ = 8'b11010010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????? :
        _3353_ = 8'b00100010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????? :
        _3353_ = 8'b00101011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????? :
        _3353_ = 8'b11101011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????? :
        _3353_ = 8'b11011001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????? :
        _3353_ = 8'b00100111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????? :
        _3353_ = 8'b00111010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????? :
        _3353_ = 8'b10011001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????? :
        _3353_ = 8'b00010111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????? :
        _3353_ = 8'b01101001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????? :
        _3353_ = 8'b10101110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????? :
        _3353_ = 8'b01101010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????? :
        _3353_ = 8'b11000010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????? :
        _3353_ = 8'b00011100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????? :
        _3353_ = 8'b11110111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????? :
        _3353_ = 8'b00000110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????? :
        _3353_ = 8'b10010000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????? :
        _3353_ = 8'b11001100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????? :
        _3353_ = 8'b01110001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????? :
        _3353_ = 8'b01111100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????? :
        _3353_ = 8'b11100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????? :
        _3353_ = 8'b00001111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????? :
        _3353_ = 8'b00001101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????? :
        _3353_ = 8'b01100001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????? :
        _3353_ = 8'b10010110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????? :
        _3353_ = 8'b00111110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????? :
        _3353_ = 8'b11101000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????? :
        _3353_ = 8'b10100001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????? :
        _3353_ = 8'b11001011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????? :
        _3353_ = 8'b10010111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????? :
        _3353_ = 8'b01110011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????? :
        _3353_ = 8'b01010111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????? :
        _3353_ = 8'b00111000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????? :
        _3353_ = 8'b01011100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????? :
        _3353_ = 8'b01001010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????? :
        _3353_ = 8'b11110000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????? :
        _3353_ = 8'b01101111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????? :
        _3353_ = 8'b00010000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b01000111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b11110100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b11001010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b11001111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b11110011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b10101100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b11011000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b01001001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b10011100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b10110001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b00000001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b11011010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b01101110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b10001011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b11010101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b11110010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b11010011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b00110001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b00111001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b11000100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b01000011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b10111101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b10011111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b10111000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b01001000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b00001100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b10010010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b00010100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b01110100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b01100100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b11011011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b10101101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b00010110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b10111100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b10100111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b00101000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b01101011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b11000111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b10001100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b00001011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b00111011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b01010100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b01000100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b10100011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b10011110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b00011001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b11000000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b11100110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b00110010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b10111010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b11001000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b01111010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b11111100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b01010101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b10010011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b00101110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b10001000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b00110101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b10111110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b11000011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b00100110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b00011000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b10000001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b10111111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b11111101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b11100101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b00100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b01000010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b10101111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b01110111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b01100011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b11110001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b01110000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b00100001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b00111111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b00000101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b10000000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b01011101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b10100010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b01001011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b00100101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b01111000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b10100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b11111110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b00000100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b11101001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b10001010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b00010001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b01100110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b10011010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b10000110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b11101101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b01001111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b11000101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b10111011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b10000101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b10110000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b10011000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b10010100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b01110010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b01100111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b10001101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b11010100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b10110110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b01111001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b11100011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b01000000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b11000001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b00000000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b10111001 ;
      256'b????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b10100110 ;
      256'b???????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b00010011 ;
      256'b??????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b01011110 ;
      256'b?????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b11011101 ;
      256'b????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b01010010 ;
      256'b???????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b01111101 ;
      256'b??????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b10110111 ;
      256'b?????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b01110110 ;
      256'b????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b10100100 ;
      256'b???????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b01011011 ;
      256'b??????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b10110100 ;
      256'b?????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b11011100 ;
      256'b????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b00110110 ;
      256'b???????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b00110100 ;
      256'b??????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b01011000 ;
      256'b?????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b00011101 ;
      256'b????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b00010010 ;
      256'b???????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b11101010 ;
      256'b??????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b01111111 ;
      256'b?????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b01001110 ;
      256'b????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b11001101 ;
      256'b???????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b11011111 ;
      256'b??????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b00011011 ;
      256'b?????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b00100100 ;
      256'b????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b00001110 ;
      256'b???????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b00101111 ;
      256'b??????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b00001010 ;
      256'b?????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b00110111 ;
      256'b????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b00110000 ;
      256'b???????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b10011101 ;
      256'b??????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b01000110 ;
      256'b?????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b10010101 ;
      256'b????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b00001000 ;
      256'b???????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b00101010 ;
      256'b??????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b01100010 ;
      256'b?????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b10101011 ;
      256'b????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b11100010 ;
      256'b???????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b11111001 ;
      256'b??????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b11010001 ;
      256'b?????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b01010001 ;
      256'b????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b01101000 ;
      256'b???????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b10000011 ;
      256'b??????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b11110101 ;
      256'b?????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b01111110 ;
      256'b????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b01101100 ;
      256'b???????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b01001100 ;
      256'b??????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b00111101 ;
      256'b?????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b11100001 ;
      256'b????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b01110101 ;
      256'b???????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b10011011 ;
      256'b??????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b11100100 ;
      256'b?????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b01010011 ;
      256'b????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b00100011 ;
      256'b???????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b01000101 ;
      256'b??????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b01011111 ;
      256'b?????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b10110011 ;
      256'b????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b01000001 ;
      256'b???????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b11111011 ;
      256'b??????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b10001110 ;
      256'b?????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b10110010 ;
      256'b????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b11101111 ;
      256'b???????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b11111010 ;
      256'b??????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b10001001 ;
      256'b?????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b00011111 ;
      256'b????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b10001111 ;
      256'b???????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b11101100 ;
      256'b??????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b01001101 ;
      256'b?????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b10110101 ;
      256'b????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b11100111 ;
      256'b???????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b01010110 ;
      256'b??????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b11001110 ;
      256'b?????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b00000010 ;
      256'b????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b01100000 ;
      256'b???????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b10010001 ;
      256'b??????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b11011110 ;
      256'b?????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b11010110 ;
      256'b????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b11111111 ;
      256'b???1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b11110110 ;
      256'b??1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b11101110 ;
      256'b?1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b11111000 ;
      256'b1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b11000110 ;
      default:
        _3353_ = \t3.t0.s4.out ;
    endcase
  end
  assign p31[31:24] = \t3.t1.s0.out ^ \t3.t1.s4.out ;
  always @(posedge clk)
      \t3.t1.s0.out <= _3354_;
  wire [255:0] fangyuan27;
  assign fangyuan27 = { _3610_, _3609_, _3608_, _3607_, _3606_, _3605_, _3604_, _3603_, _3602_, _3601_, _3600_, _3599_, _3598_, _3597_, _3596_, _3595_, _3594_, _3593_, _3592_, _3591_, _3590_, _3589_, _3588_, _3587_, _3586_, _3585_, _3584_, _3583_, _3582_, _3581_, _3580_, _3579_, _3578_, _3577_, _3576_, _3575_, _3574_, _3573_, _3572_, _3571_, _3570_, _3569_, _3568_, _3567_, _3566_, _3565_, _3564_, _3563_, _3562_, _3561_, _3560_, _3559_, _3558_, _3557_, _3556_, _3555_, _3554_, _3553_, _3552_, _3551_, _3550_, _3549_, _3548_, _3547_, _3546_, _3545_, _3544_, _3543_, _3542_, _3541_, _3540_, _3539_, _3538_, _3537_, _3536_, _3535_, _3534_, _3533_, _3532_, _3531_, _3530_, _3529_, _3528_, _3527_, _3526_, _3525_, _3524_, _3523_, _3522_, _3521_, _3520_, _3519_, _3518_, _3517_, _3516_, _3515_, _3514_, _3513_, _3512_, _3511_, _3510_, _3509_, _3508_, _3507_, _3506_, _3505_, _3504_, _3503_, _3502_, _3501_, _3500_, _3499_, _3498_, _3497_, _3496_, _3495_, _3494_, _3493_, _3492_, _3491_, _3490_, _3489_, _3488_, _3487_, _3486_, _3485_, _3484_, _3483_, _3482_, _3481_, _3480_, _3479_, _3478_, _3477_, _3476_, _3475_, _3474_, _3473_, _3472_, _3471_, _3470_, _3469_, _3468_, _3467_, _3466_, _3465_, _3464_, _3463_, _3462_, _3461_, _3460_, _3459_, _3458_, _3457_, _3456_, _3455_, _3454_, _3453_, _3452_, _3451_, _3450_, _3449_, _3448_, _3447_, _3446_, _3445_, _3444_, _3443_, _3442_, _3441_, _3440_, _3439_, _3438_, _3437_, _3436_, _3435_, _3434_, _3433_, _3432_, _3431_, _3430_, _3429_, _3428_, _3427_, _3426_, _3425_, _3424_, _3423_, _3422_, _3421_, _3420_, _3419_, _3418_, _3417_, _3416_, _3415_, _3414_, _3413_, _3412_, _3411_, _3410_, _3409_, _3408_, _3407_, _3406_, _3405_, _3404_, _3403_, _3402_, _3401_, _3400_, _3399_, _3398_, _3397_, _3396_, _3395_, _3394_, _3393_, _3392_, _3391_, _3390_, _3389_, _3388_, _3387_, _3386_, _3385_, _3384_, _3383_, _3382_, _3381_, _3380_, _3379_, _3378_, _3377_, _3376_, _3375_, _3374_, _3373_, _3372_, _3371_, _3370_, _3369_, _3368_, _3367_, _3366_, _3365_, _3364_, _3363_, _3362_, _3361_, _3360_, _3359_, _3358_, _3357_, _3356_, _3355_ };

  always @(\t3.t1.s0.out or fangyuan27) begin
    casez (fangyuan27)
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1 :
        _3354_ = 8'b00010110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1? :
        _3354_ = 8'b10111011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?? :
        _3354_ = 8'b01010100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??? :
        _3354_ = 8'b10110000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???? :
        _3354_ = 8'b00001111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????? :
        _3354_ = 8'b00101101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????? :
        _3354_ = 8'b10011001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????? :
        _3354_ = 8'b01000001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????? :
        _3354_ = 8'b01101000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????? :
        _3354_ = 8'b01000010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????? :
        _3354_ = 8'b11100110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????? :
        _3354_ = 8'b10111111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????? :
        _3354_ = 8'b00001101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????? :
        _3354_ = 8'b10001001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????? :
        _3354_ = 8'b10100001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????? :
        _3354_ = 8'b10001100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????? :
        _3354_ = 8'b11011111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????? :
        _3354_ = 8'b00101000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????? :
        _3354_ = 8'b01010101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????? :
        _3354_ = 8'b11001110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????? :
        _3354_ = 8'b11101001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????? :
        _3354_ = 8'b10000111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????? :
        _3354_ = 8'b00011110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????? :
        _3354_ = 8'b10011011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????? :
        _3354_ = 8'b10010100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????? :
        _3354_ = 8'b10001110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????? :
        _3354_ = 8'b11011001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????? :
        _3354_ = 8'b01101001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????? :
        _3354_ = 8'b00010001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????? :
        _3354_ = 8'b10011000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????? :
        _3354_ = 8'b11111000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????? :
        _3354_ = 8'b11100001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????? :
        _3354_ = 8'b10011110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????? :
        _3354_ = 8'b00011101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????? :
        _3354_ = 8'b11000001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????? :
        _3354_ = 8'b10000110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????? :
        _3354_ = 8'b10111001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????? :
        _3354_ = 8'b01010111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????? :
        _3354_ = 8'b00110101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????? :
        _3354_ = 8'b01100001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????? :
        _3354_ = 8'b00001110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????? :
        _3354_ = 8'b11110110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????? :
        _3354_ = 8'b00000011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????? :
        _3354_ = 8'b01001000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????? :
        _3354_ = 8'b01100110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????? :
        _3354_ = 8'b10110101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????? :
        _3354_ = 8'b00111110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????? :
        _3354_ = 8'b01110000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????? :
        _3354_ = 8'b10001010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????? :
        _3354_ = 8'b10001011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????? :
        _3354_ = 8'b10111101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????? :
        _3354_ = 8'b01001011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????? :
        _3354_ = 8'b00011111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????? :
        _3354_ = 8'b01110100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????? :
        _3354_ = 8'b11011101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????? :
        _3354_ = 8'b11101000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????? :
        _3354_ = 8'b11000110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????? :
        _3354_ = 8'b10110100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????? :
        _3354_ = 8'b10100110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????? :
        _3354_ = 8'b00011100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????? :
        _3354_ = 8'b00101110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????? :
        _3354_ = 8'b00100101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????? :
        _3354_ = 8'b01111000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????? :
        _3354_ = 8'b10111010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????? :
        _3354_ = 8'b00001000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b10101110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b01111010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b01100101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b11101010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b11110100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b01010110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b01101100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b10101001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b01001110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b11010101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b10001101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b01101101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b00110111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b11001000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b11100111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b01111001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b11100100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b10010101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b10010001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b01100010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b10101100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b11010011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b11000010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b01011100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b00100100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b00000110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b01001001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b00001010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b00111010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b00110010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b11100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b11011011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b00001011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b01011110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b11011110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b00010100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b10111000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b11101110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b01000110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b10001000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b10010000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b00101010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b00100010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b11011100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b01001111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b10000001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b01100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b01110011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b00011001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b01011101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b01100100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b00111101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b01111110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b10100111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b11000100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b00010111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b01000100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b10010111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b01011111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b11101100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b00010011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b00001100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b11001101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b11010010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b11110011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b11111111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b00010000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b00100001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b11011010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b10110110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b10111100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b11110101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b00111000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b10011101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b10010010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b10001111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b01000000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b10100011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b01010001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b10101000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b10011111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b00111100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b01010000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b01111111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b00000010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b11111001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b01000101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b10000101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b00110011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b01001101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b01000011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b11111011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b10101010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b11101111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b11010000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b11001111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b01011000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b01001100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b01001010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b00111001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b10111110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b11001011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b01101010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b01011011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b10110001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b11111100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b00100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b11101101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b00000000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b11010001 ;
      256'b????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b01010011 ;
      256'b???????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b10000100 ;
      256'b??????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b00101111 ;
      256'b?????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b11100011 ;
      256'b????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b00101001 ;
      256'b???????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b10110011 ;
      256'b??????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b11010110 ;
      256'b?????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b00111011 ;
      256'b????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b01010010 ;
      256'b???????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b10100000 ;
      256'b??????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b01011010 ;
      256'b?????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b01101110 ;
      256'b????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b00011011 ;
      256'b???????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b00011010 ;
      256'b??????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b00101100 ;
      256'b?????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b10000011 ;
      256'b????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b00001001 ;
      256'b???????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b01110101 ;
      256'b??????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b10110010 ;
      256'b?????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b00100111 ;
      256'b????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b11101011 ;
      256'b???????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b11100010 ;
      256'b??????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b10000000 ;
      256'b?????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b00010010 ;
      256'b????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b00000111 ;
      256'b???????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b10011010 ;
      256'b??????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b00000101 ;
      256'b?????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b10010110 ;
      256'b????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b00011000 ;
      256'b???????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b11000011 ;
      256'b??????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b00100011 ;
      256'b?????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b11000111 ;
      256'b????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b00000100 ;
      256'b???????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b00010101 ;
      256'b??????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b00110001 ;
      256'b?????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b11011000 ;
      256'b????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b01110001 ;
      256'b???????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b11110001 ;
      256'b??????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b11100101 ;
      256'b?????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b10100101 ;
      256'b????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b00110100 ;
      256'b???????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b11001100 ;
      256'b??????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b11110111 ;
      256'b?????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b00111111 ;
      256'b????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b00110110 ;
      256'b???????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b00100110 ;
      256'b??????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b10010011 ;
      256'b?????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b11111101 ;
      256'b????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b10110111 ;
      256'b???????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b11000000 ;
      256'b??????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b01110010 ;
      256'b?????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b10100100 ;
      256'b????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b10011100 ;
      256'b???????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b10101111 ;
      256'b??????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b10100010 ;
      256'b?????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b11010100 ;
      256'b????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b10101101 ;
      256'b???????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b11110000 ;
      256'b??????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b01000111 ;
      256'b?????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b01011001 ;
      256'b????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b11111010 ;
      256'b???????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b01111101 ;
      256'b??????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b11001001 ;
      256'b?????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b10000010 ;
      256'b????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b11001010 ;
      256'b???????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b01110110 ;
      256'b??????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b10101011 ;
      256'b?????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b11010111 ;
      256'b????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b11111110 ;
      256'b???????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b00101011 ;
      256'b??????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b01100111 ;
      256'b?????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b00000001 ;
      256'b????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b00110000 ;
      256'b???????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b11000101 ;
      256'b??????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b01101111 ;
      256'b?????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b01101011 ;
      256'b????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b11110010 ;
      256'b???1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b01111011 ;
      256'b??1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b01110111 ;
      256'b?1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b01111100 ;
      256'b1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b01100011 ;
      default:
        _3354_ = \t3.t1.s0.out ;
    endcase
  end
  assign _3355_ = state_in[23:16] == 8'b11111111;
  assign _3356_ = state_in[23:16] == 8'b11111110;
  assign _3357_ = state_in[23:16] == 8'b11111101;
  assign _3358_ = state_in[23:16] == 8'b11111100;
  assign _3359_ = state_in[23:16] == 8'b11111011;
  assign _3360_ = state_in[23:16] == 8'b11111010;
  assign _3361_ = state_in[23:16] == 8'b11111001;
  assign _3362_ = state_in[23:16] == 8'b11111000;
  assign _3363_ = state_in[23:16] == 8'b11110111;
  assign _3364_ = state_in[23:16] == 8'b11110110;
  assign _3365_ = state_in[23:16] == 8'b11110101;
  assign _3366_ = state_in[23:16] == 8'b11110100;
  assign _3367_ = state_in[23:16] == 8'b11110011;
  assign _3368_ = state_in[23:16] == 8'b11110010;
  assign _3369_ = state_in[23:16] == 8'b11110001;
  assign _3370_ = state_in[23:16] == 8'b11110000;
  assign _3371_ = state_in[23:16] == 8'b11101111;
  assign _3372_ = state_in[23:16] == 8'b11101110;
  assign _3373_ = state_in[23:16] == 8'b11101101;
  assign _3374_ = state_in[23:16] == 8'b11101100;
  assign _3375_ = state_in[23:16] == 8'b11101011;
  assign _3376_ = state_in[23:16] == 8'b11101010;
  assign _3377_ = state_in[23:16] == 8'b11101001;
  assign _3378_ = state_in[23:16] == 8'b11101000;
  assign _3379_ = state_in[23:16] == 8'b11100111;
  assign _3380_ = state_in[23:16] == 8'b11100110;
  assign _3381_ = state_in[23:16] == 8'b11100101;
  assign _3382_ = state_in[23:16] == 8'b11100100;
  assign _3383_ = state_in[23:16] == 8'b11100011;
  assign _3384_ = state_in[23:16] == 8'b11100010;
  assign _3385_ = state_in[23:16] == 8'b11100001;
  assign _3386_ = state_in[23:16] == 8'b11100000;
  assign _3387_ = state_in[23:16] == 8'b11011111;
  assign _3388_ = state_in[23:16] == 8'b11011110;
  assign _3389_ = state_in[23:16] == 8'b11011101;
  assign _3390_ = state_in[23:16] == 8'b11011100;
  assign _3391_ = state_in[23:16] == 8'b11011011;
  assign _3392_ = state_in[23:16] == 8'b11011010;
  assign _3393_ = state_in[23:16] == 8'b11011001;
  assign _3394_ = state_in[23:16] == 8'b11011000;
  assign _3395_ = state_in[23:16] == 8'b11010111;
  assign _3396_ = state_in[23:16] == 8'b11010110;
  assign _3397_ = state_in[23:16] == 8'b11010101;
  assign _3398_ = state_in[23:16] == 8'b11010100;
  assign _3399_ = state_in[23:16] == 8'b11010011;
  assign _3400_ = state_in[23:16] == 8'b11010010;
  assign _3401_ = state_in[23:16] == 8'b11010001;
  assign _3402_ = state_in[23:16] == 8'b11010000;
  assign _3403_ = state_in[23:16] == 8'b11001111;
  assign _3404_ = state_in[23:16] == 8'b11001110;
  assign _3405_ = state_in[23:16] == 8'b11001101;
  assign _3406_ = state_in[23:16] == 8'b11001100;
  assign _3407_ = state_in[23:16] == 8'b11001011;
  assign _3408_ = state_in[23:16] == 8'b11001010;
  assign _3409_ = state_in[23:16] == 8'b11001001;
  assign _3410_ = state_in[23:16] == 8'b11001000;
  assign _3411_ = state_in[23:16] == 8'b11000111;
  assign _3412_ = state_in[23:16] == 8'b11000110;
  assign _3413_ = state_in[23:16] == 8'b11000101;
  assign _3414_ = state_in[23:16] == 8'b11000100;
  assign _3415_ = state_in[23:16] == 8'b11000011;
  assign _3416_ = state_in[23:16] == 8'b11000010;
  assign _3417_ = state_in[23:16] == 8'b11000001;
  assign _3418_ = state_in[23:16] == 8'b11000000;
  assign _3419_ = state_in[23:16] == 8'b10111111;
  assign _3420_ = state_in[23:16] == 8'b10111110;
  assign _3421_ = state_in[23:16] == 8'b10111101;
  assign _3422_ = state_in[23:16] == 8'b10111100;
  assign _3423_ = state_in[23:16] == 8'b10111011;
  assign _3424_ = state_in[23:16] == 8'b10111010;
  assign _3425_ = state_in[23:16] == 8'b10111001;
  assign _3426_ = state_in[23:16] == 8'b10111000;
  assign _3427_ = state_in[23:16] == 8'b10110111;
  assign _3428_ = state_in[23:16] == 8'b10110110;
  assign _3429_ = state_in[23:16] == 8'b10110101;
  assign _3430_ = state_in[23:16] == 8'b10110100;
  assign _3431_ = state_in[23:16] == 8'b10110011;
  assign _3432_ = state_in[23:16] == 8'b10110010;
  assign _3433_ = state_in[23:16] == 8'b10110001;
  assign _3434_ = state_in[23:16] == 8'b10110000;
  assign _3435_ = state_in[23:16] == 8'b10101111;
  assign _3436_ = state_in[23:16] == 8'b10101110;
  assign _3437_ = state_in[23:16] == 8'b10101101;
  assign _3438_ = state_in[23:16] == 8'b10101100;
  assign _3439_ = state_in[23:16] == 8'b10101011;
  assign _3440_ = state_in[23:16] == 8'b10101010;
  assign _3441_ = state_in[23:16] == 8'b10101001;
  assign _3442_ = state_in[23:16] == 8'b10101000;
  assign _3443_ = state_in[23:16] == 8'b10100111;
  assign _3444_ = state_in[23:16] == 8'b10100110;
  assign _3445_ = state_in[23:16] == 8'b10100101;
  assign _3446_ = state_in[23:16] == 8'b10100100;
  assign _3447_ = state_in[23:16] == 8'b10100011;
  assign _3448_ = state_in[23:16] == 8'b10100010;
  assign _3449_ = state_in[23:16] == 8'b10100001;
  assign _3450_ = state_in[23:16] == 8'b10100000;
  assign _3451_ = state_in[23:16] == 8'b10011111;
  assign _3452_ = state_in[23:16] == 8'b10011110;
  assign _3453_ = state_in[23:16] == 8'b10011101;
  assign _3454_ = state_in[23:16] == 8'b10011100;
  assign _3455_ = state_in[23:16] == 8'b10011011;
  assign _3456_ = state_in[23:16] == 8'b10011010;
  assign _3457_ = state_in[23:16] == 8'b10011001;
  assign _3458_ = state_in[23:16] == 8'b10011000;
  assign _3459_ = state_in[23:16] == 8'b10010111;
  assign _3460_ = state_in[23:16] == 8'b10010110;
  assign _3461_ = state_in[23:16] == 8'b10010101;
  assign _3462_ = state_in[23:16] == 8'b10010100;
  assign _3463_ = state_in[23:16] == 8'b10010011;
  assign _3464_ = state_in[23:16] == 8'b10010010;
  assign _3465_ = state_in[23:16] == 8'b10010001;
  assign _3466_ = state_in[23:16] == 8'b10010000;
  assign _3467_ = state_in[23:16] == 8'b10001111;
  assign _3468_ = state_in[23:16] == 8'b10001110;
  assign _3469_ = state_in[23:16] == 8'b10001101;
  assign _3470_ = state_in[23:16] == 8'b10001100;
  assign _3471_ = state_in[23:16] == 8'b10001011;
  assign _3472_ = state_in[23:16] == 8'b10001010;
  assign _3473_ = state_in[23:16] == 8'b10001001;
  assign _3474_ = state_in[23:16] == 8'b10001000;
  assign _3475_ = state_in[23:16] == 8'b10000111;
  assign _3476_ = state_in[23:16] == 8'b10000110;
  assign _3477_ = state_in[23:16] == 8'b10000101;
  assign _3478_ = state_in[23:16] == 8'b10000100;
  assign _3479_ = state_in[23:16] == 8'b10000011;
  assign _3480_ = state_in[23:16] == 8'b10000010;
  assign _3481_ = state_in[23:16] == 8'b10000001;
  assign _3482_ = state_in[23:16] == 8'b10000000;
  assign _3483_ = state_in[23:16] == 7'b1111111;
  assign _3484_ = state_in[23:16] == 7'b1111110;
  assign _3485_ = state_in[23:16] == 7'b1111101;
  assign _3486_ = state_in[23:16] == 7'b1111100;
  assign _3487_ = state_in[23:16] == 7'b1111011;
  assign _3488_ = state_in[23:16] == 7'b1111010;
  assign _3489_ = state_in[23:16] == 7'b1111001;
  assign _3490_ = state_in[23:16] == 7'b1111000;
  assign _3491_ = state_in[23:16] == 7'b1110111;
  assign _3492_ = state_in[23:16] == 7'b1110110;
  assign _3493_ = state_in[23:16] == 7'b1110101;
  assign _3494_ = state_in[23:16] == 7'b1110100;
  assign _3495_ = state_in[23:16] == 7'b1110011;
  assign _3496_ = state_in[23:16] == 7'b1110010;
  assign _3497_ = state_in[23:16] == 7'b1110001;
  assign _3498_ = state_in[23:16] == 7'b1110000;
  assign _3499_ = state_in[23:16] == 7'b1101111;
  assign _3500_ = state_in[23:16] == 7'b1101110;
  assign _3501_ = state_in[23:16] == 7'b1101101;
  assign _3502_ = state_in[23:16] == 7'b1101100;
  assign _3503_ = state_in[23:16] == 7'b1101011;
  assign _3504_ = state_in[23:16] == 7'b1101010;
  assign _3505_ = state_in[23:16] == 7'b1101001;
  assign _3506_ = state_in[23:16] == 7'b1101000;
  assign _3507_ = state_in[23:16] == 7'b1100111;
  assign _3508_ = state_in[23:16] == 7'b1100110;
  assign _3509_ = state_in[23:16] == 7'b1100101;
  assign _3510_ = state_in[23:16] == 7'b1100100;
  assign _3511_ = state_in[23:16] == 7'b1100011;
  assign _3512_ = state_in[23:16] == 7'b1100010;
  assign _3513_ = state_in[23:16] == 7'b1100001;
  assign _3514_ = state_in[23:16] == 7'b1100000;
  assign _3515_ = state_in[23:16] == 7'b1011111;
  assign _3516_ = state_in[23:16] == 7'b1011110;
  assign _3517_ = state_in[23:16] == 7'b1011101;
  assign _3518_ = state_in[23:16] == 7'b1011100;
  assign _3519_ = state_in[23:16] == 7'b1011011;
  assign _3520_ = state_in[23:16] == 7'b1011010;
  assign _3521_ = state_in[23:16] == 7'b1011001;
  assign _3522_ = state_in[23:16] == 7'b1011000;
  assign _3523_ = state_in[23:16] == 7'b1010111;
  assign _3524_ = state_in[23:16] == 7'b1010110;
  assign _3525_ = state_in[23:16] == 7'b1010101;
  assign _3526_ = state_in[23:16] == 7'b1010100;
  assign _3527_ = state_in[23:16] == 7'b1010011;
  assign _3528_ = state_in[23:16] == 7'b1010010;
  assign _3529_ = state_in[23:16] == 7'b1010001;
  assign _3530_ = state_in[23:16] == 7'b1010000;
  assign _3531_ = state_in[23:16] == 7'b1001111;
  assign _3532_ = state_in[23:16] == 7'b1001110;
  assign _3533_ = state_in[23:16] == 7'b1001101;
  assign _3534_ = state_in[23:16] == 7'b1001100;
  assign _3535_ = state_in[23:16] == 7'b1001011;
  assign _3536_ = state_in[23:16] == 7'b1001010;
  assign _3537_ = state_in[23:16] == 7'b1001001;
  assign _3538_ = state_in[23:16] == 7'b1001000;
  assign _3539_ = state_in[23:16] == 7'b1000111;
  assign _3540_ = state_in[23:16] == 7'b1000110;
  assign _3541_ = state_in[23:16] == 7'b1000101;
  assign _3542_ = state_in[23:16] == 7'b1000100;
  assign _3543_ = state_in[23:16] == 7'b1000011;
  assign _3544_ = state_in[23:16] == 7'b1000010;
  assign _3545_ = state_in[23:16] == 7'b1000001;
  assign _3546_ = state_in[23:16] == 7'b1000000;
  assign _3547_ = state_in[23:16] == 6'b111111;
  assign _3548_ = state_in[23:16] == 6'b111110;
  assign _3549_ = state_in[23:16] == 6'b111101;
  assign _3550_ = state_in[23:16] == 6'b111100;
  assign _3551_ = state_in[23:16] == 6'b111011;
  assign _3552_ = state_in[23:16] == 6'b111010;
  assign _3553_ = state_in[23:16] == 6'b111001;
  assign _3554_ = state_in[23:16] == 6'b111000;
  assign _3555_ = state_in[23:16] == 6'b110111;
  assign _3556_ = state_in[23:16] == 6'b110110;
  assign _3557_ = state_in[23:16] == 6'b110101;
  assign _3558_ = state_in[23:16] == 6'b110100;
  assign _3559_ = state_in[23:16] == 6'b110011;
  assign _3560_ = state_in[23:16] == 6'b110010;
  assign _3561_ = state_in[23:16] == 6'b110001;
  assign _3562_ = state_in[23:16] == 6'b110000;
  assign _3563_ = state_in[23:16] == 6'b101111;
  assign _3564_ = state_in[23:16] == 6'b101110;
  assign _3565_ = state_in[23:16] == 6'b101101;
  assign _3566_ = state_in[23:16] == 6'b101100;
  assign _3567_ = state_in[23:16] == 6'b101011;
  assign _3568_ = state_in[23:16] == 6'b101010;
  assign _3569_ = state_in[23:16] == 6'b101001;
  assign _3570_ = state_in[23:16] == 6'b101000;
  assign _3571_ = state_in[23:16] == 6'b100111;
  assign _3572_ = state_in[23:16] == 6'b100110;
  assign _3573_ = state_in[23:16] == 6'b100101;
  assign _3574_ = state_in[23:16] == 6'b100100;
  assign _3575_ = state_in[23:16] == 6'b100011;
  assign _3576_ = state_in[23:16] == 6'b100010;
  assign _3577_ = state_in[23:16] == 6'b100001;
  assign _3578_ = state_in[23:16] == 6'b100000;
  assign _3579_ = state_in[23:16] == 5'b11111;
  assign _3580_ = state_in[23:16] == 5'b11110;
  assign _3581_ = state_in[23:16] == 5'b11101;
  assign _3582_ = state_in[23:16] == 5'b11100;
  assign _3583_ = state_in[23:16] == 5'b11011;
  assign _3584_ = state_in[23:16] == 5'b11010;
  assign _3585_ = state_in[23:16] == 5'b11001;
  assign _3586_ = state_in[23:16] == 5'b11000;
  assign _3587_ = state_in[23:16] == 5'b10111;
  assign _3588_ = state_in[23:16] == 5'b10110;
  assign _3589_ = state_in[23:16] == 5'b10101;
  assign _3590_ = state_in[23:16] == 5'b10100;
  assign _3591_ = state_in[23:16] == 5'b10011;
  assign _3592_ = state_in[23:16] == 5'b10010;
  assign _3593_ = state_in[23:16] == 5'b10001;
  assign _3594_ = state_in[23:16] == 5'b10000;
  assign _3595_ = state_in[23:16] == 4'b1111;
  assign _3596_ = state_in[23:16] == 4'b1110;
  assign _3597_ = state_in[23:16] == 4'b1101;
  assign _3598_ = state_in[23:16] == 4'b1100;
  assign _3599_ = state_in[23:16] == 4'b1011;
  assign _3600_ = state_in[23:16] == 4'b1010;
  assign _3601_ = state_in[23:16] == 4'b1001;
  assign _3602_ = state_in[23:16] == 4'b1000;
  assign _3603_ = state_in[23:16] == 3'b111;
  assign _3604_ = state_in[23:16] == 3'b110;
  assign _3605_ = state_in[23:16] == 3'b101;
  assign _3606_ = state_in[23:16] == 3'b100;
  assign _3607_ = state_in[23:16] == 2'b11;
  assign _3608_ = state_in[23:16] == 2'b10;
  assign _3609_ = state_in[23:16] == 1'b1;
  assign _3610_ = ! state_in[23:16];
  always @(posedge clk)
      \t3.t1.s4.out <= _3611_;
  wire [255:0] fangyuan28;
  assign fangyuan28 = { _3610_, _3609_, _3608_, _3607_, _3606_, _3605_, _3604_, _3603_, _3602_, _3601_, _3600_, _3599_, _3598_, _3597_, _3596_, _3595_, _3594_, _3593_, _3592_, _3591_, _3590_, _3589_, _3588_, _3587_, _3586_, _3585_, _3584_, _3583_, _3582_, _3581_, _3580_, _3579_, _3578_, _3577_, _3576_, _3575_, _3574_, _3573_, _3572_, _3571_, _3570_, _3569_, _3568_, _3567_, _3566_, _3565_, _3564_, _3563_, _3562_, _3561_, _3560_, _3559_, _3558_, _3557_, _3556_, _3555_, _3554_, _3553_, _3552_, _3551_, _3550_, _3549_, _3548_, _3547_, _3546_, _3545_, _3544_, _3543_, _3542_, _3541_, _3540_, _3539_, _3538_, _3537_, _3536_, _3535_, _3534_, _3533_, _3532_, _3531_, _3530_, _3529_, _3528_, _3527_, _3526_, _3525_, _3524_, _3523_, _3522_, _3521_, _3520_, _3519_, _3518_, _3517_, _3516_, _3515_, _3514_, _3513_, _3512_, _3511_, _3510_, _3509_, _3508_, _3507_, _3506_, _3505_, _3504_, _3503_, _3502_, _3501_, _3500_, _3499_, _3498_, _3497_, _3496_, _3495_, _3494_, _3493_, _3492_, _3491_, _3490_, _3489_, _3488_, _3487_, _3486_, _3485_, _3484_, _3483_, _3482_, _3481_, _3480_, _3479_, _3478_, _3477_, _3476_, _3475_, _3474_, _3473_, _3472_, _3471_, _3470_, _3469_, _3468_, _3467_, _3466_, _3465_, _3464_, _3463_, _3462_, _3461_, _3460_, _3459_, _3458_, _3457_, _3456_, _3455_, _3454_, _3453_, _3452_, _3451_, _3450_, _3449_, _3448_, _3447_, _3446_, _3445_, _3444_, _3443_, _3442_, _3441_, _3440_, _3439_, _3438_, _3437_, _3436_, _3435_, _3434_, _3433_, _3432_, _3431_, _3430_, _3429_, _3428_, _3427_, _3426_, _3425_, _3424_, _3423_, _3422_, _3421_, _3420_, _3419_, _3418_, _3417_, _3416_, _3415_, _3414_, _3413_, _3412_, _3411_, _3410_, _3409_, _3408_, _3407_, _3406_, _3405_, _3404_, _3403_, _3402_, _3401_, _3400_, _3399_, _3398_, _3397_, _3396_, _3395_, _3394_, _3393_, _3392_, _3391_, _3390_, _3389_, _3388_, _3387_, _3386_, _3385_, _3384_, _3383_, _3382_, _3381_, _3380_, _3379_, _3378_, _3377_, _3376_, _3375_, _3374_, _3373_, _3372_, _3371_, _3370_, _3369_, _3368_, _3367_, _3366_, _3365_, _3364_, _3363_, _3362_, _3361_, _3360_, _3359_, _3358_, _3357_, _3356_, _3355_ };

  always @(\t3.t1.s4.out or fangyuan28) begin
    casez (fangyuan28)
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1 :
        _3611_ = 8'b00101100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1? :
        _3611_ = 8'b01101101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?? :
        _3611_ = 8'b10101000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??? :
        _3611_ = 8'b01111011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???? :
        _3611_ = 8'b00011110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????? :
        _3611_ = 8'b01011010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????? :
        _3611_ = 8'b00101001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????? :
        _3611_ = 8'b10000010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????? :
        _3611_ = 8'b11010000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????? :
        _3611_ = 8'b10000100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????? :
        _3611_ = 8'b11010111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????? :
        _3611_ = 8'b01100101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????? :
        _3611_ = 8'b00011010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????? :
        _3611_ = 8'b00001001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????? :
        _3611_ = 8'b01011001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????? :
        _3611_ = 8'b00000011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????? :
        _3611_ = 8'b10100101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????? :
        _3611_ = 8'b01010000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????? :
        _3611_ = 8'b10101010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????? :
        _3611_ = 8'b10000111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????? :
        _3611_ = 8'b11001001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????? :
        _3611_ = 8'b00010101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????? :
        _3611_ = 8'b00111100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????? :
        _3611_ = 8'b00101101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????? :
        _3611_ = 8'b00110011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????? :
        _3611_ = 8'b00000111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????? :
        _3611_ = 8'b10101001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????? :
        _3611_ = 8'b11010010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????? :
        _3611_ = 8'b00100010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????? :
        _3611_ = 8'b00101011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????? :
        _3611_ = 8'b11101011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????? :
        _3611_ = 8'b11011001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????? :
        _3611_ = 8'b00100111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????? :
        _3611_ = 8'b00111010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????? :
        _3611_ = 8'b10011001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????? :
        _3611_ = 8'b00010111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????? :
        _3611_ = 8'b01101001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????? :
        _3611_ = 8'b10101110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????? :
        _3611_ = 8'b01101010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????? :
        _3611_ = 8'b11000010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????? :
        _3611_ = 8'b00011100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????? :
        _3611_ = 8'b11110111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????? :
        _3611_ = 8'b00000110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????? :
        _3611_ = 8'b10010000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????? :
        _3611_ = 8'b11001100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????? :
        _3611_ = 8'b01110001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????? :
        _3611_ = 8'b01111100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????? :
        _3611_ = 8'b11100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????? :
        _3611_ = 8'b00001111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????? :
        _3611_ = 8'b00001101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????? :
        _3611_ = 8'b01100001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????? :
        _3611_ = 8'b10010110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????? :
        _3611_ = 8'b00111110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????? :
        _3611_ = 8'b11101000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????? :
        _3611_ = 8'b10100001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????? :
        _3611_ = 8'b11001011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????? :
        _3611_ = 8'b10010111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????? :
        _3611_ = 8'b01110011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????? :
        _3611_ = 8'b01010111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????? :
        _3611_ = 8'b00111000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????? :
        _3611_ = 8'b01011100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????? :
        _3611_ = 8'b01001010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????? :
        _3611_ = 8'b11110000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????? :
        _3611_ = 8'b01101111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????? :
        _3611_ = 8'b00010000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b01000111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b11110100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b11001010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b11001111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b11110011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b10101100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b11011000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b01001001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b10011100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b10110001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b00000001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b11011010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b01101110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b10001011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b11010101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b11110010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b11010011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b00110001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b00111001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b11000100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b01000011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b10111101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b10011111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b10111000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b01001000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b00001100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b10010010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b00010100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b01110100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b01100100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b11011011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b10101101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b00010110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b10111100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b10100111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b00101000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b01101011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b11000111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b10001100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b00001011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b00111011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b01010100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b01000100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b10100011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b10011110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b00011001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b11000000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b11100110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b00110010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b10111010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b11001000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b01111010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b11111100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b01010101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b10010011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b00101110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b10001000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b00110101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b10111110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b11000011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b00100110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b00011000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b10000001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b10111111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b11111101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b11100101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b00100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b01000010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b10101111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b01110111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b01100011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b11110001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b01110000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b00100001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b00111111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b00000101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b10000000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b01011101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b10100010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b01001011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b00100101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b01111000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b10100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b11111110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b00000100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b11101001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b10001010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b00010001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b01100110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b10011010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b10000110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b11101101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b01001111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b11000101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b10111011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b10000101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b10110000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b10011000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b10010100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b01110010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b01100111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b10001101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b11010100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b10110110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b01111001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b11100011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b01000000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b11000001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b00000000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b10111001 ;
      256'b????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b10100110 ;
      256'b???????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b00010011 ;
      256'b??????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b01011110 ;
      256'b?????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b11011101 ;
      256'b????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b01010010 ;
      256'b???????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b01111101 ;
      256'b??????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b10110111 ;
      256'b?????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b01110110 ;
      256'b????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b10100100 ;
      256'b???????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b01011011 ;
      256'b??????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b10110100 ;
      256'b?????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b11011100 ;
      256'b????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b00110110 ;
      256'b???????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b00110100 ;
      256'b??????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b01011000 ;
      256'b?????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b00011101 ;
      256'b????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b00010010 ;
      256'b???????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b11101010 ;
      256'b??????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b01111111 ;
      256'b?????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b01001110 ;
      256'b????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b11001101 ;
      256'b???????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b11011111 ;
      256'b??????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b00011011 ;
      256'b?????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b00100100 ;
      256'b????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b00001110 ;
      256'b???????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b00101111 ;
      256'b??????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b00001010 ;
      256'b?????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b00110111 ;
      256'b????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b00110000 ;
      256'b???????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b10011101 ;
      256'b??????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b01000110 ;
      256'b?????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b10010101 ;
      256'b????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b00001000 ;
      256'b???????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b00101010 ;
      256'b??????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b01100010 ;
      256'b?????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b10101011 ;
      256'b????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b11100010 ;
      256'b???????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b11111001 ;
      256'b??????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b11010001 ;
      256'b?????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b01010001 ;
      256'b????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b01101000 ;
      256'b???????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b10000011 ;
      256'b??????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b11110101 ;
      256'b?????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b01111110 ;
      256'b????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b01101100 ;
      256'b???????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b01001100 ;
      256'b??????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b00111101 ;
      256'b?????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b11100001 ;
      256'b????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b01110101 ;
      256'b???????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b10011011 ;
      256'b??????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b11100100 ;
      256'b?????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b01010011 ;
      256'b????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b00100011 ;
      256'b???????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b01000101 ;
      256'b??????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b01011111 ;
      256'b?????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b10110011 ;
      256'b????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b01000001 ;
      256'b???????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b11111011 ;
      256'b??????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b10001110 ;
      256'b?????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b10110010 ;
      256'b????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b11101111 ;
      256'b???????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b11111010 ;
      256'b??????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b10001001 ;
      256'b?????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b00011111 ;
      256'b????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b10001111 ;
      256'b???????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b11101100 ;
      256'b??????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b01001101 ;
      256'b?????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b10110101 ;
      256'b????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b11100111 ;
      256'b???????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b01010110 ;
      256'b??????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b11001110 ;
      256'b?????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b00000010 ;
      256'b????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b01100000 ;
      256'b???????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b10010001 ;
      256'b??????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b11011110 ;
      256'b?????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b11010110 ;
      256'b????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b11111111 ;
      256'b???1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b11110110 ;
      256'b??1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b11101110 ;
      256'b?1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b11111000 ;
      256'b1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b11000110 ;
      default:
        _3611_ = \t3.t1.s4.out ;
    endcase
  end
  assign p32[23:16] = \t3.t2.s0.out ^ \t3.t2.s4.out ;
  always @(posedge clk)
      \t3.t2.s0.out <= _3612_;
  wire [255:0] fangyuan29;
  assign fangyuan29 = { _3868_, _3867_, _3866_, _3865_, _3864_, _3863_, _3862_, _3861_, _3860_, _3859_, _3858_, _3857_, _3856_, _3855_, _3854_, _3853_, _3852_, _3851_, _3850_, _3849_, _3848_, _3847_, _3846_, _3845_, _3844_, _3843_, _3842_, _3841_, _3840_, _3839_, _3838_, _3837_, _3836_, _3835_, _3834_, _3833_, _3832_, _3831_, _3830_, _3829_, _3828_, _3827_, _3826_, _3825_, _3824_, _3823_, _3822_, _3821_, _3820_, _3819_, _3818_, _3817_, _3816_, _3815_, _3814_, _3813_, _3812_, _3811_, _3810_, _3809_, _3808_, _3807_, _3806_, _3805_, _3804_, _3803_, _3802_, _3801_, _3800_, _3799_, _3798_, _3797_, _3796_, _3795_, _3794_, _3793_, _3792_, _3791_, _3790_, _3789_, _3788_, _3787_, _3786_, _3785_, _3784_, _3783_, _3782_, _3781_, _3780_, _3779_, _3778_, _3777_, _3776_, _3775_, _3774_, _3773_, _3772_, _3771_, _3770_, _3769_, _3768_, _3767_, _3766_, _3765_, _3764_, _3763_, _3762_, _3761_, _3760_, _3759_, _3758_, _3757_, _3756_, _3755_, _3754_, _3753_, _3752_, _3751_, _3750_, _3749_, _3748_, _3747_, _3746_, _3745_, _3744_, _3743_, _3742_, _3741_, _3740_, _3739_, _3738_, _3737_, _3736_, _3735_, _3734_, _3733_, _3732_, _3731_, _3730_, _3729_, _3728_, _3727_, _3726_, _3725_, _3724_, _3723_, _3722_, _3721_, _3720_, _3719_, _3718_, _3717_, _3716_, _3715_, _3714_, _3713_, _3712_, _3711_, _3710_, _3709_, _3708_, _3707_, _3706_, _3705_, _3704_, _3703_, _3702_, _3701_, _3700_, _3699_, _3698_, _3697_, _3696_, _3695_, _3694_, _3693_, _3692_, _3691_, _3690_, _3689_, _3688_, _3687_, _3686_, _3685_, _3684_, _3683_, _3682_, _3681_, _3680_, _3679_, _3678_, _3677_, _3676_, _3675_, _3674_, _3673_, _3672_, _3671_, _3670_, _3669_, _3668_, _3667_, _3666_, _3665_, _3664_, _3663_, _3662_, _3661_, _3660_, _3659_, _3658_, _3657_, _3656_, _3655_, _3654_, _3653_, _3652_, _3651_, _3650_, _3649_, _3648_, _3647_, _3646_, _3645_, _3644_, _3643_, _3642_, _3641_, _3640_, _3639_, _3638_, _3637_, _3636_, _3635_, _3634_, _3633_, _3632_, _3631_, _3630_, _3629_, _3628_, _3627_, _3626_, _3625_, _3624_, _3623_, _3622_, _3621_, _3620_, _3619_, _3618_, _3617_, _3616_, _3615_, _3614_, _3613_ };

  always @(\t3.t2.s0.out or fangyuan29) begin
    casez (fangyuan29)
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1 :
        _3612_ = 8'b00010110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1? :
        _3612_ = 8'b10111011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?? :
        _3612_ = 8'b01010100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??? :
        _3612_ = 8'b10110000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???? :
        _3612_ = 8'b00001111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????? :
        _3612_ = 8'b00101101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????? :
        _3612_ = 8'b10011001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????? :
        _3612_ = 8'b01000001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????? :
        _3612_ = 8'b01101000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????? :
        _3612_ = 8'b01000010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????? :
        _3612_ = 8'b11100110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????? :
        _3612_ = 8'b10111111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????? :
        _3612_ = 8'b00001101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????? :
        _3612_ = 8'b10001001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????? :
        _3612_ = 8'b10100001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????? :
        _3612_ = 8'b10001100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????? :
        _3612_ = 8'b11011111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????? :
        _3612_ = 8'b00101000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????? :
        _3612_ = 8'b01010101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????? :
        _3612_ = 8'b11001110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????? :
        _3612_ = 8'b11101001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????? :
        _3612_ = 8'b10000111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????? :
        _3612_ = 8'b00011110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????? :
        _3612_ = 8'b10011011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????? :
        _3612_ = 8'b10010100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????? :
        _3612_ = 8'b10001110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????? :
        _3612_ = 8'b11011001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????? :
        _3612_ = 8'b01101001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????? :
        _3612_ = 8'b00010001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????? :
        _3612_ = 8'b10011000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????? :
        _3612_ = 8'b11111000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????? :
        _3612_ = 8'b11100001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????? :
        _3612_ = 8'b10011110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????? :
        _3612_ = 8'b00011101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????? :
        _3612_ = 8'b11000001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????? :
        _3612_ = 8'b10000110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????? :
        _3612_ = 8'b10111001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????? :
        _3612_ = 8'b01010111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????? :
        _3612_ = 8'b00110101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????? :
        _3612_ = 8'b01100001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????? :
        _3612_ = 8'b00001110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????? :
        _3612_ = 8'b11110110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????? :
        _3612_ = 8'b00000011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????? :
        _3612_ = 8'b01001000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????? :
        _3612_ = 8'b01100110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????? :
        _3612_ = 8'b10110101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????? :
        _3612_ = 8'b00111110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????? :
        _3612_ = 8'b01110000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????? :
        _3612_ = 8'b10001010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????? :
        _3612_ = 8'b10001011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????? :
        _3612_ = 8'b10111101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????? :
        _3612_ = 8'b01001011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????? :
        _3612_ = 8'b00011111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????? :
        _3612_ = 8'b01110100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????? :
        _3612_ = 8'b11011101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????? :
        _3612_ = 8'b11101000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????? :
        _3612_ = 8'b11000110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????? :
        _3612_ = 8'b10110100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????? :
        _3612_ = 8'b10100110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????? :
        _3612_ = 8'b00011100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????? :
        _3612_ = 8'b00101110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????? :
        _3612_ = 8'b00100101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????? :
        _3612_ = 8'b01111000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????? :
        _3612_ = 8'b10111010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????? :
        _3612_ = 8'b00001000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b10101110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b01111010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b01100101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b11101010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b11110100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b01010110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b01101100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b10101001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b01001110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b11010101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b10001101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b01101101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b00110111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b11001000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b11100111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b01111001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b11100100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b10010101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b10010001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b01100010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b10101100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b11010011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b11000010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b01011100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b00100100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b00000110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b01001001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b00001010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b00111010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b00110010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b11100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b11011011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b00001011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b01011110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b11011110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b00010100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b10111000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b11101110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b01000110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b10001000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b10010000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b00101010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b00100010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b11011100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b01001111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b10000001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b01100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b01110011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b00011001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b01011101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b01100100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b00111101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b01111110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b10100111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b11000100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b00010111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b01000100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b10010111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b01011111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b11101100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b00010011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b00001100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b11001101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b11010010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b11110011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b11111111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b00010000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b00100001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b11011010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b10110110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b10111100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b11110101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b00111000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b10011101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b10010010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b10001111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b01000000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b10100011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b01010001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b10101000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b10011111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b00111100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b01010000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b01111111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b00000010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b11111001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b01000101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b10000101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b00110011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b01001101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b01000011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b11111011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b10101010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b11101111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b11010000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b11001111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b01011000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b01001100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b01001010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b00111001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b10111110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b11001011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b01101010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b01011011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b10110001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b11111100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b00100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b11101101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b00000000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b11010001 ;
      256'b????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b01010011 ;
      256'b???????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b10000100 ;
      256'b??????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b00101111 ;
      256'b?????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b11100011 ;
      256'b????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b00101001 ;
      256'b???????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b10110011 ;
      256'b??????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b11010110 ;
      256'b?????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b00111011 ;
      256'b????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b01010010 ;
      256'b???????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b10100000 ;
      256'b??????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b01011010 ;
      256'b?????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b01101110 ;
      256'b????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b00011011 ;
      256'b???????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b00011010 ;
      256'b??????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b00101100 ;
      256'b?????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b10000011 ;
      256'b????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b00001001 ;
      256'b???????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b01110101 ;
      256'b??????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b10110010 ;
      256'b?????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b00100111 ;
      256'b????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b11101011 ;
      256'b???????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b11100010 ;
      256'b??????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b10000000 ;
      256'b?????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b00010010 ;
      256'b????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b00000111 ;
      256'b???????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b10011010 ;
      256'b??????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b00000101 ;
      256'b?????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b10010110 ;
      256'b????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b00011000 ;
      256'b???????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b11000011 ;
      256'b??????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b00100011 ;
      256'b?????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b11000111 ;
      256'b????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b00000100 ;
      256'b???????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b00010101 ;
      256'b??????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b00110001 ;
      256'b?????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b11011000 ;
      256'b????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b01110001 ;
      256'b???????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b11110001 ;
      256'b??????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b11100101 ;
      256'b?????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b10100101 ;
      256'b????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b00110100 ;
      256'b???????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b11001100 ;
      256'b??????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b11110111 ;
      256'b?????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b00111111 ;
      256'b????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b00110110 ;
      256'b???????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b00100110 ;
      256'b??????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b10010011 ;
      256'b?????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b11111101 ;
      256'b????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b10110111 ;
      256'b???????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b11000000 ;
      256'b??????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b01110010 ;
      256'b?????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b10100100 ;
      256'b????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b10011100 ;
      256'b???????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b10101111 ;
      256'b??????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b10100010 ;
      256'b?????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b11010100 ;
      256'b????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b10101101 ;
      256'b???????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b11110000 ;
      256'b??????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b01000111 ;
      256'b?????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b01011001 ;
      256'b????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b11111010 ;
      256'b???????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b01111101 ;
      256'b??????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b11001001 ;
      256'b?????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b10000010 ;
      256'b????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b11001010 ;
      256'b???????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b01110110 ;
      256'b??????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b10101011 ;
      256'b?????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b11010111 ;
      256'b????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b11111110 ;
      256'b???????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b00101011 ;
      256'b??????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b01100111 ;
      256'b?????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b00000001 ;
      256'b????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b00110000 ;
      256'b???????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b11000101 ;
      256'b??????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b01101111 ;
      256'b?????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b01101011 ;
      256'b????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b11110010 ;
      256'b???1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b01111011 ;
      256'b??1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b01110111 ;
      256'b?1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b01111100 ;
      256'b1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b01100011 ;
      default:
        _3612_ = \t3.t2.s0.out ;
    endcase
  end
  assign _3613_ = state_in[15:8] == 8'b11111111;
  assign _3614_ = state_in[15:8] == 8'b11111110;
  assign _3615_ = state_in[15:8] == 8'b11111101;
  assign _3616_ = state_in[15:8] == 8'b11111100;
  assign _3617_ = state_in[15:8] == 8'b11111011;
  assign _3618_ = state_in[15:8] == 8'b11111010;
  assign _3619_ = state_in[15:8] == 8'b11111001;
  assign _3620_ = state_in[15:8] == 8'b11111000;
  assign _3621_ = state_in[15:8] == 8'b11110111;
  assign _3622_ = state_in[15:8] == 8'b11110110;
  assign _3623_ = state_in[15:8] == 8'b11110101;
  assign _3624_ = state_in[15:8] == 8'b11110100;
  assign _3625_ = state_in[15:8] == 8'b11110011;
  assign _3626_ = state_in[15:8] == 8'b11110010;
  assign _3627_ = state_in[15:8] == 8'b11110001;
  assign _3628_ = state_in[15:8] == 8'b11110000;
  assign _3629_ = state_in[15:8] == 8'b11101111;
  assign _3630_ = state_in[15:8] == 8'b11101110;
  assign _3631_ = state_in[15:8] == 8'b11101101;
  assign _3632_ = state_in[15:8] == 8'b11101100;
  assign _3633_ = state_in[15:8] == 8'b11101011;
  assign _3634_ = state_in[15:8] == 8'b11101010;
  assign _3635_ = state_in[15:8] == 8'b11101001;
  assign _3636_ = state_in[15:8] == 8'b11101000;
  assign _3637_ = state_in[15:8] == 8'b11100111;
  assign _3638_ = state_in[15:8] == 8'b11100110;
  assign _3639_ = state_in[15:8] == 8'b11100101;
  assign _3640_ = state_in[15:8] == 8'b11100100;
  assign _3641_ = state_in[15:8] == 8'b11100011;
  assign _3642_ = state_in[15:8] == 8'b11100010;
  assign _3643_ = state_in[15:8] == 8'b11100001;
  assign _3644_ = state_in[15:8] == 8'b11100000;
  assign _3645_ = state_in[15:8] == 8'b11011111;
  assign _3646_ = state_in[15:8] == 8'b11011110;
  assign _3647_ = state_in[15:8] == 8'b11011101;
  assign _3648_ = state_in[15:8] == 8'b11011100;
  assign _3649_ = state_in[15:8] == 8'b11011011;
  assign _3650_ = state_in[15:8] == 8'b11011010;
  assign _3651_ = state_in[15:8] == 8'b11011001;
  assign _3652_ = state_in[15:8] == 8'b11011000;
  assign _3653_ = state_in[15:8] == 8'b11010111;
  assign _3654_ = state_in[15:8] == 8'b11010110;
  assign _3655_ = state_in[15:8] == 8'b11010101;
  assign _3656_ = state_in[15:8] == 8'b11010100;
  assign _3657_ = state_in[15:8] == 8'b11010011;
  assign _3658_ = state_in[15:8] == 8'b11010010;
  assign _3659_ = state_in[15:8] == 8'b11010001;
  assign _3660_ = state_in[15:8] == 8'b11010000;
  assign _3661_ = state_in[15:8] == 8'b11001111;
  assign _3662_ = state_in[15:8] == 8'b11001110;
  assign _3663_ = state_in[15:8] == 8'b11001101;
  assign _3664_ = state_in[15:8] == 8'b11001100;
  assign _3665_ = state_in[15:8] == 8'b11001011;
  assign _3666_ = state_in[15:8] == 8'b11001010;
  assign _3667_ = state_in[15:8] == 8'b11001001;
  assign _3668_ = state_in[15:8] == 8'b11001000;
  assign _3669_ = state_in[15:8] == 8'b11000111;
  assign _3670_ = state_in[15:8] == 8'b11000110;
  assign _3671_ = state_in[15:8] == 8'b11000101;
  assign _3672_ = state_in[15:8] == 8'b11000100;
  assign _3673_ = state_in[15:8] == 8'b11000011;
  assign _3674_ = state_in[15:8] == 8'b11000010;
  assign _3675_ = state_in[15:8] == 8'b11000001;
  assign _3676_ = state_in[15:8] == 8'b11000000;
  assign _3677_ = state_in[15:8] == 8'b10111111;
  assign _3678_ = state_in[15:8] == 8'b10111110;
  assign _3679_ = state_in[15:8] == 8'b10111101;
  assign _3680_ = state_in[15:8] == 8'b10111100;
  assign _3681_ = state_in[15:8] == 8'b10111011;
  assign _3682_ = state_in[15:8] == 8'b10111010;
  assign _3683_ = state_in[15:8] == 8'b10111001;
  assign _3684_ = state_in[15:8] == 8'b10111000;
  assign _3685_ = state_in[15:8] == 8'b10110111;
  assign _3686_ = state_in[15:8] == 8'b10110110;
  assign _3687_ = state_in[15:8] == 8'b10110101;
  assign _3688_ = state_in[15:8] == 8'b10110100;
  assign _3689_ = state_in[15:8] == 8'b10110011;
  assign _3690_ = state_in[15:8] == 8'b10110010;
  assign _3691_ = state_in[15:8] == 8'b10110001;
  assign _3692_ = state_in[15:8] == 8'b10110000;
  assign _3693_ = state_in[15:8] == 8'b10101111;
  assign _3694_ = state_in[15:8] == 8'b10101110;
  assign _3695_ = state_in[15:8] == 8'b10101101;
  assign _3696_ = state_in[15:8] == 8'b10101100;
  assign _3697_ = state_in[15:8] == 8'b10101011;
  assign _3698_ = state_in[15:8] == 8'b10101010;
  assign _3699_ = state_in[15:8] == 8'b10101001;
  assign _3700_ = state_in[15:8] == 8'b10101000;
  assign _3701_ = state_in[15:8] == 8'b10100111;
  assign _3702_ = state_in[15:8] == 8'b10100110;
  assign _3703_ = state_in[15:8] == 8'b10100101;
  assign _3704_ = state_in[15:8] == 8'b10100100;
  assign _3705_ = state_in[15:8] == 8'b10100011;
  assign _3706_ = state_in[15:8] == 8'b10100010;
  assign _3707_ = state_in[15:8] == 8'b10100001;
  assign _3708_ = state_in[15:8] == 8'b10100000;
  assign _3709_ = state_in[15:8] == 8'b10011111;
  assign _3710_ = state_in[15:8] == 8'b10011110;
  assign _3711_ = state_in[15:8] == 8'b10011101;
  assign _3712_ = state_in[15:8] == 8'b10011100;
  assign _3713_ = state_in[15:8] == 8'b10011011;
  assign _3714_ = state_in[15:8] == 8'b10011010;
  assign _3715_ = state_in[15:8] == 8'b10011001;
  assign _3716_ = state_in[15:8] == 8'b10011000;
  assign _3717_ = state_in[15:8] == 8'b10010111;
  assign _3718_ = state_in[15:8] == 8'b10010110;
  assign _3719_ = state_in[15:8] == 8'b10010101;
  assign _3720_ = state_in[15:8] == 8'b10010100;
  assign _3721_ = state_in[15:8] == 8'b10010011;
  assign _3722_ = state_in[15:8] == 8'b10010010;
  assign _3723_ = state_in[15:8] == 8'b10010001;
  assign _3724_ = state_in[15:8] == 8'b10010000;
  assign _3725_ = state_in[15:8] == 8'b10001111;
  assign _3726_ = state_in[15:8] == 8'b10001110;
  assign _3727_ = state_in[15:8] == 8'b10001101;
  assign _3728_ = state_in[15:8] == 8'b10001100;
  assign _3729_ = state_in[15:8] == 8'b10001011;
  assign _3730_ = state_in[15:8] == 8'b10001010;
  assign _3731_ = state_in[15:8] == 8'b10001001;
  assign _3732_ = state_in[15:8] == 8'b10001000;
  assign _3733_ = state_in[15:8] == 8'b10000111;
  assign _3734_ = state_in[15:8] == 8'b10000110;
  assign _3735_ = state_in[15:8] == 8'b10000101;
  assign _3736_ = state_in[15:8] == 8'b10000100;
  assign _3737_ = state_in[15:8] == 8'b10000011;
  assign _3738_ = state_in[15:8] == 8'b10000010;
  assign _3739_ = state_in[15:8] == 8'b10000001;
  assign _3740_ = state_in[15:8] == 8'b10000000;
  assign _3741_ = state_in[15:8] == 7'b1111111;
  assign _3742_ = state_in[15:8] == 7'b1111110;
  assign _3743_ = state_in[15:8] == 7'b1111101;
  assign _3744_ = state_in[15:8] == 7'b1111100;
  assign _3745_ = state_in[15:8] == 7'b1111011;
  assign _3746_ = state_in[15:8] == 7'b1111010;
  assign _3747_ = state_in[15:8] == 7'b1111001;
  assign _3748_ = state_in[15:8] == 7'b1111000;
  assign _3749_ = state_in[15:8] == 7'b1110111;
  assign _3750_ = state_in[15:8] == 7'b1110110;
  assign _3751_ = state_in[15:8] == 7'b1110101;
  assign _3752_ = state_in[15:8] == 7'b1110100;
  assign _3753_ = state_in[15:8] == 7'b1110011;
  assign _3754_ = state_in[15:8] == 7'b1110010;
  assign _3755_ = state_in[15:8] == 7'b1110001;
  assign _3756_ = state_in[15:8] == 7'b1110000;
  assign _3757_ = state_in[15:8] == 7'b1101111;
  assign _3758_ = state_in[15:8] == 7'b1101110;
  assign _3759_ = state_in[15:8] == 7'b1101101;
  assign _3760_ = state_in[15:8] == 7'b1101100;
  assign _3761_ = state_in[15:8] == 7'b1101011;
  assign _3762_ = state_in[15:8] == 7'b1101010;
  assign _3763_ = state_in[15:8] == 7'b1101001;
  assign _3764_ = state_in[15:8] == 7'b1101000;
  assign _3765_ = state_in[15:8] == 7'b1100111;
  assign _3766_ = state_in[15:8] == 7'b1100110;
  assign _3767_ = state_in[15:8] == 7'b1100101;
  assign _3768_ = state_in[15:8] == 7'b1100100;
  assign _3769_ = state_in[15:8] == 7'b1100011;
  assign _3770_ = state_in[15:8] == 7'b1100010;
  assign _3771_ = state_in[15:8] == 7'b1100001;
  assign _3772_ = state_in[15:8] == 7'b1100000;
  assign _3773_ = state_in[15:8] == 7'b1011111;
  assign _3774_ = state_in[15:8] == 7'b1011110;
  assign _3775_ = state_in[15:8] == 7'b1011101;
  assign _3776_ = state_in[15:8] == 7'b1011100;
  assign _3777_ = state_in[15:8] == 7'b1011011;
  assign _3778_ = state_in[15:8] == 7'b1011010;
  assign _3779_ = state_in[15:8] == 7'b1011001;
  assign _3780_ = state_in[15:8] == 7'b1011000;
  assign _3781_ = state_in[15:8] == 7'b1010111;
  assign _3782_ = state_in[15:8] == 7'b1010110;
  assign _3783_ = state_in[15:8] == 7'b1010101;
  assign _3784_ = state_in[15:8] == 7'b1010100;
  assign _3785_ = state_in[15:8] == 7'b1010011;
  assign _3786_ = state_in[15:8] == 7'b1010010;
  assign _3787_ = state_in[15:8] == 7'b1010001;
  assign _3788_ = state_in[15:8] == 7'b1010000;
  assign _3789_ = state_in[15:8] == 7'b1001111;
  assign _3790_ = state_in[15:8] == 7'b1001110;
  assign _3791_ = state_in[15:8] == 7'b1001101;
  assign _3792_ = state_in[15:8] == 7'b1001100;
  assign _3793_ = state_in[15:8] == 7'b1001011;
  assign _3794_ = state_in[15:8] == 7'b1001010;
  assign _3795_ = state_in[15:8] == 7'b1001001;
  assign _3796_ = state_in[15:8] == 7'b1001000;
  assign _3797_ = state_in[15:8] == 7'b1000111;
  assign _3798_ = state_in[15:8] == 7'b1000110;
  assign _3799_ = state_in[15:8] == 7'b1000101;
  assign _3800_ = state_in[15:8] == 7'b1000100;
  assign _3801_ = state_in[15:8] == 7'b1000011;
  assign _3802_ = state_in[15:8] == 7'b1000010;
  assign _3803_ = state_in[15:8] == 7'b1000001;
  assign _3804_ = state_in[15:8] == 7'b1000000;
  assign _3805_ = state_in[15:8] == 6'b111111;
  assign _3806_ = state_in[15:8] == 6'b111110;
  assign _3807_ = state_in[15:8] == 6'b111101;
  assign _3808_ = state_in[15:8] == 6'b111100;
  assign _3809_ = state_in[15:8] == 6'b111011;
  assign _3810_ = state_in[15:8] == 6'b111010;
  assign _3811_ = state_in[15:8] == 6'b111001;
  assign _3812_ = state_in[15:8] == 6'b111000;
  assign _3813_ = state_in[15:8] == 6'b110111;
  assign _3814_ = state_in[15:8] == 6'b110110;
  assign _3815_ = state_in[15:8] == 6'b110101;
  assign _3816_ = state_in[15:8] == 6'b110100;
  assign _3817_ = state_in[15:8] == 6'b110011;
  assign _3818_ = state_in[15:8] == 6'b110010;
  assign _3819_ = state_in[15:8] == 6'b110001;
  assign _3820_ = state_in[15:8] == 6'b110000;
  assign _3821_ = state_in[15:8] == 6'b101111;
  assign _3822_ = state_in[15:8] == 6'b101110;
  assign _3823_ = state_in[15:8] == 6'b101101;
  assign _3824_ = state_in[15:8] == 6'b101100;
  assign _3825_ = state_in[15:8] == 6'b101011;
  assign _3826_ = state_in[15:8] == 6'b101010;
  assign _3827_ = state_in[15:8] == 6'b101001;
  assign _3828_ = state_in[15:8] == 6'b101000;
  assign _3829_ = state_in[15:8] == 6'b100111;
  assign _3830_ = state_in[15:8] == 6'b100110;
  assign _3831_ = state_in[15:8] == 6'b100101;
  assign _3832_ = state_in[15:8] == 6'b100100;
  assign _3833_ = state_in[15:8] == 6'b100011;
  assign _3834_ = state_in[15:8] == 6'b100010;
  assign _3835_ = state_in[15:8] == 6'b100001;
  assign _3836_ = state_in[15:8] == 6'b100000;
  assign _3837_ = state_in[15:8] == 5'b11111;
  assign _3838_ = state_in[15:8] == 5'b11110;
  assign _3839_ = state_in[15:8] == 5'b11101;
  assign _3840_ = state_in[15:8] == 5'b11100;
  assign _3841_ = state_in[15:8] == 5'b11011;
  assign _3842_ = state_in[15:8] == 5'b11010;
  assign _3843_ = state_in[15:8] == 5'b11001;
  assign _3844_ = state_in[15:8] == 5'b11000;
  assign _3845_ = state_in[15:8] == 5'b10111;
  assign _3846_ = state_in[15:8] == 5'b10110;
  assign _3847_ = state_in[15:8] == 5'b10101;
  assign _3848_ = state_in[15:8] == 5'b10100;
  assign _3849_ = state_in[15:8] == 5'b10011;
  assign _3850_ = state_in[15:8] == 5'b10010;
  assign _3851_ = state_in[15:8] == 5'b10001;
  assign _3852_ = state_in[15:8] == 5'b10000;
  assign _3853_ = state_in[15:8] == 4'b1111;
  assign _3854_ = state_in[15:8] == 4'b1110;
  assign _3855_ = state_in[15:8] == 4'b1101;
  assign _3856_ = state_in[15:8] == 4'b1100;
  assign _3857_ = state_in[15:8] == 4'b1011;
  assign _3858_ = state_in[15:8] == 4'b1010;
  assign _3859_ = state_in[15:8] == 4'b1001;
  assign _3860_ = state_in[15:8] == 4'b1000;
  assign _3861_ = state_in[15:8] == 3'b111;
  assign _3862_ = state_in[15:8] == 3'b110;
  assign _3863_ = state_in[15:8] == 3'b101;
  assign _3864_ = state_in[15:8] == 3'b100;
  assign _3865_ = state_in[15:8] == 2'b11;
  assign _3866_ = state_in[15:8] == 2'b10;
  assign _3867_ = state_in[15:8] == 1'b1;
  assign _3868_ = ! state_in[15:8];
  always @(posedge clk)
      \t3.t2.s4.out <= _3869_;
  wire [255:0] fangyuan30;
  assign fangyuan30 = { _3868_, _3867_, _3866_, _3865_, _3864_, _3863_, _3862_, _3861_, _3860_, _3859_, _3858_, _3857_, _3856_, _3855_, _3854_, _3853_, _3852_, _3851_, _3850_, _3849_, _3848_, _3847_, _3846_, _3845_, _3844_, _3843_, _3842_, _3841_, _3840_, _3839_, _3838_, _3837_, _3836_, _3835_, _3834_, _3833_, _3832_, _3831_, _3830_, _3829_, _3828_, _3827_, _3826_, _3825_, _3824_, _3823_, _3822_, _3821_, _3820_, _3819_, _3818_, _3817_, _3816_, _3815_, _3814_, _3813_, _3812_, _3811_, _3810_, _3809_, _3808_, _3807_, _3806_, _3805_, _3804_, _3803_, _3802_, _3801_, _3800_, _3799_, _3798_, _3797_, _3796_, _3795_, _3794_, _3793_, _3792_, _3791_, _3790_, _3789_, _3788_, _3787_, _3786_, _3785_, _3784_, _3783_, _3782_, _3781_, _3780_, _3779_, _3778_, _3777_, _3776_, _3775_, _3774_, _3773_, _3772_, _3771_, _3770_, _3769_, _3768_, _3767_, _3766_, _3765_, _3764_, _3763_, _3762_, _3761_, _3760_, _3759_, _3758_, _3757_, _3756_, _3755_, _3754_, _3753_, _3752_, _3751_, _3750_, _3749_, _3748_, _3747_, _3746_, _3745_, _3744_, _3743_, _3742_, _3741_, _3740_, _3739_, _3738_, _3737_, _3736_, _3735_, _3734_, _3733_, _3732_, _3731_, _3730_, _3729_, _3728_, _3727_, _3726_, _3725_, _3724_, _3723_, _3722_, _3721_, _3720_, _3719_, _3718_, _3717_, _3716_, _3715_, _3714_, _3713_, _3712_, _3711_, _3710_, _3709_, _3708_, _3707_, _3706_, _3705_, _3704_, _3703_, _3702_, _3701_, _3700_, _3699_, _3698_, _3697_, _3696_, _3695_, _3694_, _3693_, _3692_, _3691_, _3690_, _3689_, _3688_, _3687_, _3686_, _3685_, _3684_, _3683_, _3682_, _3681_, _3680_, _3679_, _3678_, _3677_, _3676_, _3675_, _3674_, _3673_, _3672_, _3671_, _3670_, _3669_, _3668_, _3667_, _3666_, _3665_, _3664_, _3663_, _3662_, _3661_, _3660_, _3659_, _3658_, _3657_, _3656_, _3655_, _3654_, _3653_, _3652_, _3651_, _3650_, _3649_, _3648_, _3647_, _3646_, _3645_, _3644_, _3643_, _3642_, _3641_, _3640_, _3639_, _3638_, _3637_, _3636_, _3635_, _3634_, _3633_, _3632_, _3631_, _3630_, _3629_, _3628_, _3627_, _3626_, _3625_, _3624_, _3623_, _3622_, _3621_, _3620_, _3619_, _3618_, _3617_, _3616_, _3615_, _3614_, _3613_ };

  always @(\t3.t2.s4.out or fangyuan30) begin
    casez (fangyuan30)
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1 :
        _3869_ = 8'b00101100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1? :
        _3869_ = 8'b01101101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?? :
        _3869_ = 8'b10101000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??? :
        _3869_ = 8'b01111011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???? :
        _3869_ = 8'b00011110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????? :
        _3869_ = 8'b01011010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????? :
        _3869_ = 8'b00101001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????? :
        _3869_ = 8'b10000010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????? :
        _3869_ = 8'b11010000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????? :
        _3869_ = 8'b10000100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????? :
        _3869_ = 8'b11010111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????? :
        _3869_ = 8'b01100101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????? :
        _3869_ = 8'b00011010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????? :
        _3869_ = 8'b00001001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????? :
        _3869_ = 8'b01011001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????? :
        _3869_ = 8'b00000011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????? :
        _3869_ = 8'b10100101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????? :
        _3869_ = 8'b01010000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????? :
        _3869_ = 8'b10101010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????? :
        _3869_ = 8'b10000111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????? :
        _3869_ = 8'b11001001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????? :
        _3869_ = 8'b00010101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????? :
        _3869_ = 8'b00111100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????? :
        _3869_ = 8'b00101101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????? :
        _3869_ = 8'b00110011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????? :
        _3869_ = 8'b00000111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????? :
        _3869_ = 8'b10101001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????? :
        _3869_ = 8'b11010010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????? :
        _3869_ = 8'b00100010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????? :
        _3869_ = 8'b00101011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????? :
        _3869_ = 8'b11101011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????? :
        _3869_ = 8'b11011001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????? :
        _3869_ = 8'b00100111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????? :
        _3869_ = 8'b00111010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????? :
        _3869_ = 8'b10011001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????? :
        _3869_ = 8'b00010111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????? :
        _3869_ = 8'b01101001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????? :
        _3869_ = 8'b10101110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????? :
        _3869_ = 8'b01101010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????? :
        _3869_ = 8'b11000010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????? :
        _3869_ = 8'b00011100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????? :
        _3869_ = 8'b11110111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????? :
        _3869_ = 8'b00000110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????? :
        _3869_ = 8'b10010000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????? :
        _3869_ = 8'b11001100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????? :
        _3869_ = 8'b01110001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????? :
        _3869_ = 8'b01111100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????? :
        _3869_ = 8'b11100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????? :
        _3869_ = 8'b00001111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????? :
        _3869_ = 8'b00001101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????? :
        _3869_ = 8'b01100001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????? :
        _3869_ = 8'b10010110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????? :
        _3869_ = 8'b00111110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????? :
        _3869_ = 8'b11101000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????? :
        _3869_ = 8'b10100001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????? :
        _3869_ = 8'b11001011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????? :
        _3869_ = 8'b10010111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????? :
        _3869_ = 8'b01110011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????? :
        _3869_ = 8'b01010111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????? :
        _3869_ = 8'b00111000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????? :
        _3869_ = 8'b01011100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????? :
        _3869_ = 8'b01001010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????? :
        _3869_ = 8'b11110000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????? :
        _3869_ = 8'b01101111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????? :
        _3869_ = 8'b00010000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b01000111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b11110100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b11001010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b11001111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b11110011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b10101100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b11011000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b01001001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b10011100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b10110001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b00000001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b11011010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b01101110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b10001011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b11010101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b11110010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b11010011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b00110001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b00111001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b11000100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b01000011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b10111101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b10011111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b10111000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b01001000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b00001100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b10010010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b00010100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b01110100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b01100100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b11011011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b10101101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b00010110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b10111100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b10100111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b00101000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b01101011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b11000111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b10001100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b00001011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b00111011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b01010100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b01000100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b10100011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b10011110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b00011001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b11000000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b11100110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b00110010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b10111010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b11001000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b01111010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b11111100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b01010101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b10010011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b00101110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b10001000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b00110101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b10111110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b11000011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b00100110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b00011000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b10000001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b10111111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b11111101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b11100101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b00100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b01000010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b10101111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b01110111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b01100011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b11110001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b01110000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b00100001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b00111111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b00000101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b10000000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b01011101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b10100010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b01001011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b00100101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b01111000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b10100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b11111110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b00000100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b11101001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b10001010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b00010001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b01100110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b10011010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b10000110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b11101101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b01001111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b11000101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b10111011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b10000101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b10110000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b10011000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b10010100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b01110010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b01100111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b10001101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b11010100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b10110110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b01111001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b11100011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b01000000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b11000001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b00000000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b10111001 ;
      256'b????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b10100110 ;
      256'b???????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b00010011 ;
      256'b??????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b01011110 ;
      256'b?????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b11011101 ;
      256'b????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b01010010 ;
      256'b???????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b01111101 ;
      256'b??????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b10110111 ;
      256'b?????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b01110110 ;
      256'b????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b10100100 ;
      256'b???????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b01011011 ;
      256'b??????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b10110100 ;
      256'b?????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b11011100 ;
      256'b????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b00110110 ;
      256'b???????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b00110100 ;
      256'b??????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b01011000 ;
      256'b?????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b00011101 ;
      256'b????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b00010010 ;
      256'b???????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b11101010 ;
      256'b??????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b01111111 ;
      256'b?????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b01001110 ;
      256'b????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b11001101 ;
      256'b???????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b11011111 ;
      256'b??????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b00011011 ;
      256'b?????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b00100100 ;
      256'b????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b00001110 ;
      256'b???????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b00101111 ;
      256'b??????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b00001010 ;
      256'b?????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b00110111 ;
      256'b????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b00110000 ;
      256'b???????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b10011101 ;
      256'b??????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b01000110 ;
      256'b?????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b10010101 ;
      256'b????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b00001000 ;
      256'b???????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b00101010 ;
      256'b??????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b01100010 ;
      256'b?????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b10101011 ;
      256'b????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b11100010 ;
      256'b???????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b11111001 ;
      256'b??????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b11010001 ;
      256'b?????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b01010001 ;
      256'b????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b01101000 ;
      256'b???????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b10000011 ;
      256'b??????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b11110101 ;
      256'b?????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b01111110 ;
      256'b????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b01101100 ;
      256'b???????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b01001100 ;
      256'b??????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b00111101 ;
      256'b?????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b11100001 ;
      256'b????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b01110101 ;
      256'b???????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b10011011 ;
      256'b??????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b11100100 ;
      256'b?????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b01010011 ;
      256'b????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b00100011 ;
      256'b???????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b01000101 ;
      256'b??????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b01011111 ;
      256'b?????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b10110011 ;
      256'b????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b01000001 ;
      256'b???????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b11111011 ;
      256'b??????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b10001110 ;
      256'b?????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b10110010 ;
      256'b????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b11101111 ;
      256'b???????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b11111010 ;
      256'b??????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b10001001 ;
      256'b?????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b00011111 ;
      256'b????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b10001111 ;
      256'b???????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b11101100 ;
      256'b??????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b01001101 ;
      256'b?????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b10110101 ;
      256'b????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b11100111 ;
      256'b???????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b01010110 ;
      256'b??????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b11001110 ;
      256'b?????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b00000010 ;
      256'b????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b01100000 ;
      256'b???????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b10010001 ;
      256'b??????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b11011110 ;
      256'b?????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b11010110 ;
      256'b????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b11111111 ;
      256'b???1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b11110110 ;
      256'b??1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b11101110 ;
      256'b?1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b11111000 ;
      256'b1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b11000110 ;
      default:
        _3869_ = \t3.t2.s4.out ;
    endcase
  end
  assign p33[15:8] = \t3.t3.s0.out ^ \t3.t3.s4.out ;
  always @(posedge clk)
      \t3.t3.s0.out <= _3870_;
  wire [255:0] fangyuan31;
  assign fangyuan31 = { _4126_, _4125_, _4124_, _4123_, _4122_, _4121_, _4120_, _4119_, _4118_, _4117_, _4116_, _4115_, _4114_, _4113_, _4112_, _4111_, _4110_, _4109_, _4108_, _4107_, _4106_, _4105_, _4104_, _4103_, _4102_, _4101_, _4100_, _4099_, _4098_, _4097_, _4096_, _4095_, _4094_, _4093_, _4092_, _4091_, _4090_, _4089_, _4088_, _4087_, _4086_, _4085_, _4084_, _4083_, _4082_, _4081_, _4080_, _4079_, _4078_, _4077_, _4076_, _4075_, _4074_, _4073_, _4072_, _4071_, _4070_, _4069_, _4068_, _4067_, _4066_, _4065_, _4064_, _4063_, _4062_, _4061_, _4060_, _4059_, _4058_, _4057_, _4056_, _4055_, _4054_, _4053_, _4052_, _4051_, _4050_, _4049_, _4048_, _4047_, _4046_, _4045_, _4044_, _4043_, _4042_, _4041_, _4040_, _4039_, _4038_, _4037_, _4036_, _4035_, _4034_, _4033_, _4032_, _4031_, _4030_, _4029_, _4028_, _4027_, _4026_, _4025_, _4024_, _4023_, _4022_, _4021_, _4020_, _4019_, _4018_, _4017_, _4016_, _4015_, _4014_, _4013_, _4012_, _4011_, _4010_, _4009_, _4008_, _4007_, _4006_, _4005_, _4004_, _4003_, _4002_, _4001_, _4000_, _3999_, _3998_, _3997_, _3996_, _3995_, _3994_, _3993_, _3992_, _3991_, _3990_, _3989_, _3988_, _3987_, _3986_, _3985_, _3984_, _3983_, _3982_, _3981_, _3980_, _3979_, _3978_, _3977_, _3976_, _3975_, _3974_, _3973_, _3972_, _3971_, _3970_, _3969_, _3968_, _3967_, _3966_, _3965_, _3964_, _3963_, _3962_, _3961_, _3960_, _3959_, _3958_, _3957_, _3956_, _3955_, _3954_, _3953_, _3952_, _3951_, _3950_, _3949_, _3948_, _3947_, _3946_, _3945_, _3944_, _3943_, _3942_, _3941_, _3940_, _3939_, _3938_, _3937_, _3936_, _3935_, _3934_, _3933_, _3932_, _3931_, _3930_, _3929_, _3928_, _3927_, _3926_, _3925_, _3924_, _3923_, _3922_, _3921_, _3920_, _3919_, _3918_, _3917_, _3916_, _3915_, _3914_, _3913_, _3912_, _3911_, _3910_, _3909_, _3908_, _3907_, _3906_, _3905_, _3904_, _3903_, _3902_, _3901_, _3900_, _3899_, _3898_, _3897_, _3896_, _3895_, _3894_, _3893_, _3892_, _3891_, _3890_, _3889_, _3888_, _3887_, _3886_, _3885_, _3884_, _3883_, _3882_, _3881_, _3880_, _3879_, _3878_, _3877_, _3876_, _3875_, _3874_, _3873_, _3872_, _3871_ };

  always @(\t3.t3.s0.out or fangyuan31) begin
    casez (fangyuan31)
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1 :
        _3870_ = 8'b00010110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1? :
        _3870_ = 8'b10111011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?? :
        _3870_ = 8'b01010100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??? :
        _3870_ = 8'b10110000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???? :
        _3870_ = 8'b00001111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????? :
        _3870_ = 8'b00101101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????? :
        _3870_ = 8'b10011001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????? :
        _3870_ = 8'b01000001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????? :
        _3870_ = 8'b01101000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????? :
        _3870_ = 8'b01000010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????? :
        _3870_ = 8'b11100110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????? :
        _3870_ = 8'b10111111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????? :
        _3870_ = 8'b00001101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????? :
        _3870_ = 8'b10001001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????? :
        _3870_ = 8'b10100001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????? :
        _3870_ = 8'b10001100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????? :
        _3870_ = 8'b11011111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????? :
        _3870_ = 8'b00101000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????? :
        _3870_ = 8'b01010101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????? :
        _3870_ = 8'b11001110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????? :
        _3870_ = 8'b11101001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????? :
        _3870_ = 8'b10000111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????? :
        _3870_ = 8'b00011110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????? :
        _3870_ = 8'b10011011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????? :
        _3870_ = 8'b10010100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????? :
        _3870_ = 8'b10001110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????? :
        _3870_ = 8'b11011001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????? :
        _3870_ = 8'b01101001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????? :
        _3870_ = 8'b00010001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????? :
        _3870_ = 8'b10011000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????? :
        _3870_ = 8'b11111000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????? :
        _3870_ = 8'b11100001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????? :
        _3870_ = 8'b10011110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????? :
        _3870_ = 8'b00011101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????? :
        _3870_ = 8'b11000001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????? :
        _3870_ = 8'b10000110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????? :
        _3870_ = 8'b10111001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????? :
        _3870_ = 8'b01010111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????? :
        _3870_ = 8'b00110101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????? :
        _3870_ = 8'b01100001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????? :
        _3870_ = 8'b00001110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????? :
        _3870_ = 8'b11110110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????? :
        _3870_ = 8'b00000011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????? :
        _3870_ = 8'b01001000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????? :
        _3870_ = 8'b01100110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????? :
        _3870_ = 8'b10110101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????? :
        _3870_ = 8'b00111110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????? :
        _3870_ = 8'b01110000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????? :
        _3870_ = 8'b10001010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????? :
        _3870_ = 8'b10001011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????? :
        _3870_ = 8'b10111101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????? :
        _3870_ = 8'b01001011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????? :
        _3870_ = 8'b00011111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????? :
        _3870_ = 8'b01110100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????? :
        _3870_ = 8'b11011101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????? :
        _3870_ = 8'b11101000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????? :
        _3870_ = 8'b11000110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????? :
        _3870_ = 8'b10110100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????? :
        _3870_ = 8'b10100110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????? :
        _3870_ = 8'b00011100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????? :
        _3870_ = 8'b00101110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????? :
        _3870_ = 8'b00100101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????? :
        _3870_ = 8'b01111000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????? :
        _3870_ = 8'b10111010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????? :
        _3870_ = 8'b00001000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b10101110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b01111010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b01100101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b11101010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b11110100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b01010110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b01101100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b10101001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b01001110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b11010101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b10001101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b01101101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b00110111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b11001000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b11100111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b01111001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b11100100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b10010101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b10010001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b01100010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b10101100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b11010011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b11000010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b01011100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b00100100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b00000110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b01001001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b00001010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b00111010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b00110010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b11100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b11011011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b00001011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b01011110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b11011110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b00010100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b10111000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b11101110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b01000110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b10001000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b10010000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b00101010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b00100010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b11011100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b01001111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b10000001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b01100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b01110011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b00011001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b01011101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b01100100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b00111101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b01111110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b10100111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b11000100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b00010111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b01000100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b10010111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b01011111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b11101100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b00010011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b00001100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b11001101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b11010010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b11110011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b11111111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b00010000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b00100001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b11011010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b10110110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b10111100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b11110101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b00111000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b10011101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b10010010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b10001111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b01000000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b10100011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b01010001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b10101000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b10011111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b00111100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b01010000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b01111111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b00000010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b11111001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b01000101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b10000101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b00110011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b01001101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b01000011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b11111011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b10101010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b11101111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b11010000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b11001111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b01011000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b01001100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b01001010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b00111001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b10111110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b11001011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b01101010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b01011011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b10110001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b11111100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b00100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b11101101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b00000000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b11010001 ;
      256'b????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b01010011 ;
      256'b???????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b10000100 ;
      256'b??????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b00101111 ;
      256'b?????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b11100011 ;
      256'b????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b00101001 ;
      256'b???????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b10110011 ;
      256'b??????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b11010110 ;
      256'b?????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b00111011 ;
      256'b????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b01010010 ;
      256'b???????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b10100000 ;
      256'b??????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b01011010 ;
      256'b?????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b01101110 ;
      256'b????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b00011011 ;
      256'b???????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b00011010 ;
      256'b??????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b00101100 ;
      256'b?????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b10000011 ;
      256'b????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b00001001 ;
      256'b???????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b01110101 ;
      256'b??????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b10110010 ;
      256'b?????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b00100111 ;
      256'b????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b11101011 ;
      256'b???????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b11100010 ;
      256'b??????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b10000000 ;
      256'b?????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b00010010 ;
      256'b????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b00000111 ;
      256'b???????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b10011010 ;
      256'b??????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b00000101 ;
      256'b?????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b10010110 ;
      256'b????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b00011000 ;
      256'b???????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b11000011 ;
      256'b??????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b00100011 ;
      256'b?????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b11000111 ;
      256'b????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b00000100 ;
      256'b???????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b00010101 ;
      256'b??????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b00110001 ;
      256'b?????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b11011000 ;
      256'b????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b01110001 ;
      256'b???????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b11110001 ;
      256'b??????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b11100101 ;
      256'b?????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b10100101 ;
      256'b????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b00110100 ;
      256'b???????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b11001100 ;
      256'b??????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b11110111 ;
      256'b?????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b00111111 ;
      256'b????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b00110110 ;
      256'b???????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b00100110 ;
      256'b??????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b10010011 ;
      256'b?????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b11111101 ;
      256'b????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b10110111 ;
      256'b???????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b11000000 ;
      256'b??????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b01110010 ;
      256'b?????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b10100100 ;
      256'b????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b10011100 ;
      256'b???????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b10101111 ;
      256'b??????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b10100010 ;
      256'b?????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b11010100 ;
      256'b????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b10101101 ;
      256'b???????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b11110000 ;
      256'b??????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b01000111 ;
      256'b?????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b01011001 ;
      256'b????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b11111010 ;
      256'b???????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b01111101 ;
      256'b??????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b11001001 ;
      256'b?????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b10000010 ;
      256'b????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b11001010 ;
      256'b???????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b01110110 ;
      256'b??????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b10101011 ;
      256'b?????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b11010111 ;
      256'b????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b11111110 ;
      256'b???????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b00101011 ;
      256'b??????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b01100111 ;
      256'b?????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b00000001 ;
      256'b????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b00110000 ;
      256'b???????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b11000101 ;
      256'b??????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b01101111 ;
      256'b?????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b01101011 ;
      256'b????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b11110010 ;
      256'b???1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b01111011 ;
      256'b??1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b01110111 ;
      256'b?1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b01111100 ;
      256'b1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b01100011 ;
      default:
        _3870_ = \t3.t3.s0.out ;
    endcase
  end
  assign _3871_ = state_in[7:0] == 8'b11111111;
  assign _3872_ = state_in[7:0] == 8'b11111110;
  assign _3873_ = state_in[7:0] == 8'b11111101;
  assign _3874_ = state_in[7:0] == 8'b11111100;
  assign _3875_ = state_in[7:0] == 8'b11111011;
  assign _3876_ = state_in[7:0] == 8'b11111010;
  assign _3877_ = state_in[7:0] == 8'b11111001;
  assign _3878_ = state_in[7:0] == 8'b11111000;
  assign _3879_ = state_in[7:0] == 8'b11110111;
  assign _3880_ = state_in[7:0] == 8'b11110110;
  assign _3881_ = state_in[7:0] == 8'b11110101;
  assign _3882_ = state_in[7:0] == 8'b11110100;
  assign _3883_ = state_in[7:0] == 8'b11110011;
  assign _3884_ = state_in[7:0] == 8'b11110010;
  assign _3885_ = state_in[7:0] == 8'b11110001;
  assign _3886_ = state_in[7:0] == 8'b11110000;
  assign _3887_ = state_in[7:0] == 8'b11101111;
  assign _3888_ = state_in[7:0] == 8'b11101110;
  assign _3889_ = state_in[7:0] == 8'b11101101;
  assign _3890_ = state_in[7:0] == 8'b11101100;
  assign _3891_ = state_in[7:0] == 8'b11101011;
  assign _3892_ = state_in[7:0] == 8'b11101010;
  assign _3893_ = state_in[7:0] == 8'b11101001;
  assign _3894_ = state_in[7:0] == 8'b11101000;
  assign _3895_ = state_in[7:0] == 8'b11100111;
  assign _3896_ = state_in[7:0] == 8'b11100110;
  assign _3897_ = state_in[7:0] == 8'b11100101;
  assign _3898_ = state_in[7:0] == 8'b11100100;
  assign _3899_ = state_in[7:0] == 8'b11100011;
  assign _3900_ = state_in[7:0] == 8'b11100010;
  assign _3901_ = state_in[7:0] == 8'b11100001;
  assign _3902_ = state_in[7:0] == 8'b11100000;
  assign _3903_ = state_in[7:0] == 8'b11011111;
  assign _3904_ = state_in[7:0] == 8'b11011110;
  assign _3905_ = state_in[7:0] == 8'b11011101;
  assign _3906_ = state_in[7:0] == 8'b11011100;
  assign _3907_ = state_in[7:0] == 8'b11011011;
  assign _3908_ = state_in[7:0] == 8'b11011010;
  assign _3909_ = state_in[7:0] == 8'b11011001;
  assign _3910_ = state_in[7:0] == 8'b11011000;
  assign _3911_ = state_in[7:0] == 8'b11010111;
  assign _3912_ = state_in[7:0] == 8'b11010110;
  assign _3913_ = state_in[7:0] == 8'b11010101;
  assign _3914_ = state_in[7:0] == 8'b11010100;
  assign _3915_ = state_in[7:0] == 8'b11010011;
  assign _3916_ = state_in[7:0] == 8'b11010010;
  assign _3917_ = state_in[7:0] == 8'b11010001;
  assign _3918_ = state_in[7:0] == 8'b11010000;
  assign _3919_ = state_in[7:0] == 8'b11001111;
  assign _3920_ = state_in[7:0] == 8'b11001110;
  assign _3921_ = state_in[7:0] == 8'b11001101;
  assign _3922_ = state_in[7:0] == 8'b11001100;
  assign _3923_ = state_in[7:0] == 8'b11001011;
  assign _3924_ = state_in[7:0] == 8'b11001010;
  assign _3925_ = state_in[7:0] == 8'b11001001;
  assign _3926_ = state_in[7:0] == 8'b11001000;
  assign _3927_ = state_in[7:0] == 8'b11000111;
  assign _3928_ = state_in[7:0] == 8'b11000110;
  assign _3929_ = state_in[7:0] == 8'b11000101;
  assign _3930_ = state_in[7:0] == 8'b11000100;
  assign _3931_ = state_in[7:0] == 8'b11000011;
  assign _3932_ = state_in[7:0] == 8'b11000010;
  assign _3933_ = state_in[7:0] == 8'b11000001;
  assign _3934_ = state_in[7:0] == 8'b11000000;
  assign _3935_ = state_in[7:0] == 8'b10111111;
  assign _3936_ = state_in[7:0] == 8'b10111110;
  assign _3937_ = state_in[7:0] == 8'b10111101;
  assign _3938_ = state_in[7:0] == 8'b10111100;
  assign _3939_ = state_in[7:0] == 8'b10111011;
  assign _3940_ = state_in[7:0] == 8'b10111010;
  assign _3941_ = state_in[7:0] == 8'b10111001;
  assign _3942_ = state_in[7:0] == 8'b10111000;
  assign _3943_ = state_in[7:0] == 8'b10110111;
  assign _3944_ = state_in[7:0] == 8'b10110110;
  assign _3945_ = state_in[7:0] == 8'b10110101;
  assign _3946_ = state_in[7:0] == 8'b10110100;
  assign _3947_ = state_in[7:0] == 8'b10110011;
  assign _3948_ = state_in[7:0] == 8'b10110010;
  assign _3949_ = state_in[7:0] == 8'b10110001;
  assign _3950_ = state_in[7:0] == 8'b10110000;
  assign _3951_ = state_in[7:0] == 8'b10101111;
  assign _3952_ = state_in[7:0] == 8'b10101110;
  assign _3953_ = state_in[7:0] == 8'b10101101;
  assign _3954_ = state_in[7:0] == 8'b10101100;
  assign _3955_ = state_in[7:0] == 8'b10101011;
  assign _3956_ = state_in[7:0] == 8'b10101010;
  assign _3957_ = state_in[7:0] == 8'b10101001;
  assign _3958_ = state_in[7:0] == 8'b10101000;
  assign _3959_ = state_in[7:0] == 8'b10100111;
  assign _3960_ = state_in[7:0] == 8'b10100110;
  assign _3961_ = state_in[7:0] == 8'b10100101;
  assign _3962_ = state_in[7:0] == 8'b10100100;
  assign _3963_ = state_in[7:0] == 8'b10100011;
  assign _3964_ = state_in[7:0] == 8'b10100010;
  assign _3965_ = state_in[7:0] == 8'b10100001;
  assign _3966_ = state_in[7:0] == 8'b10100000;
  assign _3967_ = state_in[7:0] == 8'b10011111;
  assign _3968_ = state_in[7:0] == 8'b10011110;
  assign _3969_ = state_in[7:0] == 8'b10011101;
  assign _3970_ = state_in[7:0] == 8'b10011100;
  assign _3971_ = state_in[7:0] == 8'b10011011;
  assign _3972_ = state_in[7:0] == 8'b10011010;
  assign _3973_ = state_in[7:0] == 8'b10011001;
  assign _3974_ = state_in[7:0] == 8'b10011000;
  assign _3975_ = state_in[7:0] == 8'b10010111;
  assign _3976_ = state_in[7:0] == 8'b10010110;
  assign _3977_ = state_in[7:0] == 8'b10010101;
  assign _3978_ = state_in[7:0] == 8'b10010100;
  assign _3979_ = state_in[7:0] == 8'b10010011;
  assign _3980_ = state_in[7:0] == 8'b10010010;
  assign _3981_ = state_in[7:0] == 8'b10010001;
  assign _3982_ = state_in[7:0] == 8'b10010000;
  assign _3983_ = state_in[7:0] == 8'b10001111;
  assign _3984_ = state_in[7:0] == 8'b10001110;
  assign _3985_ = state_in[7:0] == 8'b10001101;
  assign _3986_ = state_in[7:0] == 8'b10001100;
  assign _3987_ = state_in[7:0] == 8'b10001011;
  assign _3988_ = state_in[7:0] == 8'b10001010;
  assign _3989_ = state_in[7:0] == 8'b10001001;
  assign _3990_ = state_in[7:0] == 8'b10001000;
  assign _3991_ = state_in[7:0] == 8'b10000111;
  assign _3992_ = state_in[7:0] == 8'b10000110;
  assign _3993_ = state_in[7:0] == 8'b10000101;
  assign _3994_ = state_in[7:0] == 8'b10000100;
  assign _3995_ = state_in[7:0] == 8'b10000011;
  assign _3996_ = state_in[7:0] == 8'b10000010;
  assign _3997_ = state_in[7:0] == 8'b10000001;
  assign _3998_ = state_in[7:0] == 8'b10000000;
  assign _3999_ = state_in[7:0] == 7'b1111111;
  assign _4000_ = state_in[7:0] == 7'b1111110;
  assign _4001_ = state_in[7:0] == 7'b1111101;
  assign _4002_ = state_in[7:0] == 7'b1111100;
  assign _4003_ = state_in[7:0] == 7'b1111011;
  assign _4004_ = state_in[7:0] == 7'b1111010;
  assign _4005_ = state_in[7:0] == 7'b1111001;
  assign _4006_ = state_in[7:0] == 7'b1111000;
  assign _4007_ = state_in[7:0] == 7'b1110111;
  assign _4008_ = state_in[7:0] == 7'b1110110;
  assign _4009_ = state_in[7:0] == 7'b1110101;
  assign _4010_ = state_in[7:0] == 7'b1110100;
  assign _4011_ = state_in[7:0] == 7'b1110011;
  assign _4012_ = state_in[7:0] == 7'b1110010;
  assign _4013_ = state_in[7:0] == 7'b1110001;
  assign _4014_ = state_in[7:0] == 7'b1110000;
  assign _4015_ = state_in[7:0] == 7'b1101111;
  assign _4016_ = state_in[7:0] == 7'b1101110;
  assign _4017_ = state_in[7:0] == 7'b1101101;
  assign _4018_ = state_in[7:0] == 7'b1101100;
  assign _4019_ = state_in[7:0] == 7'b1101011;
  assign _4020_ = state_in[7:0] == 7'b1101010;
  assign _4021_ = state_in[7:0] == 7'b1101001;
  assign _4022_ = state_in[7:0] == 7'b1101000;
  assign _4023_ = state_in[7:0] == 7'b1100111;
  assign _4024_ = state_in[7:0] == 7'b1100110;
  assign _4025_ = state_in[7:0] == 7'b1100101;
  assign _4026_ = state_in[7:0] == 7'b1100100;
  assign _4027_ = state_in[7:0] == 7'b1100011;
  assign _4028_ = state_in[7:0] == 7'b1100010;
  assign _4029_ = state_in[7:0] == 7'b1100001;
  assign _4030_ = state_in[7:0] == 7'b1100000;
  assign _4031_ = state_in[7:0] == 7'b1011111;
  assign _4032_ = state_in[7:0] == 7'b1011110;
  assign _4033_ = state_in[7:0] == 7'b1011101;
  assign _4034_ = state_in[7:0] == 7'b1011100;
  assign _4035_ = state_in[7:0] == 7'b1011011;
  assign _4036_ = state_in[7:0] == 7'b1011010;
  assign _4037_ = state_in[7:0] == 7'b1011001;
  assign _4038_ = state_in[7:0] == 7'b1011000;
  assign _4039_ = state_in[7:0] == 7'b1010111;
  assign _4040_ = state_in[7:0] == 7'b1010110;
  assign _4041_ = state_in[7:0] == 7'b1010101;
  assign _4042_ = state_in[7:0] == 7'b1010100;
  assign _4043_ = state_in[7:0] == 7'b1010011;
  assign _4044_ = state_in[7:0] == 7'b1010010;
  assign _4045_ = state_in[7:0] == 7'b1010001;
  assign _4046_ = state_in[7:0] == 7'b1010000;
  assign _4047_ = state_in[7:0] == 7'b1001111;
  assign _4048_ = state_in[7:0] == 7'b1001110;
  assign _4049_ = state_in[7:0] == 7'b1001101;
  assign _4050_ = state_in[7:0] == 7'b1001100;
  assign _4051_ = state_in[7:0] == 7'b1001011;
  assign _4052_ = state_in[7:0] == 7'b1001010;
  assign _4053_ = state_in[7:0] == 7'b1001001;
  assign _4054_ = state_in[7:0] == 7'b1001000;
  assign _4055_ = state_in[7:0] == 7'b1000111;
  assign _4056_ = state_in[7:0] == 7'b1000110;
  assign _4057_ = state_in[7:0] == 7'b1000101;
  assign _4058_ = state_in[7:0] == 7'b1000100;
  assign _4059_ = state_in[7:0] == 7'b1000011;
  assign _4060_ = state_in[7:0] == 7'b1000010;
  assign _4061_ = state_in[7:0] == 7'b1000001;
  assign _4062_ = state_in[7:0] == 7'b1000000;
  assign _4063_ = state_in[7:0] == 6'b111111;
  assign _4064_ = state_in[7:0] == 6'b111110;
  assign _4065_ = state_in[7:0] == 6'b111101;
  assign _4066_ = state_in[7:0] == 6'b111100;
  assign _4067_ = state_in[7:0] == 6'b111011;
  assign _4068_ = state_in[7:0] == 6'b111010;
  assign _4069_ = state_in[7:0] == 6'b111001;
  assign _4070_ = state_in[7:0] == 6'b111000;
  assign _4071_ = state_in[7:0] == 6'b110111;
  assign _4072_ = state_in[7:0] == 6'b110110;
  assign _4073_ = state_in[7:0] == 6'b110101;
  assign _4074_ = state_in[7:0] == 6'b110100;
  assign _4075_ = state_in[7:0] == 6'b110011;
  assign _4076_ = state_in[7:0] == 6'b110010;
  assign _4077_ = state_in[7:0] == 6'b110001;
  assign _4078_ = state_in[7:0] == 6'b110000;
  assign _4079_ = state_in[7:0] == 6'b101111;
  assign _4080_ = state_in[7:0] == 6'b101110;
  assign _4081_ = state_in[7:0] == 6'b101101;
  assign _4082_ = state_in[7:0] == 6'b101100;
  assign _4083_ = state_in[7:0] == 6'b101011;
  assign _4084_ = state_in[7:0] == 6'b101010;
  assign _4085_ = state_in[7:0] == 6'b101001;
  assign _4086_ = state_in[7:0] == 6'b101000;
  assign _4087_ = state_in[7:0] == 6'b100111;
  assign _4088_ = state_in[7:0] == 6'b100110;
  assign _4089_ = state_in[7:0] == 6'b100101;
  assign _4090_ = state_in[7:0] == 6'b100100;
  assign _4091_ = state_in[7:0] == 6'b100011;
  assign _4092_ = state_in[7:0] == 6'b100010;
  assign _4093_ = state_in[7:0] == 6'b100001;
  assign _4094_ = state_in[7:0] == 6'b100000;
  assign _4095_ = state_in[7:0] == 5'b11111;
  assign _4096_ = state_in[7:0] == 5'b11110;
  assign _4097_ = state_in[7:0] == 5'b11101;
  assign _4098_ = state_in[7:0] == 5'b11100;
  assign _4099_ = state_in[7:0] == 5'b11011;
  assign _4100_ = state_in[7:0] == 5'b11010;
  assign _4101_ = state_in[7:0] == 5'b11001;
  assign _4102_ = state_in[7:0] == 5'b11000;
  assign _4103_ = state_in[7:0] == 5'b10111;
  assign _4104_ = state_in[7:0] == 5'b10110;
  assign _4105_ = state_in[7:0] == 5'b10101;
  assign _4106_ = state_in[7:0] == 5'b10100;
  assign _4107_ = state_in[7:0] == 5'b10011;
  assign _4108_ = state_in[7:0] == 5'b10010;
  assign _4109_ = state_in[7:0] == 5'b10001;
  assign _4110_ = state_in[7:0] == 5'b10000;
  assign _4111_ = state_in[7:0] == 4'b1111;
  assign _4112_ = state_in[7:0] == 4'b1110;
  assign _4113_ = state_in[7:0] == 4'b1101;
  assign _4114_ = state_in[7:0] == 4'b1100;
  assign _4115_ = state_in[7:0] == 4'b1011;
  assign _4116_ = state_in[7:0] == 4'b1010;
  assign _4117_ = state_in[7:0] == 4'b1001;
  assign _4118_ = state_in[7:0] == 4'b1000;
  assign _4119_ = state_in[7:0] == 3'b111;
  assign _4120_ = state_in[7:0] == 3'b110;
  assign _4121_ = state_in[7:0] == 3'b101;
  assign _4122_ = state_in[7:0] == 3'b100;
  assign _4123_ = state_in[7:0] == 2'b11;
  assign _4124_ = state_in[7:0] == 2'b10;
  assign _4125_ = state_in[7:0] == 1'b1;
  assign _4126_ = ! state_in[7:0];
  always @(posedge clk)
      \t3.t3.s4.out <= _4127_;
  wire [255:0] fangyuan32;
  assign fangyuan32 = { _4126_, _4125_, _4124_, _4123_, _4122_, _4121_, _4120_, _4119_, _4118_, _4117_, _4116_, _4115_, _4114_, _4113_, _4112_, _4111_, _4110_, _4109_, _4108_, _4107_, _4106_, _4105_, _4104_, _4103_, _4102_, _4101_, _4100_, _4099_, _4098_, _4097_, _4096_, _4095_, _4094_, _4093_, _4092_, _4091_, _4090_, _4089_, _4088_, _4087_, _4086_, _4085_, _4084_, _4083_, _4082_, _4081_, _4080_, _4079_, _4078_, _4077_, _4076_, _4075_, _4074_, _4073_, _4072_, _4071_, _4070_, _4069_, _4068_, _4067_, _4066_, _4065_, _4064_, _4063_, _4062_, _4061_, _4060_, _4059_, _4058_, _4057_, _4056_, _4055_, _4054_, _4053_, _4052_, _4051_, _4050_, _4049_, _4048_, _4047_, _4046_, _4045_, _4044_, _4043_, _4042_, _4041_, _4040_, _4039_, _4038_, _4037_, _4036_, _4035_, _4034_, _4033_, _4032_, _4031_, _4030_, _4029_, _4028_, _4027_, _4026_, _4025_, _4024_, _4023_, _4022_, _4021_, _4020_, _4019_, _4018_, _4017_, _4016_, _4015_, _4014_, _4013_, _4012_, _4011_, _4010_, _4009_, _4008_, _4007_, _4006_, _4005_, _4004_, _4003_, _4002_, _4001_, _4000_, _3999_, _3998_, _3997_, _3996_, _3995_, _3994_, _3993_, _3992_, _3991_, _3990_, _3989_, _3988_, _3987_, _3986_, _3985_, _3984_, _3983_, _3982_, _3981_, _3980_, _3979_, _3978_, _3977_, _3976_, _3975_, _3974_, _3973_, _3972_, _3971_, _3970_, _3969_, _3968_, _3967_, _3966_, _3965_, _3964_, _3963_, _3962_, _3961_, _3960_, _3959_, _3958_, _3957_, _3956_, _3955_, _3954_, _3953_, _3952_, _3951_, _3950_, _3949_, _3948_, _3947_, _3946_, _3945_, _3944_, _3943_, _3942_, _3941_, _3940_, _3939_, _3938_, _3937_, _3936_, _3935_, _3934_, _3933_, _3932_, _3931_, _3930_, _3929_, _3928_, _3927_, _3926_, _3925_, _3924_, _3923_, _3922_, _3921_, _3920_, _3919_, _3918_, _3917_, _3916_, _3915_, _3914_, _3913_, _3912_, _3911_, _3910_, _3909_, _3908_, _3907_, _3906_, _3905_, _3904_, _3903_, _3902_, _3901_, _3900_, _3899_, _3898_, _3897_, _3896_, _3895_, _3894_, _3893_, _3892_, _3891_, _3890_, _3889_, _3888_, _3887_, _3886_, _3885_, _3884_, _3883_, _3882_, _3881_, _3880_, _3879_, _3878_, _3877_, _3876_, _3875_, _3874_, _3873_, _3872_, _3871_ };

  always @(\t3.t3.s4.out or fangyuan32) begin
    casez (fangyuan32)
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1 :
        _4127_ = 8'b00101100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1? :
        _4127_ = 8'b01101101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?? :
        _4127_ = 8'b10101000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??? :
        _4127_ = 8'b01111011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???? :
        _4127_ = 8'b00011110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????? :
        _4127_ = 8'b01011010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????? :
        _4127_ = 8'b00101001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????? :
        _4127_ = 8'b10000010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????? :
        _4127_ = 8'b11010000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????? :
        _4127_ = 8'b10000100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????? :
        _4127_ = 8'b11010111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????? :
        _4127_ = 8'b01100101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????? :
        _4127_ = 8'b00011010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????? :
        _4127_ = 8'b00001001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????? :
        _4127_ = 8'b01011001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????? :
        _4127_ = 8'b00000011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????? :
        _4127_ = 8'b10100101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????? :
        _4127_ = 8'b01010000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????? :
        _4127_ = 8'b10101010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????? :
        _4127_ = 8'b10000111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????? :
        _4127_ = 8'b11001001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????? :
        _4127_ = 8'b00010101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????? :
        _4127_ = 8'b00111100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????? :
        _4127_ = 8'b00101101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????? :
        _4127_ = 8'b00110011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????? :
        _4127_ = 8'b00000111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????? :
        _4127_ = 8'b10101001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????? :
        _4127_ = 8'b11010010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????? :
        _4127_ = 8'b00100010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????? :
        _4127_ = 8'b00101011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????? :
        _4127_ = 8'b11101011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????? :
        _4127_ = 8'b11011001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????? :
        _4127_ = 8'b00100111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????? :
        _4127_ = 8'b00111010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????? :
        _4127_ = 8'b10011001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????? :
        _4127_ = 8'b00010111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????? :
        _4127_ = 8'b01101001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????? :
        _4127_ = 8'b10101110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????? :
        _4127_ = 8'b01101010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????? :
        _4127_ = 8'b11000010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????? :
        _4127_ = 8'b00011100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????? :
        _4127_ = 8'b11110111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????? :
        _4127_ = 8'b00000110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????? :
        _4127_ = 8'b10010000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????? :
        _4127_ = 8'b11001100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????? :
        _4127_ = 8'b01110001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????? :
        _4127_ = 8'b01111100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????? :
        _4127_ = 8'b11100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????? :
        _4127_ = 8'b00001111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????? :
        _4127_ = 8'b00001101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????? :
        _4127_ = 8'b01100001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????? :
        _4127_ = 8'b10010110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????? :
        _4127_ = 8'b00111110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????? :
        _4127_ = 8'b11101000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????? :
        _4127_ = 8'b10100001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????? :
        _4127_ = 8'b11001011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????? :
        _4127_ = 8'b10010111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????? :
        _4127_ = 8'b01110011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????? :
        _4127_ = 8'b01010111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????? :
        _4127_ = 8'b00111000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????? :
        _4127_ = 8'b01011100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????? :
        _4127_ = 8'b01001010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????? :
        _4127_ = 8'b11110000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????? :
        _4127_ = 8'b01101111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????? :
        _4127_ = 8'b00010000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b01000111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b11110100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b11001010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b11001111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b11110011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b10101100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b11011000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b01001001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b10011100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b10110001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b00000001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b11011010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b01101110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b10001011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b11010101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b11110010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b11010011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b00110001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b00111001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b11000100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b01000011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b10111101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b10011111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b10111000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b01001000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b00001100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b10010010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b00010100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b01110100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b01100100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b11011011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b10101101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b00010110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b10111100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b10100111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b00101000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b01101011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b11000111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b10001100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b00001011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b00111011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b01010100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b01000100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b10100011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b10011110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b00011001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b11000000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b11100110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b00110010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b10111010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b11001000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b01111010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b11111100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b01010101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b10010011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b00101110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b10001000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b00110101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b10111110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b11000011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b00100110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b00011000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b10000001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b10111111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b11111101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b11100101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b00100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b01000010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b10101111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b01110111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b01100011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b11110001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b01110000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b00100001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b00111111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b00000101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b10000000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b01011101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b10100010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b01001011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b00100101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b01111000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b10100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b11111110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b00000100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b11101001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b10001010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b00010001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b01100110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b10011010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b10000110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b11101101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b01001111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b11000101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b10111011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b10000101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b10110000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b10011000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b10010100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b01110010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b01100111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b10001101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b11010100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b10110110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b01111001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b11100011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b01000000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b11000001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b00000000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b10111001 ;
      256'b????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b10100110 ;
      256'b???????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b00010011 ;
      256'b??????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b01011110 ;
      256'b?????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b11011101 ;
      256'b????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b01010010 ;
      256'b???????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b01111101 ;
      256'b??????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b10110111 ;
      256'b?????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b01110110 ;
      256'b????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b10100100 ;
      256'b???????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b01011011 ;
      256'b??????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b10110100 ;
      256'b?????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b11011100 ;
      256'b????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b00110110 ;
      256'b???????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b00110100 ;
      256'b??????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b01011000 ;
      256'b?????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b00011101 ;
      256'b????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b00010010 ;
      256'b???????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b11101010 ;
      256'b??????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b01111111 ;
      256'b?????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b01001110 ;
      256'b????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b11001101 ;
      256'b???????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b11011111 ;
      256'b??????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b00011011 ;
      256'b?????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b00100100 ;
      256'b????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b00001110 ;
      256'b???????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b00101111 ;
      256'b??????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b00001010 ;
      256'b?????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b00110111 ;
      256'b????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b00110000 ;
      256'b???????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b10011101 ;
      256'b??????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b01000110 ;
      256'b?????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b10010101 ;
      256'b????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b00001000 ;
      256'b???????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b00101010 ;
      256'b??????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b01100010 ;
      256'b?????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b10101011 ;
      256'b????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b11100010 ;
      256'b???????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b11111001 ;
      256'b??????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b11010001 ;
      256'b?????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b01010001 ;
      256'b????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b01101000 ;
      256'b???????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b10000011 ;
      256'b??????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b11110101 ;
      256'b?????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b01111110 ;
      256'b????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b01101100 ;
      256'b???????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b01001100 ;
      256'b??????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b00111101 ;
      256'b?????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b11100001 ;
      256'b????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b01110101 ;
      256'b???????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b10011011 ;
      256'b??????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b11100100 ;
      256'b?????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b01010011 ;
      256'b????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b00100011 ;
      256'b???????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b01000101 ;
      256'b??????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b01011111 ;
      256'b?????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b10110011 ;
      256'b????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b01000001 ;
      256'b???????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b11111011 ;
      256'b??????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b10001110 ;
      256'b?????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b10110010 ;
      256'b????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b11101111 ;
      256'b???????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b11111010 ;
      256'b??????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b10001001 ;
      256'b?????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b00011111 ;
      256'b????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b10001111 ;
      256'b???????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b11101100 ;
      256'b??????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b01001101 ;
      256'b?????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b10110101 ;
      256'b????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b11100111 ;
      256'b???????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b01010110 ;
      256'b??????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b11001110 ;
      256'b?????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b00000010 ;
      256'b????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b01100000 ;
      256'b???????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b10010001 ;
      256'b??????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b11011110 ;
      256'b?????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b11010110 ;
      256'b????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b11111111 ;
      256'b???1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b11110110 ;
      256'b??1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b11101110 ;
      256'b?1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b11111000 ;
      256'b1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b11000110 ;
      default:
        _4127_ = \t3.t3.s4.out ;
    endcase
  end
  wire [31:0] fangyuan33;
  assign fangyuan33 = { \t0.t0.s4.out , \t0.t0.s0.out , \t0.t0.s0.out , p00[7:0] };
  wire [31:0] fangyuan34;
  assign fangyuan34 = { p11[31:24], \t1.t1.s4.out , \t1.t1.s0.out , \t1.t1.s0.out };

  assign _4128_ = fangyuan33 ^ fangyuan34;
  wire [31:0] fangyuan35;
  assign fangyuan35 = { \t2.t2.s0.out , p22[23:16], \t2.t2.s4.out , \t2.t2.s0.out };

  assign _4129_ = _4128_ ^ fangyuan35;
  wire [31:0] fangyuan36;
  assign fangyuan36 = { \t3.t3.s0.out , \t3.t3.s0.out , p33[15:8], \t3.t3.s4.out };

  assign _4130_ = _4129_ ^ fangyuan36;
  assign z0 = _4130_ ^ key[127:96];
  wire [31:0] fangyuan37;
  assign fangyuan37 = { \t0.t3.s0.out , \t0.t3.s0.out , p03[15:8], \t0.t3.s4.out };
  wire [31:0] fangyuan38;
  assign fangyuan38 = { \t1.t0.s4.out , \t1.t0.s0.out , \t1.t0.s0.out , p10[7:0] };

  assign _4131_ = fangyuan37 ^ fangyuan38;
  wire [31:0] fangyuan39;
  assign fangyuan39 = { p21[31:24], \t2.t1.s4.out , \t2.t1.s0.out , \t2.t1.s0.out };

  assign _4132_ = _4131_ ^ fangyuan39;
  wire [31:0] fangyuan40;
  assign fangyuan40 = { \t3.t2.s0.out , p32[23:16], \t3.t2.s4.out , \t3.t2.s0.out };

  assign _4133_ = _4132_ ^ fangyuan40;
  assign z1 = _4133_ ^ key[95:64];
  wire [31:0] fangyuan41;
  assign fangyuan41 = { \t2.t0.s4.out , \t2.t0.s0.out , \t2.t0.s0.out , p20[7:0] };

  assign _4134_ = _4136_ ^ fangyuan41;
  wire [31:0] fangyuan42;
  assign fangyuan42 = { p31[31:24], \t3.t1.s4.out , \t3.t1.s0.out , \t3.t1.s0.out };

  assign _4135_ = _4134_ ^ fangyuan42;
  assign z2 = _4135_ ^ key[63:32];
  wire [31:0] fangyuan43;
  assign fangyuan43 = { \t0.t2.s0.out , p02[23:16], \t0.t2.s4.out , \t0.t2.s0.out };
  wire [31:0] fangyuan44;
  assign fangyuan44 = { \t1.t3.s0.out , \t1.t3.s0.out , p13[15:8], \t1.t3.s4.out };

  assign _4136_ = fangyuan43 ^ fangyuan44;
  wire [31:0] fangyuan45;
  assign fangyuan45 = { p01[31:24], \t0.t1.s4.out , \t0.t1.s0.out , \t0.t1.s0.out };
  wire [31:0] fangyuan46;
  assign fangyuan46 = { \t1.t2.s0.out , p12[23:16], \t1.t2.s4.out , \t1.t2.s0.out };

  assign _4137_ = fangyuan45 ^ fangyuan46;
  wire [31:0] fangyuan47;
  assign fangyuan47 = { \t2.t3.s0.out , \t2.t3.s0.out , p23[15:8], \t2.t3.s4.out };

  assign _4138_ = _4137_ ^ fangyuan47;
  wire [31:0] fangyuan48;
  assign fangyuan48 = { \t3.t0.s4.out , \t3.t0.s0.out , \t3.t0.s0.out , p30[7:0] };

  assign _4139_ = _4138_ ^ fangyuan48;
  assign z3 = _4139_ ^ key[31:0];
  assign k0 = key[127:96];
  assign k1 = key[95:64];
  assign k2 = key[63:32];
  assign k3 = key[31:0];
  assign p00[31:8] = { \t0.t0.s4.out , \t0.t0.s0.out , \t0.t0.s0.out };
  assign p01[23:0] = { \t0.t1.s4.out , \t0.t1.s0.out , \t0.t1.s0.out };
  assign p02[31:24] = { \t0.t2.s0.out };
  assign p02[15:0] = { \t0.t2.s4.out, \t0.t2.s0.out };
  assign p03[31:16] = { \t0.t3.s0.out, \t0.t3.s0.out };
  assign p03[7:0] = { \t0.t3.s4.out };
  assign p10[31:8] = { \t1.t0.s4.out , \t1.t0.s0.out , \t1.t0.s0.out };
  assign p11[23:0] = { \t1.t1.s4.out , \t1.t1.s0.out , \t1.t1.s0.out };
  assign p12[31:24] = { \t1.t2.s0.out };
  assign p12[15:0] = { \t1.t2.s4.out, \t1.t2.s0.out };
  assign p13[31:16] = { \t1.t3.s0.out, \t1.t3.s0.out };
  assign p13[7:0] = { \t1.t3.s4.out };
  assign p20[31:8] = { \t2.t0.s4.out , \t2.t0.s0.out , \t2.t0.s0.out };
  assign p21[23:0] = { \t2.t1.s4.out , \t2.t1.s0.out , \t2.t1.s0.out };
  assign p22[31:24] = { \t2.t2.s0.out };
  assign p22[15:0] = { \t2.t2.s4.out, \t2.t2.s0.out };
  assign p23[31:16] = { \t2.t3.s0.out, \t2.t3.s0.out };
  assign p23[7:0] = { \t2.t3.s4.out };
  assign p30[31:8] = { \t3.t0.s4.out , \t3.t0.s0.out , \t3.t0.s0.out };
  assign p31[23:0] = { \t3.t1.s4.out , \t3.t1.s0.out , \t3.t1.s0.out };
  assign p32[31:24] = { \t3.t2.s0.out };
  assign p32[15:0] = { \t3.t2.s4.out, \t3.t2.s0.out };
  assign p33[31:16] = { \t3.t3.s0.out, \t3.t3.s0.out };
  assign p33[7:0] = { \t3.t3.s4.out };
  assign s0 = state_in[127:96];
  assign s1 = state_in[95:64];
  assign s2 = state_in[63:32];
  assign s3 = state_in[31:0];
  assign \t0.b0 = state_in[127:120];
  assign \t0.b1 = state_in[119:112];
  assign \t0.b2 = state_in[111:104];
  assign \t0.b3 = state_in[103:96];
  assign \t0.clk = clk;
  assign \t0.p0 = { \t0.t0.s4.out , \t0.t0.s0.out , \t0.t0.s0.out , p00[7:0] };
  assign \t0.p1 = { p01[31:24], \t0.t1.s4.out , \t0.t1.s0.out , \t0.t1.s0.out };
  assign \t0.p2 = { \t0.t2.s0.out , p02[23:16], \t0.t2.s4.out , \t0.t2.s0.out };
  assign \t0.p3 = { \t0.t3.s0.out , \t0.t3.s0.out , p03[15:8], \t0.t3.s4.out };
  assign \t0.state = state_in[127:96];
  assign \t0.t0.clk = clk;
  assign \t0.t0.in = state_in[127:120];
  assign \t0.t0.out = { \t0.t0.s0.out , \t0.t0.s0.out , p00[7:0], \t0.t0.s4.out };
  assign \t0.t0.s0.clk = clk;
  assign \t0.t0.s0.in = state_in[127:120];
  assign \t0.t0.s4.clk = clk;
  assign \t0.t0.s4.in = state_in[127:120];
  assign \t0.t1.clk = clk;
  assign \t0.t1.in = state_in[119:112];
  assign \t0.t1.out = { \t0.t1.s0.out , \t0.t1.s0.out , p01[31:24], \t0.t1.s4.out };
  assign \t0.t1.s0.clk = clk;
  assign \t0.t1.s0.in = state_in[119:112];
  assign \t0.t1.s4.clk = clk;
  assign \t0.t1.s4.in = state_in[119:112];
  assign \t0.t2.clk = clk;
  assign \t0.t2.in = state_in[111:104];
  assign \t0.t2.out = { \t0.t2.s0.out , \t0.t2.s0.out , p02[23:16], \t0.t2.s4.out };
  assign \t0.t2.s0.clk = clk;
  assign \t0.t2.s0.in = state_in[111:104];
  assign \t0.t2.s4.clk = clk;
  assign \t0.t2.s4.in = state_in[111:104];
  assign \t0.t3.clk = clk;
  assign \t0.t3.in = state_in[103:96];
  assign \t0.t3.out = { \t0.t3.s0.out , \t0.t3.s0.out , p03[15:8], \t0.t3.s4.out };
  assign \t0.t3.s0.clk = clk;
  assign \t0.t3.s0.in = state_in[103:96];
  assign \t0.t3.s4.clk = clk;
  assign \t0.t3.s4.in = state_in[103:96];
  assign \t1.b0 = state_in[95:88];
  assign \t1.b1 = state_in[87:80];
  assign \t1.b2 = state_in[79:72];
  assign \t1.b3 = state_in[71:64];
  assign \t1.clk = clk;
  assign \t1.p0 = { \t1.t0.s4.out , \t1.t0.s0.out , \t1.t0.s0.out , p10[7:0] };
  assign \t1.p1 = { p11[31:24], \t1.t1.s4.out , \t1.t1.s0.out , \t1.t1.s0.out };
  assign \t1.p2 = { \t1.t2.s0.out , p12[23:16], \t1.t2.s4.out , \t1.t2.s0.out };
  assign \t1.p3 = { \t1.t3.s0.out , \t1.t3.s0.out , p13[15:8], \t1.t3.s4.out };
  assign \t1.state = state_in[95:64];
  assign \t1.t0.clk = clk;
  assign \t1.t0.in = state_in[95:88];
  assign \t1.t0.out = { \t1.t0.s0.out , \t1.t0.s0.out , p10[7:0], \t1.t0.s4.out };
  assign \t1.t0.s0.clk = clk;
  assign \t1.t0.s0.in = state_in[95:88];
  assign \t1.t0.s4.clk = clk;
  assign \t1.t0.s4.in = state_in[95:88];
  assign \t1.t1.clk = clk;
  assign \t1.t1.in = state_in[87:80];
  assign \t1.t1.out = { \t1.t1.s0.out , \t1.t1.s0.out , p11[31:24], \t1.t1.s4.out };
  assign \t1.t1.s0.clk = clk;
  assign \t1.t1.s0.in = state_in[87:80];
  assign \t1.t1.s4.clk = clk;
  assign \t1.t1.s4.in = state_in[87:80];
  assign \t1.t2.clk = clk;
  assign \t1.t2.in = state_in[79:72];
  assign \t1.t2.out = { \t1.t2.s0.out , \t1.t2.s0.out , p12[23:16], \t1.t2.s4.out };
  assign \t1.t2.s0.clk = clk;
  assign \t1.t2.s0.in = state_in[79:72];
  assign \t1.t2.s4.clk = clk;
  assign \t1.t2.s4.in = state_in[79:72];
  assign \t1.t3.clk = clk;
  assign \t1.t3.in = state_in[71:64];
  assign \t1.t3.out = { \t1.t3.s0.out , \t1.t3.s0.out , p13[15:8], \t1.t3.s4.out };
  assign \t1.t3.s0.clk = clk;
  assign \t1.t3.s0.in = state_in[71:64];
  assign \t1.t3.s4.clk = clk;
  assign \t1.t3.s4.in = state_in[71:64];
  assign \t2.b0 = state_in[63:56];
  assign \t2.b1 = state_in[55:48];
  assign \t2.b2 = state_in[47:40];
  assign \t2.b3 = state_in[39:32];
  assign \t2.clk = clk;
  assign \t2.p0 = { \t2.t0.s4.out , \t2.t0.s0.out , \t2.t0.s0.out , p20[7:0] };
  assign \t2.p1 = { p21[31:24], \t2.t1.s4.out , \t2.t1.s0.out , \t2.t1.s0.out };
  assign \t2.p2 = { \t2.t2.s0.out , p22[23:16], \t2.t2.s4.out , \t2.t2.s0.out };
  assign \t2.p3 = { \t2.t3.s0.out , \t2.t3.s0.out , p23[15:8], \t2.t3.s4.out };
  assign \t2.state = state_in[63:32];
  assign \t2.t0.clk = clk;
  assign \t2.t0.in = state_in[63:56];
  assign \t2.t0.out = { \t2.t0.s0.out , \t2.t0.s0.out , p20[7:0], \t2.t0.s4.out };
  assign \t2.t0.s0.clk = clk;
  assign \t2.t0.s0.in = state_in[63:56];
  assign \t2.t0.s4.clk = clk;
  assign \t2.t0.s4.in = state_in[63:56];
  assign \t2.t1.clk = clk;
  assign \t2.t1.in = state_in[55:48];
  assign \t2.t1.out = { \t2.t1.s0.out , \t2.t1.s0.out , p21[31:24], \t2.t1.s4.out };
  assign \t2.t1.s0.clk = clk;
  assign \t2.t1.s0.in = state_in[55:48];
  assign \t2.t1.s4.clk = clk;
  assign \t2.t1.s4.in = state_in[55:48];
  assign \t2.t2.clk = clk;
  assign \t2.t2.in = state_in[47:40];
  assign \t2.t2.out = { \t2.t2.s0.out , \t2.t2.s0.out , p22[23:16], \t2.t2.s4.out };
  assign \t2.t2.s0.clk = clk;
  assign \t2.t2.s0.in = state_in[47:40];
  assign \t2.t2.s4.clk = clk;
  assign \t2.t2.s4.in = state_in[47:40];
  assign \t2.t3.clk = clk;
  assign \t2.t3.in = state_in[39:32];
  assign \t2.t3.out = { \t2.t3.s0.out , \t2.t3.s0.out , p23[15:8], \t2.t3.s4.out };
  assign \t2.t3.s0.clk = clk;
  assign \t2.t3.s0.in = state_in[39:32];
  assign \t2.t3.s4.clk = clk;
  assign \t2.t3.s4.in = state_in[39:32];
  assign \t3.b0 = state_in[31:24];
  assign \t3.b1 = state_in[23:16];
  assign \t3.b2 = state_in[15:8];
  assign \t3.b3 = state_in[7:0];
  assign \t3.clk = clk;
  assign \t3.p0 = { \t3.t0.s4.out , \t3.t0.s0.out , \t3.t0.s0.out , p30[7:0] };
  assign \t3.p1 = { p31[31:24], \t3.t1.s4.out , \t3.t1.s0.out , \t3.t1.s0.out };
  assign \t3.p2 = { \t3.t2.s0.out , p32[23:16], \t3.t2.s4.out , \t3.t2.s0.out };
  assign \t3.p3 = { \t3.t3.s0.out , \t3.t3.s0.out , p33[15:8], \t3.t3.s4.out };
  assign \t3.state = state_in[31:0];
  assign \t3.t0.clk = clk;
  assign \t3.t0.in = state_in[31:24];
  assign \t3.t0.out = { \t3.t0.s0.out , \t3.t0.s0.out , p30[7:0], \t3.t0.s4.out };
  assign \t3.t0.s0.clk = clk;
  assign \t3.t0.s0.in = state_in[31:24];
  assign \t3.t0.s4.clk = clk;
  assign \t3.t0.s4.in = state_in[31:24];
  assign \t3.t1.clk = clk;
  assign \t3.t1.in = state_in[23:16];
  assign \t3.t1.out = { \t3.t1.s0.out , \t3.t1.s0.out , p31[31:24], \t3.t1.s4.out };
  assign \t3.t1.s0.clk = clk;
  assign \t3.t1.s0.in = state_in[23:16];
  assign \t3.t1.s4.clk = clk;
  assign \t3.t1.s4.in = state_in[23:16];
  assign \t3.t2.clk = clk;
  assign \t3.t2.in = state_in[15:8];
  assign \t3.t2.out = { \t3.t2.s0.out , \t3.t2.s0.out , p32[23:16], \t3.t2.s4.out };
  assign \t3.t2.s0.clk = clk;
  assign \t3.t2.s0.in = state_in[15:8];
  assign \t3.t2.s4.clk = clk;
  assign \t3.t2.s4.in = state_in[15:8];
  assign \t3.t3.clk = clk;
  assign \t3.t3.in = state_in[7:0];
  assign \t3.t3.out = { \t3.t3.s0.out , \t3.t3.s0.out , p33[15:8], \t3.t3.s4.out };
  assign \t3.t3.s0.clk = clk;
  assign \t3.t3.s0.in = state_in[7:0];
  assign \t3.t3.s4.clk = clk;
  assign \t3.t3.s4.in = state_in[7:0];
endmodule
