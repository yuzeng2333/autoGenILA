module NV_NVDLA_CDP_DP_lut(nvdla_core_clk, nvdla_core_clk_orig, nvdla_core_rstn, dp2lut_X_entry_0, dp2lut_X_entry_1, dp2lut_X_entry_2, dp2lut_X_entry_3, dp2lut_X_entry_4, dp2lut_X_entry_5, dp2lut_X_entry_6, dp2lut_X_entry_7, dp2lut_Xinfo_0, dp2lut_Xinfo_1, dp2lut_Xinfo_2, dp2lut_Xinfo_3, dp2lut_Xinfo_4, dp2lut_Xinfo_5, dp2lut_Xinfo_6, dp2lut_Xinfo_7, dp2lut_Y_entry_0, dp2lut_Y_entry_1, dp2lut_Y_entry_2, dp2lut_Y_entry_3, dp2lut_Y_entry_4, dp2lut_Y_entry_5, dp2lut_Y_entry_6, dp2lut_Y_entry_7, dp2lut_Yinfo_0, dp2lut_Yinfo_1, dp2lut_Yinfo_2, dp2lut_Yinfo_3, dp2lut_Yinfo_4, dp2lut_Yinfo_5, dp2lut_Yinfo_6, dp2lut_Yinfo_7, dp2lut_pvld, int8_en, lut2intp_prdy, nvdla_op_gated_clk_fp16, reg2dp_input_data_type, reg2dp_lut_access_type, reg2dp_lut_addr, reg2dp_lut_data, reg2dp_lut_data_trigger, reg2dp_lut_hybrid_priority, reg2dp_lut_oflow_priority, reg2dp_lut_table_id, reg2dp_lut_uflow_priority, dp2lut_prdy, dp2reg_lut_data, lut2intp_X_data_00, lut2intp_X_data_00_17b, lut2intp_X_data_01, lut2intp_X_data_10, lut2intp_X_data_10_17b, lut2intp_X_data_11, lut2intp_X_data_20, lut2intp_X_data_20_17b, lut2intp_X_data_21, lut2intp_X_data_30, lut2intp_X_data_30_17b, lut2intp_X_data_31, lut2intp_X_data_40, lut2intp_X_data_40_17b, lut2intp_X_data_41, lut2intp_X_data_50, lut2intp_X_data_50_17b, lut2intp_X_data_51, lut2intp_X_data_60, lut2intp_X_data_60_17b, lut2intp_X_data_61, lut2intp_X_data_70, lut2intp_X_data_70_17b, lut2intp_X_data_71, lut2intp_X_info_0, lut2intp_X_info_1, lut2intp_X_info_2, lut2intp_X_info_3, lut2intp_X_info_4, lut2intp_X_info_5, lut2intp_X_info_6, lut2intp_X_info_7, lut2intp_X_sel, lut2intp_Y_sel, lut2intp_pvld);
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4030" *)
  wire [15:0] _0000_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1318" *)
  wire [15:0] _0001_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2318" *)
  wire [15:0] _0002_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2328" *)
  wire [15:0] _0003_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2338" *)
  wire [15:0] _0004_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2348" *)
  wire [15:0] _0005_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2358" *)
  wire [15:0] _0006_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2368" *)
  wire [15:0] _0007_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2378" *)
  wire [15:0] _0008_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2388" *)
  wire [15:0] _0009_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2398" *)
  wire [15:0] _0010_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2408" *)
  wire [15:0] _0011_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1418" *)
  wire [15:0] _0012_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2418" *)
  wire [15:0] _0013_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2428" *)
  wire [15:0] _0014_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2438" *)
  wire [15:0] _0015_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2448" *)
  wire [15:0] _0016_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2458" *)
  wire [15:0] _0017_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2468" *)
  wire [15:0] _0018_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2478" *)
  wire [15:0] _0019_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2488" *)
  wire [15:0] _0020_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2498" *)
  wire [15:0] _0021_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2508" *)
  wire [15:0] _0022_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1428" *)
  wire [15:0] _0023_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2518" *)
  wire [15:0] _0024_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2528" *)
  wire [15:0] _0025_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2538" *)
  wire [15:0] _0026_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2548" *)
  wire [15:0] _0027_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2558" *)
  wire [15:0] _0028_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2568" *)
  wire [15:0] _0029_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2578" *)
  wire [15:0] _0030_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2588" *)
  wire [15:0] _0031_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2598" *)
  wire [15:0] _0032_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2608" *)
  wire [15:0] _0033_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1438" *)
  wire [15:0] _0034_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2618" *)
  wire [15:0] _0035_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2628" *)
  wire [15:0] _0036_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2638" *)
  wire [15:0] _0037_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2648" *)
  wire [15:0] _0038_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2658" *)
  wire [15:0] _0039_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2668" *)
  wire [15:0] _0040_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2678" *)
  wire [15:0] _0041_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2688" *)
  wire [15:0] _0042_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2698" *)
  wire [15:0] _0043_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2708" *)
  wire [15:0] _0044_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1448" *)
  wire [15:0] _0045_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2718" *)
  wire [15:0] _0046_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2728" *)
  wire [15:0] _0047_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2738" *)
  wire [15:0] _0048_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2748" *)
  wire [15:0] _0049_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2758" *)
  wire [15:0] _0050_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2768" *)
  wire [15:0] _0051_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2778" *)
  wire [15:0] _0052_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2788" *)
  wire [15:0] _0053_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2798" *)
  wire [15:0] _0054_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2808" *)
  wire [15:0] _0055_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1458" *)
  wire [15:0] _0056_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2818" *)
  wire [15:0] _0057_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2828" *)
  wire [15:0] _0058_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2838" *)
  wire [15:0] _0059_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2848" *)
  wire [15:0] _0060_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2858" *)
  wire [15:0] _0061_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2868" *)
  wire [15:0] _0062_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2878" *)
  wire [15:0] _0063_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2888" *)
  wire [15:0] _0064_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2898" *)
  wire [15:0] _0065_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2908" *)
  wire [15:0] _0066_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1468" *)
  wire [15:0] _0067_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2918" *)
  wire [15:0] _0068_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2928" *)
  wire [15:0] _0069_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2938" *)
  wire [15:0] _0070_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2948" *)
  wire [15:0] _0071_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2958" *)
  wire [15:0] _0072_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2968" *)
  wire [15:0] _0073_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2978" *)
  wire [15:0] _0074_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2988" *)
  wire [15:0] _0075_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2998" *)
  wire [15:0] _0076_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3008" *)
  wire [15:0] _0077_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1478" *)
  wire [15:0] _0078_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3018" *)
  wire [15:0] _0079_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3028" *)
  wire [15:0] _0080_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3038" *)
  wire [15:0] _0081_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3048" *)
  wire [15:0] _0082_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3058" *)
  wire [15:0] _0083_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3068" *)
  wire [15:0] _0084_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3078" *)
  wire [15:0] _0085_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3088" *)
  wire [15:0] _0086_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3098" *)
  wire [15:0] _0087_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3108" *)
  wire [15:0] _0088_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1488" *)
  wire [15:0] _0089_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3118" *)
  wire [15:0] _0090_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3128" *)
  wire [15:0] _0091_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3138" *)
  wire [15:0] _0092_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3148" *)
  wire [15:0] _0093_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3158" *)
  wire [15:0] _0094_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3168" *)
  wire [15:0] _0095_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3178" *)
  wire [15:0] _0096_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3188" *)
  wire [15:0] _0097_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3198" *)
  wire [15:0] _0098_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3208" *)
  wire [15:0] _0099_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1498" *)
  wire [15:0] _0100_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3218" *)
  wire [15:0] _0101_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3228" *)
  wire [15:0] _0102_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3238" *)
  wire [15:0] _0103_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3248" *)
  wire [15:0] _0104_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3258" *)
  wire [15:0] _0105_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3268" *)
  wire [15:0] _0106_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3278" *)
  wire [15:0] _0107_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3288" *)
  wire [15:0] _0108_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3298" *)
  wire [15:0] _0109_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3308" *)
  wire [15:0] _0110_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1508" *)
  wire [15:0] _0111_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1328" *)
  wire [15:0] _0112_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3318" *)
  wire [15:0] _0113_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3328" *)
  wire [15:0] _0114_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3338" *)
  wire [15:0] _0115_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3348" *)
  wire [15:0] _0116_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3358" *)
  wire [15:0] _0117_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3368" *)
  wire [15:0] _0118_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3378" *)
  wire [15:0] _0119_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3388" *)
  wire [15:0] _0120_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3398" *)
  wire [15:0] _0121_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3408" *)
  wire [15:0] _0122_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1518" *)
  wire [15:0] _0123_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3418" *)
  wire [15:0] _0124_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3428" *)
  wire [15:0] _0125_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3438" *)
  wire [15:0] _0126_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3448" *)
  wire [15:0] _0127_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3458" *)
  wire [15:0] _0128_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3468" *)
  wire [15:0] _0129_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3478" *)
  wire [15:0] _0130_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3488" *)
  wire [15:0] _0131_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3498" *)
  wire [15:0] _0132_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3508" *)
  wire [15:0] _0133_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1528" *)
  wire [15:0] _0134_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3518" *)
  wire [15:0] _0135_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3528" *)
  wire [15:0] _0136_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3538" *)
  wire [15:0] _0137_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3548" *)
  wire [15:0] _0138_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3558" *)
  wire [15:0] _0139_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3568" *)
  wire [15:0] _0140_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3578" *)
  wire [15:0] _0141_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3588" *)
  wire [15:0] _0142_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3598" *)
  wire [15:0] _0143_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3608" *)
  wire [15:0] _0144_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1538" *)
  wire [15:0] _0145_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3618" *)
  wire [15:0] _0146_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3628" *)
  wire [15:0] _0147_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3638" *)
  wire [15:0] _0148_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3648" *)
  wire [15:0] _0149_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3658" *)
  wire [15:0] _0150_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3668" *)
  wire [15:0] _0151_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3678" *)
  wire [15:0] _0152_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3688" *)
  wire [15:0] _0153_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3698" *)
  wire [15:0] _0154_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3708" *)
  wire [15:0] _0155_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1548" *)
  wire [15:0] _0156_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3718" *)
  wire [15:0] _0157_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3728" *)
  wire [15:0] _0158_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3738" *)
  wire [15:0] _0159_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3748" *)
  wire [15:0] _0160_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3758" *)
  wire [15:0] _0161_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3768" *)
  wire [15:0] _0162_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3778" *)
  wire [15:0] _0163_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3788" *)
  wire [15:0] _0164_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3798" *)
  wire [15:0] _0165_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3808" *)
  wire [15:0] _0166_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1558" *)
  wire [15:0] _0167_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3818" *)
  wire [15:0] _0168_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3828" *)
  wire [15:0] _0169_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3838" *)
  wire [15:0] _0170_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3848" *)
  wire [15:0] _0171_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3858" *)
  wire [15:0] _0172_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3868" *)
  wire [15:0] _0173_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3878" *)
  wire [15:0] _0174_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1568" *)
  wire [15:0] _0175_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1578" *)
  wire [15:0] _0176_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1588" *)
  wire [15:0] _0177_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1598" *)
  wire [15:0] _0178_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1608" *)
  wire [15:0] _0179_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1338" *)
  wire [15:0] _0180_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1618" *)
  wire [15:0] _0181_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1628" *)
  wire [15:0] _0182_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1638" *)
  wire [15:0] _0183_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1648" *)
  wire [15:0] _0184_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1658" *)
  wire [15:0] _0185_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1668" *)
  wire [15:0] _0186_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1678" *)
  wire [15:0] _0187_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1688" *)
  wire [15:0] _0188_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1698" *)
  wire [15:0] _0189_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1708" *)
  wire [15:0] _0190_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1348" *)
  wire [15:0] _0191_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1718" *)
  wire [15:0] _0192_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1728" *)
  wire [15:0] _0193_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1738" *)
  wire [15:0] _0194_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1748" *)
  wire [15:0] _0195_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1758" *)
  wire [15:0] _0196_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1768" *)
  wire [15:0] _0197_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1778" *)
  wire [15:0] _0198_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1788" *)
  wire [15:0] _0199_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1798" *)
  wire [15:0] _0200_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1808" *)
  wire [15:0] _0201_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1358" *)
  wire [15:0] _0202_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1818" *)
  wire [15:0] _0203_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1828" *)
  wire [15:0] _0204_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1838" *)
  wire [15:0] _0205_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1848" *)
  wire [15:0] _0206_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1858" *)
  wire [15:0] _0207_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1868" *)
  wire [15:0] _0208_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1878" *)
  wire [15:0] _0209_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1888" *)
  wire [15:0] _0210_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1898" *)
  wire [15:0] _0211_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1908" *)
  wire [15:0] _0212_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1368" *)
  wire [15:0] _0213_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1918" *)
  wire [15:0] _0214_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1928" *)
  wire [15:0] _0215_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1938" *)
  wire [15:0] _0216_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1948" *)
  wire [15:0] _0217_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1958" *)
  wire [15:0] _0218_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1968" *)
  wire [15:0] _0219_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1978" *)
  wire [15:0] _0220_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1988" *)
  wire [15:0] _0221_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1998" *)
  wire [15:0] _0222_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2008" *)
  wire [15:0] _0223_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1378" *)
  wire [15:0] _0224_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2018" *)
  wire [15:0] _0225_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2028" *)
  wire [15:0] _0226_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2038" *)
  wire [15:0] _0227_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2048" *)
  wire [15:0] _0228_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2058" *)
  wire [15:0] _0229_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2068" *)
  wire [15:0] _0230_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2078" *)
  wire [15:0] _0231_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2088" *)
  wire [15:0] _0232_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2098" *)
  wire [15:0] _0233_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2108" *)
  wire [15:0] _0234_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1388" *)
  wire [15:0] _0235_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2118" *)
  wire [15:0] _0236_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2128" *)
  wire [15:0] _0237_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2138" *)
  wire [15:0] _0238_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2148" *)
  wire [15:0] _0239_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2158" *)
  wire [15:0] _0240_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2168" *)
  wire [15:0] _0241_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2178" *)
  wire [15:0] _0242_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2188" *)
  wire [15:0] _0243_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2198" *)
  wire [15:0] _0244_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2208" *)
  wire [15:0] _0245_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1398" *)
  wire [15:0] _0246_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2218" *)
  wire [15:0] _0247_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2228" *)
  wire [15:0] _0248_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2238" *)
  wire [15:0] _0249_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2248" *)
  wire [15:0] _0250_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2258" *)
  wire [15:0] _0251_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2268" *)
  wire [15:0] _0252_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2278" *)
  wire [15:0] _0253_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2288" *)
  wire [15:0] _0254_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2298" *)
  wire [15:0] _0255_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2308" *)
  wire [15:0] _0256_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1408" *)
  wire [15:0] _0257_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:16750" *)
  wire _0258_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:16106" *)
  wire [7:0] _0259_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:16655" *)
  wire [7:0] _0260_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4945" *)
  wire [15:0] _0261_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4945" *)
  wire [15:0] _0262_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5228" *)
  wire [15:0] _0263_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5228" *)
  wire [15:0] _0264_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5511" *)
  wire [15:0] _0265_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5511" *)
  wire [15:0] _0266_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5794" *)
  wire [15:0] _0267_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5794" *)
  wire [15:0] _0268_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6077" *)
  wire [15:0] _0269_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6077" *)
  wire [15:0] _0270_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6360" *)
  wire [15:0] _0271_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6360" *)
  wire [15:0] _0272_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6643" *)
  wire [15:0] _0273_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6643" *)
  wire [15:0] _0274_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6926" *)
  wire [15:0] _0275_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6926" *)
  wire [15:0] _0276_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:15618" *)
  wire [17:0] _0277_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:15679" *)
  wire [17:0] _0278_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:15740" *)
  wire [17:0] _0279_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:15801" *)
  wire [17:0] _0280_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:15862" *)
  wire [17:0] _0281_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:15923" *)
  wire [17:0] _0282_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:15984" *)
  wire [17:0] _0283_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:16045" *)
  wire [17:0] _0284_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7210" *)
  wire [15:0] _0285_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7210" *)
  wire [15:0] _0286_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8261" *)
  wire [15:0] _0287_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8261" *)
  wire [15:0] _0288_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9312" *)
  wire [15:0] _0289_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9312" *)
  wire [15:0] _0290_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10363" *)
  wire [15:0] _0291_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10363" *)
  wire [15:0] _0292_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11414" *)
  wire [15:0] _0293_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11414" *)
  wire [15:0] _0294_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12465" *)
  wire [15:0] _0295_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12465" *)
  wire [15:0] _0296_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13516" *)
  wire [15:0] _0297_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13516" *)
  wire [15:0] _0298_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14567" *)
  wire [15:0] _0299_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14567" *)
  wire [15:0] _0300_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:16167" *)
  wire [17:0] _0301_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:16228" *)
  wire [17:0] _0302_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:16289" *)
  wire [17:0] _0303_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:16350" *)
  wire [17:0] _0304_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:16411" *)
  wire [17:0] _0305_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:16472" *)
  wire [17:0] _0306_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:16533" *)
  wire [17:0] _0307_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:16594" *)
  wire [17:0] _0308_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:16740" *)
  wire _0309_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3891" *)
  wire [15:0] _0310_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:667" *)
  wire [15:0] _0311_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:767" *)
  wire [15:0] _0312_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:777" *)
  wire [15:0] _0313_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:787" *)
  wire [15:0] _0314_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:797" *)
  wire [15:0] _0315_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:807" *)
  wire [15:0] _0316_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:817" *)
  wire [15:0] _0317_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:827" *)
  wire [15:0] _0318_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:837" *)
  wire [15:0] _0319_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:847" *)
  wire [15:0] _0320_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:857" *)
  wire [15:0] _0321_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:677" *)
  wire [15:0] _0322_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:867" *)
  wire [15:0] _0323_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:877" *)
  wire [15:0] _0324_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:887" *)
  wire [15:0] _0325_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:897" *)
  wire [15:0] _0326_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:907" *)
  wire [15:0] _0327_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:917" *)
  wire [15:0] _0328_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:927" *)
  wire [15:0] _0329_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:937" *)
  wire [15:0] _0330_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:947" *)
  wire [15:0] _0331_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:957" *)
  wire [15:0] _0332_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:687" *)
  wire [15:0] _0333_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:967" *)
  wire [15:0] _0334_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:977" *)
  wire [15:0] _0335_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:987" *)
  wire [15:0] _0336_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:997" *)
  wire [15:0] _0337_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1007" *)
  wire [15:0] _0338_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1017" *)
  wire [15:0] _0339_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1027" *)
  wire [15:0] _0340_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1037" *)
  wire [15:0] _0341_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1047" *)
  wire [15:0] _0342_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1057" *)
  wire [15:0] _0343_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:697" *)
  wire [15:0] _0344_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1067" *)
  wire [15:0] _0345_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1077" *)
  wire [15:0] _0346_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1087" *)
  wire [15:0] _0347_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1097" *)
  wire [15:0] _0348_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1107" *)
  wire [15:0] _0349_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1117" *)
  wire [15:0] _0350_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1127" *)
  wire [15:0] _0351_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1137" *)
  wire [15:0] _0352_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1147" *)
  wire [15:0] _0353_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1157" *)
  wire [15:0] _0354_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:707" *)
  wire [15:0] _0355_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1167" *)
  wire [15:0] _0356_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1177" *)
  wire [15:0] _0357_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1187" *)
  wire [15:0] _0358_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1197" *)
  wire [15:0] _0359_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1207" *)
  wire [15:0] _0360_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1217" *)
  wire [15:0] _0361_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1227" *)
  wire [15:0] _0362_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1237" *)
  wire [15:0] _0363_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1247" *)
  wire [15:0] _0364_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1257" *)
  wire [15:0] _0365_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:717" *)
  wire [15:0] _0366_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1267" *)
  wire [15:0] _0367_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1277" *)
  wire [15:0] _0368_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1287" *)
  wire [15:0] _0369_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1297" *)
  wire [15:0] _0370_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1307" *)
  wire [15:0] _0371_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:727" *)
  wire [15:0] _0372_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:737" *)
  wire [15:0] _0373_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:747" *)
  wire [15:0] _0374_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:757" *)
  wire [15:0] _0375_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4630" *)
  wire _0376_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4650" *)
  wire _0377_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4670" *)
  wire _0378_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4690" *)
  wire _0379_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4774" *)
  wire _0380_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4794" *)
  wire _0381_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4814" *)
  wire _0382_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4834" *)
  wire _0383_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1001" *)
  wire _0384_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10368" *)
  wire _0385_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11419" *)
  wire _0386_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11419" *)
  wire _0387_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12470" *)
  wire _0388_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1322" *)
  wire _0389_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13521" *)
  wire _0390_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14572" *)
  wire _0391_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4950" *)
  wire _0392_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5233" *)
  wire _0393_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5516" *)
  wire _0394_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5799" *)
  wire _0395_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6082" *)
  wire _0396_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6365" *)
  wire _0397_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6648" *)
  wire _0398_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6931" *)
  wire _0399_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7215" *)
  wire _0400_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8266" *)
  wire _0401_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9317" *)
  wire _0402_;
  wire _0403_;
  wire _0404_;
  wire _0405_;
  wire _0406_;
  wire _0407_;
  wire _0408_;
  wire _0409_;
  wire _0410_;
  wire _0411_;
  wire _0412_;
  wire _0413_;
  wire _0414_;
  wire _0415_;
  wire _0416_;
  wire _0417_;
  wire _0418_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1002" *)
  wire _0419_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1012" *)
  wire _0420_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1022" *)
  wire _0421_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1032" *)
  wire _0422_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1042" *)
  wire _0423_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1052" *)
  wire _0424_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1062" *)
  wire _0425_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1072" *)
  wire _0426_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1082" *)
  wire _0427_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1092" *)
  wire _0428_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1102" *)
  wire _0429_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1112" *)
  wire _0430_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1122" *)
  wire _0431_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1132" *)
  wire _0432_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1142" *)
  wire _0433_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1152" *)
  wire _0434_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1162" *)
  wire _0435_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1172" *)
  wire _0436_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1182" *)
  wire _0437_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1192" *)
  wire _0438_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1202" *)
  wire _0439_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1212" *)
  wire _0440_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1222" *)
  wire _0441_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1232" *)
  wire _0442_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1242" *)
  wire _0443_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1252" *)
  wire _0444_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1262" *)
  wire _0445_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1272" *)
  wire _0446_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1282" *)
  wire _0447_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1292" *)
  wire _0448_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1302" *)
  wire _0449_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1312" *)
  wire _0450_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1323" *)
  wire _0451_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1333" *)
  wire _0452_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1343" *)
  wire _0453_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1353" *)
  wire _0454_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1363" *)
  wire _0455_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1373" *)
  wire _0456_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1383" *)
  wire _0457_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1393" *)
  wire _0458_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1403" *)
  wire _0459_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1413" *)
  wire _0460_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1423" *)
  wire _0461_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1433" *)
  wire _0462_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1443" *)
  wire _0463_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1453" *)
  wire _0464_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1463" *)
  wire _0465_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1473" *)
  wire _0466_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1483" *)
  wire _0467_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1493" *)
  wire _0468_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1503" *)
  wire _0469_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1513" *)
  wire _0470_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1523" *)
  wire _0471_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1533" *)
  wire _0472_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1543" *)
  wire _0473_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1553" *)
  wire _0474_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1563" *)
  wire _0475_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1573" *)
  wire _0476_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1583" *)
  wire _0477_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1593" *)
  wire _0478_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1603" *)
  wire _0479_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1613" *)
  wire _0480_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1623" *)
  wire _0481_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1633" *)
  wire _0482_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1643" *)
  wire _0483_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1973" *)
  wire _0484_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1983" *)
  wire _0485_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1993" *)
  wire _0486_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2003" *)
  wire _0487_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2013" *)
  wire _0488_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2023" *)
  wire _0489_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2033" *)
  wire _0490_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2043" *)
  wire _0491_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2053" *)
  wire _0492_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2063" *)
  wire _0493_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2073" *)
  wire _0494_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2083" *)
  wire _0495_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2093" *)
  wire _0496_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2103" *)
  wire _0497_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2113" *)
  wire _0498_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2123" *)
  wire _0499_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2133" *)
  wire _0500_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2143" *)
  wire _0501_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2153" *)
  wire _0502_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2163" *)
  wire _0503_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2173" *)
  wire _0504_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2183" *)
  wire _0505_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2193" *)
  wire _0506_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2203" *)
  wire _0507_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2213" *)
  wire _0508_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2223" *)
  wire _0509_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2233" *)
  wire _0510_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2243" *)
  wire _0511_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2253" *)
  wire _0512_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2263" *)
  wire _0513_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2273" *)
  wire _0514_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2283" *)
  wire _0515_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2293" *)
  wire _0516_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2303" *)
  wire _0517_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2313" *)
  wire _0518_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2323" *)
  wire _0519_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2333" *)
  wire _0520_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2343" *)
  wire _0521_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2353" *)
  wire _0522_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2363" *)
  wire _0523_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2373" *)
  wire _0524_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2383" *)
  wire _0525_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2393" *)
  wire _0526_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2403" *)
  wire _0527_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2413" *)
  wire _0528_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2423" *)
  wire _0529_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2433" *)
  wire _0530_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2443" *)
  wire _0531_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2453" *)
  wire _0532_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2463" *)
  wire _0533_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2473" *)
  wire _0534_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2483" *)
  wire _0535_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2493" *)
  wire _0536_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2503" *)
  wire _0537_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2513" *)
  wire _0538_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2523" *)
  wire _0539_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2533" *)
  wire _0540_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2543" *)
  wire _0541_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2553" *)
  wire _0542_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2563" *)
  wire _0543_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2573" *)
  wire _0544_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2583" *)
  wire _0545_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2593" *)
  wire _0546_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2603" *)
  wire _0547_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2613" *)
  wire _0548_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2623" *)
  wire _0549_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2633" *)
  wire _0550_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2643" *)
  wire _0551_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2653" *)
  wire _0552_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2663" *)
  wire _0553_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2673" *)
  wire _0554_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2683" *)
  wire _0555_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2693" *)
  wire _0556_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2703" *)
  wire _0557_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2713" *)
  wire _0558_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2723" *)
  wire _0559_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2733" *)
  wire _0560_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2743" *)
  wire _0561_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2753" *)
  wire _0562_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2763" *)
  wire _0563_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2773" *)
  wire _0564_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2783" *)
  wire _0565_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2793" *)
  wire _0566_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2803" *)
  wire _0567_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2813" *)
  wire _0568_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2823" *)
  wire _0569_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2833" *)
  wire _0570_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2843" *)
  wire _0571_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2853" *)
  wire _0572_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2863" *)
  wire _0573_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2873" *)
  wire _0574_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2883" *)
  wire _0575_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2893" *)
  wire _0576_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2903" *)
  wire _0577_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2913" *)
  wire _0578_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2923" *)
  wire _0579_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2933" *)
  wire _0580_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2943" *)
  wire _0581_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2953" *)
  wire _0582_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2963" *)
  wire _0583_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2973" *)
  wire _0584_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2983" *)
  wire _0585_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2993" *)
  wire _0586_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3003" *)
  wire _0587_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3013" *)
  wire _0588_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3023" *)
  wire _0589_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3033" *)
  wire _0590_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3043" *)
  wire _0591_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3053" *)
  wire _0592_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3063" *)
  wire _0593_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3073" *)
  wire _0594_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3083" *)
  wire _0595_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3093" *)
  wire _0596_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3103" *)
  wire _0597_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3113" *)
  wire _0598_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3123" *)
  wire _0599_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3133" *)
  wire _0600_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3143" *)
  wire _0601_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3153" *)
  wire _0602_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3163" *)
  wire _0603_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3173" *)
  wire _0604_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3183" *)
  wire _0605_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3193" *)
  wire _0606_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3203" *)
  wire _0607_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3213" *)
  wire _0608_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3223" *)
  wire _0609_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3233" *)
  wire _0610_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3243" *)
  wire _0611_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3253" *)
  wire _0612_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3263" *)
  wire _0613_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3273" *)
  wire _0614_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3283" *)
  wire _0615_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3293" *)
  wire _0616_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3303" *)
  wire _0617_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3313" *)
  wire _0618_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3323" *)
  wire _0619_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3333" *)
  wire _0620_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3343" *)
  wire _0621_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3353" *)
  wire _0622_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3363" *)
  wire _0623_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3373" *)
  wire _0624_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3383" *)
  wire _0625_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3393" *)
  wire _0626_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3403" *)
  wire _0627_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3413" *)
  wire _0628_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3423" *)
  wire _0629_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3433" *)
  wire _0630_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3443" *)
  wire _0631_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3453" *)
  wire _0632_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3463" *)
  wire _0633_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3473" *)
  wire _0634_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3483" *)
  wire _0635_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3493" *)
  wire _0636_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3503" *)
  wire _0637_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3513" *)
  wire _0638_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3523" *)
  wire _0639_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3533" *)
  wire _0640_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3543" *)
  wire _0641_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3553" *)
  wire _0642_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3563" *)
  wire _0643_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3573" *)
  wire _0644_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3583" *)
  wire _0645_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3593" *)
  wire _0646_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3603" *)
  wire _0647_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3613" *)
  wire _0648_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3623" *)
  wire _0649_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3633" *)
  wire _0650_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3643" *)
  wire _0651_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3653" *)
  wire _0652_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3663" *)
  wire _0653_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3673" *)
  wire _0654_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3683" *)
  wire _0655_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3693" *)
  wire _0656_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3703" *)
  wire _0657_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3713" *)
  wire _0658_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3723" *)
  wire _0659_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3733" *)
  wire _0660_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3743" *)
  wire _0661_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3753" *)
  wire _0662_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3763" *)
  wire _0663_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3773" *)
  wire _0664_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3783" *)
  wire _0665_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3793" *)
  wire _0666_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3803" *)
  wire _0667_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3813" *)
  wire _0668_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3823" *)
  wire _0669_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3833" *)
  wire _0670_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3843" *)
  wire _0671_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3853" *)
  wire _0672_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3863" *)
  wire _0673_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3873" *)
  wire _0674_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3883" *)
  wire _0675_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4558" *)
  wire _0676_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4574" *)
  wire _0677_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4577" *)
  wire _0678_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4578" *)
  wire _0679_;
  wire _0680_;
  wire [15:0] _0681_;
  wire _0682_;
  wire _0683_;
  wire _0684_;
  wire _0685_;
  wire _0686_;
  wire _0687_;
  wire _0688_;
  wire _0689_;
  wire _0690_;
  wire _0691_;
  wire _0692_;
  wire _0693_;
  wire _0694_;
  wire _0695_;
  wire _0696_;
  wire _0697_;
  wire _0698_;
  wire _0699_;
  wire _0700_;
  wire _0701_;
  wire _0702_;
  wire _0703_;
  wire _0704_;
  wire _0705_;
  wire _0706_;
  wire _0707_;
  wire _0708_;
  wire _0709_;
  wire _0710_;
  wire _0711_;
  wire _0712_;
  wire _0713_;
  wire _0714_;
  wire _0715_;
  wire _0716_;
  wire _0717_;
  wire _0718_;
  wire _0719_;
  wire _0720_;
  wire _0721_;
  wire _0722_;
  wire _0723_;
  wire _0724_;
  wire _0725_;
  wire _0726_;
  wire _0727_;
  wire _0728_;
  wire _0729_;
  wire _0730_;
  wire _0731_;
  wire _0732_;
  wire _0733_;
  wire _0734_;
  wire _0735_;
  wire _0736_;
  wire _0737_;
  wire _0738_;
  wire _0739_;
  wire _0740_;
  wire _0741_;
  wire _0742_;
  wire _0743_;
  wire _0744_;
  wire _0745_;
  wire _0746_;
  wire _0747_;
  wire _0748_;
  wire _0749_;
  wire _0750_;
  wire _0751_;
  wire _0752_;
  wire _0753_;
  wire _0754_;
  wire _0755_;
  wire _0756_;
  wire _0757_;
  wire _0758_;
  wire _0759_;
  wire _0760_;
  wire _0761_;
  wire _0762_;
  wire _0763_;
  wire _0764_;
  wire _0765_;
  wire _0766_;
  wire _0767_;
  wire _0768_;
  wire _0769_;
  wire _0770_;
  wire _0771_;
  wire _0772_;
  wire _0773_;
  wire _0774_;
  wire _0775_;
  wire _0776_;
  wire _0777_;
  wire _0778_;
  wire _0779_;
  wire _0780_;
  wire _0781_;
  wire _0782_;
  wire _0783_;
  wire _0784_;
  wire _0785_;
  wire _0786_;
  wire _0787_;
  wire _0788_;
  wire _0789_;
  wire _0790_;
  wire _0791_;
  wire _0792_;
  wire _0793_;
  wire _0794_;
  wire _0795_;
  wire _0796_;
  wire _0797_;
  wire _0798_;
  wire _0799_;
  wire _0800_;
  wire _0801_;
  wire _0802_;
  wire _0803_;
  wire _0804_;
  wire _0805_;
  wire _0806_;
  wire _0807_;
  wire _0808_;
  wire _0809_;
  wire _0810_;
  wire _0811_;
  wire _0812_;
  wire _0813_;
  wire _0814_;
  wire _0815_;
  wire _0816_;
  wire _0817_;
  wire _0818_;
  wire _0819_;
  wire _0820_;
  wire _0821_;
  wire _0822_;
  wire _0823_;
  wire _0824_;
  wire _0825_;
  wire _0826_;
  wire _0827_;
  wire _0828_;
  wire _0829_;
  wire _0830_;
  wire _0831_;
  wire _0832_;
  wire _0833_;
  wire _0834_;
  wire _0835_;
  wire _0836_;
  wire _0837_;
  wire _0838_;
  wire _0839_;
  wire _0840_;
  wire _0841_;
  wire _0842_;
  wire _0843_;
  wire _0844_;
  wire _0845_;
  wire _0846_;
  wire _0847_;
  wire _0848_;
  wire _0849_;
  wire _0850_;
  wire _0851_;
  wire _0852_;
  wire _0853_;
  wire _0854_;
  wire _0855_;
  wire _0856_;
  wire _0857_;
  wire _0858_;
  wire _0859_;
  wire _0860_;
  wire _0861_;
  wire _0862_;
  wire _0863_;
  wire _0864_;
  wire _0865_;
  wire _0866_;
  wire _0867_;
  wire _0868_;
  wire _0869_;
  wire _0870_;
  wire _0871_;
  wire _0872_;
  wire _0873_;
  wire _0874_;
  wire _0875_;
  wire _0876_;
  wire _0877_;
  wire _0878_;
  wire _0879_;
  wire _0880_;
  wire _0881_;
  wire _0882_;
  wire _0883_;
  wire _0884_;
  wire _0885_;
  wire _0886_;
  wire _0887_;
  wire _0888_;
  wire _0889_;
  wire _0890_;
  wire _0891_;
  wire _0892_;
  wire _0893_;
  wire _0894_;
  wire _0895_;
  wire _0896_;
  wire _0897_;
  wire _0898_;
  wire _0899_;
  wire _0900_;
  wire _0901_;
  wire _0902_;
  wire _0903_;
  wire _0904_;
  wire _0905_;
  wire _0906_;
  wire _0907_;
  wire _0908_;
  wire _0909_;
  wire _0910_;
  wire _0911_;
  wire _0912_;
  wire _0913_;
  wire _0914_;
  wire _0915_;
  wire _0916_;
  wire _0917_;
  wire _0918_;
  wire _0919_;
  wire _0920_;
  wire _0921_;
  wire _0922_;
  wire _0923_;
  wire _0924_;
  wire _0925_;
  wire _0926_;
  wire _0927_;
  wire _0928_;
  wire _0929_;
  wire _0930_;
  wire _0931_;
  wire _0932_;
  wire _0933_;
  wire _0934_;
  wire _0935_;
  wire _0936_;
  wire _0937_;
  wire _0938_;
  wire [15:0] _0939_;
  wire [15:0] _0940_;
  wire [15:0] _0941_;
  wire [15:0] _0942_;
  wire [15:0] _0943_;
  wire [15:0] _0944_;
  wire _0945_;
  wire _0946_;
  wire _0947_;
  wire _0948_;
  wire _0949_;
  wire _0950_;
  wire _0951_;
  wire _0952_;
  wire _0953_;
  wire _0954_;
  wire _0955_;
  wire _0956_;
  wire _0957_;
  wire _0958_;
  wire _0959_;
  wire _0960_;
  wire _0961_;
  wire _0962_;
  wire _0963_;
  wire _0964_;
  wire _0965_;
  wire _0966_;
  wire _0967_;
  wire _0968_;
  wire _0969_;
  wire _0970_;
  wire _0971_;
  wire _0972_;
  wire _0973_;
  wire _0974_;
  wire _0975_;
  wire _0976_;
  wire _0977_;
  wire _0978_;
  wire _0979_;
  wire _0980_;
  wire _0981_;
  wire _0982_;
  wire _0983_;
  wire _0984_;
  wire _0985_;
  wire _0986_;
  wire _0987_;
  wire _0988_;
  wire _0989_;
  wire _0990_;
  wire _0991_;
  wire _0992_;
  wire _0993_;
  wire _0994_;
  wire _0995_;
  wire _0996_;
  wire _0997_;
  wire _0998_;
  wire _0999_;
  wire _1000_;
  wire _1001_;
  wire _1002_;
  wire _1003_;
  wire _1004_;
  wire _1005_;
  wire _1006_;
  wire _1007_;
  wire _1008_;
  wire _1009_;
  wire _1010_;
  wire _1011_;
  wire _1012_;
  wire _1013_;
  wire _1014_;
  wire _1015_;
  wire _1016_;
  wire _1017_;
  wire _1018_;
  wire _1019_;
  wire _1020_;
  wire _1021_;
  wire _1022_;
  wire _1023_;
  wire _1024_;
  wire _1025_;
  wire _1026_;
  wire _1027_;
  wire _1028_;
  wire _1029_;
  wire _1030_;
  wire _1031_;
  wire _1032_;
  wire _1033_;
  wire _1034_;
  wire _1035_;
  wire _1036_;
  wire _1037_;
  wire _1038_;
  wire _1039_;
  wire _1040_;
  wire _1041_;
  wire _1042_;
  wire _1043_;
  wire _1044_;
  wire _1045_;
  wire _1046_;
  wire _1047_;
  wire _1048_;
  wire _1049_;
  wire _1050_;
  wire _1051_;
  wire _1052_;
  wire _1053_;
  wire _1054_;
  wire _1055_;
  wire _1056_;
  wire _1057_;
  wire _1058_;
  wire _1059_;
  wire _1060_;
  wire _1061_;
  wire _1062_;
  wire _1063_;
  wire _1064_;
  wire _1065_;
  wire _1066_;
  wire _1067_;
  wire _1068_;
  wire _1069_;
  wire _1070_;
  wire _1071_;
  wire _1072_;
  wire _1073_;
  wire _1074_;
  wire _1075_;
  wire _1076_;
  wire _1077_;
  wire _1078_;
  wire _1079_;
  wire _1080_;
  wire _1081_;
  wire _1082_;
  wire _1083_;
  wire _1084_;
  wire _1085_;
  wire _1086_;
  wire _1087_;
  wire _1088_;
  wire _1089_;
  wire _1090_;
  wire _1091_;
  wire _1092_;
  wire _1093_;
  wire _1094_;
  wire _1095_;
  wire _1096_;
  wire _1097_;
  wire _1098_;
  wire _1099_;
  wire _1100_;
  wire _1101_;
  wire _1102_;
  wire _1103_;
  wire _1104_;
  wire _1105_;
  wire _1106_;
  wire _1107_;
  wire _1108_;
  wire _1109_;
  wire _1110_;
  wire _1111_;
  wire _1112_;
  wire _1113_;
  wire _1114_;
  wire _1115_;
  wire _1116_;
  wire _1117_;
  wire _1118_;
  wire _1119_;
  wire _1120_;
  wire _1121_;
  wire _1122_;
  wire _1123_;
  wire _1124_;
  wire _1125_;
  wire _1126_;
  wire _1127_;
  wire _1128_;
  wire _1129_;
  wire _1130_;
  wire _1131_;
  wire _1132_;
  wire _1133_;
  wire _1134_;
  wire _1135_;
  wire _1136_;
  wire _1137_;
  wire _1138_;
  wire _1139_;
  wire _1140_;
  wire _1141_;
  wire _1142_;
  wire _1143_;
  wire _1144_;
  wire _1145_;
  wire _1146_;
  wire _1147_;
  wire _1148_;
  wire _1149_;
  wire _1150_;
  wire _1151_;
  wire _1152_;
  wire _1153_;
  wire _1154_;
  wire _1155_;
  wire _1156_;
  wire _1157_;
  wire _1158_;
  wire _1159_;
  wire _1160_;
  wire _1161_;
  wire _1162_;
  wire _1163_;
  wire _1164_;
  wire _1165_;
  wire _1166_;
  wire _1167_;
  wire _1168_;
  wire _1169_;
  wire _1170_;
  wire _1171_;
  wire _1172_;
  wire _1173_;
  wire _1174_;
  wire _1175_;
  wire _1176_;
  wire _1177_;
  wire _1178_;
  wire _1179_;
  wire _1180_;
  wire _1181_;
  wire _1182_;
  wire _1183_;
  wire _1184_;
  wire _1185_;
  wire _1186_;
  wire _1187_;
  wire _1188_;
  wire _1189_;
  wire _1190_;
  wire _1191_;
  wire _1192_;
  wire _1193_;
  wire _1194_;
  wire _1195_;
  wire _1196_;
  wire _1197_;
  wire _1198_;
  wire _1199_;
  wire _1200_;
  wire _1201_;
  wire [15:0] _1202_;
  wire [15:0] _1203_;
  wire [15:0] _1204_;
  wire [15:0] _1205_;
  wire [15:0] _1206_;
  wire [15:0] _1207_;
  wire _1208_;
  wire _1209_;
  wire _1210_;
  wire _1211_;
  wire _1212_;
  wire _1213_;
  wire _1214_;
  wire _1215_;
  wire _1216_;
  wire _1217_;
  wire _1218_;
  wire _1219_;
  wire _1220_;
  wire _1221_;
  wire _1222_;
  wire _1223_;
  wire _1224_;
  wire _1225_;
  wire _1226_;
  wire _1227_;
  wire _1228_;
  wire _1229_;
  wire _1230_;
  wire _1231_;
  wire _1232_;
  wire _1233_;
  wire _1234_;
  wire _1235_;
  wire _1236_;
  wire _1237_;
  wire _1238_;
  wire _1239_;
  wire _1240_;
  wire _1241_;
  wire _1242_;
  wire _1243_;
  wire _1244_;
  wire _1245_;
  wire _1246_;
  wire _1247_;
  wire _1248_;
  wire _1249_;
  wire _1250_;
  wire _1251_;
  wire _1252_;
  wire _1253_;
  wire _1254_;
  wire _1255_;
  wire _1256_;
  wire _1257_;
  wire _1258_;
  wire _1259_;
  wire _1260_;
  wire _1261_;
  wire _1262_;
  wire _1263_;
  wire _1264_;
  wire _1265_;
  wire _1266_;
  wire _1267_;
  wire _1268_;
  wire _1269_;
  wire _1270_;
  wire _1271_;
  wire _1272_;
  wire _1273_;
  wire _1274_;
  wire _1275_;
  wire _1276_;
  wire _1277_;
  wire _1278_;
  wire _1279_;
  wire _1280_;
  wire _1281_;
  wire _1282_;
  wire _1283_;
  wire _1284_;
  wire _1285_;
  wire _1286_;
  wire _1287_;
  wire _1288_;
  wire _1289_;
  wire _1290_;
  wire _1291_;
  wire _1292_;
  wire _1293_;
  wire _1294_;
  wire _1295_;
  wire _1296_;
  wire _1297_;
  wire _1298_;
  wire _1299_;
  wire _1300_;
  wire _1301_;
  wire _1302_;
  wire _1303_;
  wire _1304_;
  wire _1305_;
  wire _1306_;
  wire _1307_;
  wire _1308_;
  wire _1309_;
  wire _1310_;
  wire _1311_;
  wire _1312_;
  wire _1313_;
  wire _1314_;
  wire _1315_;
  wire _1316_;
  wire _1317_;
  wire _1318_;
  wire _1319_;
  wire _1320_;
  wire _1321_;
  wire _1322_;
  wire _1323_;
  wire _1324_;
  wire _1325_;
  wire _1326_;
  wire _1327_;
  wire _1328_;
  wire _1329_;
  wire _1330_;
  wire _1331_;
  wire _1332_;
  wire _1333_;
  wire _1334_;
  wire _1335_;
  wire _1336_;
  wire _1337_;
  wire _1338_;
  wire _1339_;
  wire _1340_;
  wire _1341_;
  wire _1342_;
  wire _1343_;
  wire _1344_;
  wire _1345_;
  wire _1346_;
  wire _1347_;
  wire _1348_;
  wire _1349_;
  wire _1350_;
  wire _1351_;
  wire _1352_;
  wire _1353_;
  wire _1354_;
  wire _1355_;
  wire _1356_;
  wire _1357_;
  wire _1358_;
  wire _1359_;
  wire _1360_;
  wire _1361_;
  wire _1362_;
  wire _1363_;
  wire _1364_;
  wire _1365_;
  wire _1366_;
  wire _1367_;
  wire _1368_;
  wire _1369_;
  wire _1370_;
  wire _1371_;
  wire _1372_;
  wire _1373_;
  wire _1374_;
  wire _1375_;
  wire _1376_;
  wire _1377_;
  wire _1378_;
  wire _1379_;
  wire _1380_;
  wire _1381_;
  wire _1382_;
  wire _1383_;
  wire _1384_;
  wire _1385_;
  wire _1386_;
  wire _1387_;
  wire _1388_;
  wire _1389_;
  wire _1390_;
  wire _1391_;
  wire _1392_;
  wire _1393_;
  wire _1394_;
  wire _1395_;
  wire _1396_;
  wire _1397_;
  wire _1398_;
  wire _1399_;
  wire _1400_;
  wire _1401_;
  wire _1402_;
  wire _1403_;
  wire _1404_;
  wire _1405_;
  wire _1406_;
  wire _1407_;
  wire _1408_;
  wire _1409_;
  wire _1410_;
  wire _1411_;
  wire _1412_;
  wire _1413_;
  wire _1414_;
  wire _1415_;
  wire _1416_;
  wire _1417_;
  wire _1418_;
  wire _1419_;
  wire _1420_;
  wire _1421_;
  wire _1422_;
  wire _1423_;
  wire _1424_;
  wire _1425_;
  wire _1426_;
  wire _1427_;
  wire _1428_;
  wire _1429_;
  wire _1430_;
  wire _1431_;
  wire _1432_;
  wire _1433_;
  wire _1434_;
  wire _1435_;
  wire _1436_;
  wire _1437_;
  wire _1438_;
  wire _1439_;
  wire _1440_;
  wire _1441_;
  wire _1442_;
  wire _1443_;
  wire _1444_;
  wire _1445_;
  wire _1446_;
  wire _1447_;
  wire _1448_;
  wire _1449_;
  wire _1450_;
  wire _1451_;
  wire _1452_;
  wire _1453_;
  wire _1454_;
  wire _1455_;
  wire _1456_;
  wire _1457_;
  wire _1458_;
  wire _1459_;
  wire _1460_;
  wire _1461_;
  wire _1462_;
  wire _1463_;
  wire _1464_;
  wire [15:0] _1465_;
  wire [15:0] _1466_;
  wire [15:0] _1467_;
  wire [15:0] _1468_;
  wire [15:0] _1469_;
  wire [15:0] _1470_;
  wire _1471_;
  wire _1472_;
  wire _1473_;
  wire _1474_;
  wire _1475_;
  wire _1476_;
  wire _1477_;
  wire _1478_;
  wire _1479_;
  wire _1480_;
  wire _1481_;
  wire _1482_;
  wire _1483_;
  wire _1484_;
  wire _1485_;
  wire _1486_;
  wire _1487_;
  wire _1488_;
  wire _1489_;
  wire _1490_;
  wire _1491_;
  wire _1492_;
  wire _1493_;
  wire _1494_;
  wire _1495_;
  wire _1496_;
  wire _1497_;
  wire _1498_;
  wire _1499_;
  wire _1500_;
  wire _1501_;
  wire _1502_;
  wire _1503_;
  wire _1504_;
  wire _1505_;
  wire _1506_;
  wire _1507_;
  wire _1508_;
  wire _1509_;
  wire _1510_;
  wire _1511_;
  wire _1512_;
  wire _1513_;
  wire _1514_;
  wire _1515_;
  wire _1516_;
  wire _1517_;
  wire _1518_;
  wire _1519_;
  wire _1520_;
  wire _1521_;
  wire _1522_;
  wire _1523_;
  wire _1524_;
  wire _1525_;
  wire _1526_;
  wire _1527_;
  wire _1528_;
  wire _1529_;
  wire _1530_;
  wire _1531_;
  wire _1532_;
  wire _1533_;
  wire _1534_;
  wire _1535_;
  wire _1536_;
  wire _1537_;
  wire _1538_;
  wire _1539_;
  wire _1540_;
  wire _1541_;
  wire _1542_;
  wire _1543_;
  wire _1544_;
  wire _1545_;
  wire _1546_;
  wire _1547_;
  wire _1548_;
  wire _1549_;
  wire _1550_;
  wire _1551_;
  wire _1552_;
  wire _1553_;
  wire _1554_;
  wire _1555_;
  wire _1556_;
  wire _1557_;
  wire _1558_;
  wire _1559_;
  wire _1560_;
  wire _1561_;
  wire _1562_;
  wire _1563_;
  wire _1564_;
  wire _1565_;
  wire _1566_;
  wire _1567_;
  wire _1568_;
  wire _1569_;
  wire _1570_;
  wire _1571_;
  wire _1572_;
  wire _1573_;
  wire _1574_;
  wire _1575_;
  wire _1576_;
  wire _1577_;
  wire _1578_;
  wire _1579_;
  wire _1580_;
  wire _1581_;
  wire _1582_;
  wire _1583_;
  wire _1584_;
  wire _1585_;
  wire _1586_;
  wire _1587_;
  wire _1588_;
  wire _1589_;
  wire _1590_;
  wire _1591_;
  wire _1592_;
  wire _1593_;
  wire _1594_;
  wire _1595_;
  wire _1596_;
  wire _1597_;
  wire _1598_;
  wire _1599_;
  wire _1600_;
  wire _1601_;
  wire _1602_;
  wire _1603_;
  wire _1604_;
  wire _1605_;
  wire _1606_;
  wire _1607_;
  wire _1608_;
  wire _1609_;
  wire _1610_;
  wire _1611_;
  wire _1612_;
  wire _1613_;
  wire _1614_;
  wire _1615_;
  wire _1616_;
  wire _1617_;
  wire _1618_;
  wire _1619_;
  wire _1620_;
  wire _1621_;
  wire _1622_;
  wire _1623_;
  wire _1624_;
  wire _1625_;
  wire _1626_;
  wire _1627_;
  wire _1628_;
  wire _1629_;
  wire _1630_;
  wire _1631_;
  wire _1632_;
  wire _1633_;
  wire _1634_;
  wire _1635_;
  wire _1636_;
  wire _1637_;
  wire _1638_;
  wire _1639_;
  wire _1640_;
  wire _1641_;
  wire _1642_;
  wire _1643_;
  wire _1644_;
  wire _1645_;
  wire _1646_;
  wire _1647_;
  wire _1648_;
  wire _1649_;
  wire _1650_;
  wire _1651_;
  wire _1652_;
  wire _1653_;
  wire _1654_;
  wire _1655_;
  wire _1656_;
  wire _1657_;
  wire _1658_;
  wire _1659_;
  wire _1660_;
  wire _1661_;
  wire _1662_;
  wire _1663_;
  wire _1664_;
  wire _1665_;
  wire _1666_;
  wire _1667_;
  wire _1668_;
  wire _1669_;
  wire _1670_;
  wire _1671_;
  wire _1672_;
  wire _1673_;
  wire _1674_;
  wire _1675_;
  wire _1676_;
  wire _1677_;
  wire _1678_;
  wire _1679_;
  wire _1680_;
  wire _1681_;
  wire _1682_;
  wire _1683_;
  wire _1684_;
  wire _1685_;
  wire _1686_;
  wire _1687_;
  wire _1688_;
  wire _1689_;
  wire _1690_;
  wire _1691_;
  wire _1692_;
  wire _1693_;
  wire _1694_;
  wire _1695_;
  wire _1696_;
  wire _1697_;
  wire _1698_;
  wire _1699_;
  wire _1700_;
  wire _1701_;
  wire _1702_;
  wire _1703_;
  wire _1704_;
  wire _1705_;
  wire _1706_;
  wire _1707_;
  wire _1708_;
  wire _1709_;
  wire _1710_;
  wire _1711_;
  wire _1712_;
  wire _1713_;
  wire _1714_;
  wire _1715_;
  wire _1716_;
  wire _1717_;
  wire _1718_;
  wire _1719_;
  wire _1720_;
  wire _1721_;
  wire _1722_;
  wire _1723_;
  wire _1724_;
  wire _1725_;
  wire _1726_;
  wire _1727_;
  wire [15:0] _1728_;
  wire [15:0] _1729_;
  wire [15:0] _1730_;
  wire [15:0] _1731_;
  wire [15:0] _1732_;
  wire [15:0] _1733_;
  wire _1734_;
  wire _1735_;
  wire _1736_;
  wire _1737_;
  wire _1738_;
  wire _1739_;
  wire _1740_;
  wire _1741_;
  wire _1742_;
  wire _1743_;
  wire _1744_;
  wire _1745_;
  wire _1746_;
  wire _1747_;
  wire _1748_;
  wire _1749_;
  wire _1750_;
  wire _1751_;
  wire _1752_;
  wire _1753_;
  wire _1754_;
  wire _1755_;
  wire _1756_;
  wire _1757_;
  wire _1758_;
  wire _1759_;
  wire _1760_;
  wire _1761_;
  wire _1762_;
  wire _1763_;
  wire _1764_;
  wire _1765_;
  wire _1766_;
  wire _1767_;
  wire _1768_;
  wire _1769_;
  wire _1770_;
  wire _1771_;
  wire _1772_;
  wire _1773_;
  wire _1774_;
  wire _1775_;
  wire _1776_;
  wire _1777_;
  wire _1778_;
  wire _1779_;
  wire _1780_;
  wire _1781_;
  wire _1782_;
  wire _1783_;
  wire _1784_;
  wire _1785_;
  wire _1786_;
  wire _1787_;
  wire _1788_;
  wire _1789_;
  wire _1790_;
  wire _1791_;
  wire _1792_;
  wire _1793_;
  wire _1794_;
  wire _1795_;
  wire _1796_;
  wire _1797_;
  wire _1798_;
  wire _1799_;
  wire _1800_;
  wire _1801_;
  wire _1802_;
  wire _1803_;
  wire _1804_;
  wire _1805_;
  wire _1806_;
  wire _1807_;
  wire _1808_;
  wire _1809_;
  wire _1810_;
  wire _1811_;
  wire _1812_;
  wire _1813_;
  wire _1814_;
  wire _1815_;
  wire _1816_;
  wire _1817_;
  wire _1818_;
  wire _1819_;
  wire _1820_;
  wire _1821_;
  wire _1822_;
  wire _1823_;
  wire _1824_;
  wire _1825_;
  wire _1826_;
  wire _1827_;
  wire _1828_;
  wire _1829_;
  wire _1830_;
  wire _1831_;
  wire _1832_;
  wire _1833_;
  wire _1834_;
  wire _1835_;
  wire _1836_;
  wire _1837_;
  wire _1838_;
  wire _1839_;
  wire _1840_;
  wire _1841_;
  wire _1842_;
  wire _1843_;
  wire _1844_;
  wire _1845_;
  wire _1846_;
  wire _1847_;
  wire _1848_;
  wire _1849_;
  wire _1850_;
  wire _1851_;
  wire _1852_;
  wire _1853_;
  wire _1854_;
  wire _1855_;
  wire _1856_;
  wire _1857_;
  wire _1858_;
  wire _1859_;
  wire _1860_;
  wire _1861_;
  wire _1862_;
  wire _1863_;
  wire _1864_;
  wire _1865_;
  wire _1866_;
  wire _1867_;
  wire _1868_;
  wire _1869_;
  wire _1870_;
  wire _1871_;
  wire _1872_;
  wire _1873_;
  wire _1874_;
  wire _1875_;
  wire _1876_;
  wire _1877_;
  wire _1878_;
  wire _1879_;
  wire _1880_;
  wire _1881_;
  wire _1882_;
  wire _1883_;
  wire _1884_;
  wire _1885_;
  wire _1886_;
  wire _1887_;
  wire _1888_;
  wire _1889_;
  wire _1890_;
  wire _1891_;
  wire _1892_;
  wire _1893_;
  wire _1894_;
  wire _1895_;
  wire _1896_;
  wire _1897_;
  wire _1898_;
  wire _1899_;
  wire _1900_;
  wire _1901_;
  wire _1902_;
  wire _1903_;
  wire _1904_;
  wire _1905_;
  wire _1906_;
  wire _1907_;
  wire _1908_;
  wire _1909_;
  wire _1910_;
  wire _1911_;
  wire _1912_;
  wire _1913_;
  wire _1914_;
  wire _1915_;
  wire _1916_;
  wire _1917_;
  wire _1918_;
  wire _1919_;
  wire _1920_;
  wire _1921_;
  wire _1922_;
  wire _1923_;
  wire _1924_;
  wire _1925_;
  wire _1926_;
  wire _1927_;
  wire _1928_;
  wire _1929_;
  wire _1930_;
  wire _1931_;
  wire _1932_;
  wire _1933_;
  wire _1934_;
  wire _1935_;
  wire _1936_;
  wire _1937_;
  wire _1938_;
  wire _1939_;
  wire _1940_;
  wire _1941_;
  wire _1942_;
  wire _1943_;
  wire _1944_;
  wire _1945_;
  wire _1946_;
  wire _1947_;
  wire _1948_;
  wire _1949_;
  wire _1950_;
  wire _1951_;
  wire _1952_;
  wire _1953_;
  wire _1954_;
  wire _1955_;
  wire _1956_;
  wire _1957_;
  wire _1958_;
  wire _1959_;
  wire _1960_;
  wire _1961_;
  wire _1962_;
  wire _1963_;
  wire _1964_;
  wire _1965_;
  wire _1966_;
  wire _1967_;
  wire _1968_;
  wire _1969_;
  wire _1970_;
  wire _1971_;
  wire _1972_;
  wire _1973_;
  wire _1974_;
  wire _1975_;
  wire _1976_;
  wire _1977_;
  wire _1978_;
  wire _1979_;
  wire _1980_;
  wire _1981_;
  wire _1982_;
  wire _1983_;
  wire _1984_;
  wire _1985_;
  wire _1986_;
  wire _1987_;
  wire _1988_;
  wire _1989_;
  wire _1990_;
  wire [15:0] _1991_;
  wire [15:0] _1992_;
  wire [15:0] _1993_;
  wire [15:0] _1994_;
  wire [15:0] _1995_;
  wire [15:0] _1996_;
  wire _1997_;
  wire _1998_;
  wire _1999_;
  wire _2000_;
  wire _2001_;
  wire _2002_;
  wire _2003_;
  wire _2004_;
  wire _2005_;
  wire _2006_;
  wire _2007_;
  wire _2008_;
  wire _2009_;
  wire _2010_;
  wire _2011_;
  wire _2012_;
  wire _2013_;
  wire _2014_;
  wire _2015_;
  wire _2016_;
  wire _2017_;
  wire _2018_;
  wire _2019_;
  wire _2020_;
  wire _2021_;
  wire _2022_;
  wire _2023_;
  wire _2024_;
  wire _2025_;
  wire _2026_;
  wire _2027_;
  wire _2028_;
  wire _2029_;
  wire _2030_;
  wire _2031_;
  wire _2032_;
  wire _2033_;
  wire _2034_;
  wire _2035_;
  wire _2036_;
  wire _2037_;
  wire _2038_;
  wire _2039_;
  wire _2040_;
  wire _2041_;
  wire _2042_;
  wire _2043_;
  wire _2044_;
  wire _2045_;
  wire _2046_;
  wire _2047_;
  wire _2048_;
  wire _2049_;
  wire _2050_;
  wire _2051_;
  wire _2052_;
  wire _2053_;
  wire _2054_;
  wire _2055_;
  wire _2056_;
  wire _2057_;
  wire _2058_;
  wire _2059_;
  wire _2060_;
  wire _2061_;
  wire _2062_;
  wire _2063_;
  wire _2064_;
  wire _2065_;
  wire _2066_;
  wire _2067_;
  wire _2068_;
  wire _2069_;
  wire _2070_;
  wire _2071_;
  wire _2072_;
  wire _2073_;
  wire _2074_;
  wire _2075_;
  wire _2076_;
  wire _2077_;
  wire _2078_;
  wire _2079_;
  wire _2080_;
  wire _2081_;
  wire _2082_;
  wire _2083_;
  wire _2084_;
  wire _2085_;
  wire _2086_;
  wire _2087_;
  wire _2088_;
  wire _2089_;
  wire _2090_;
  wire _2091_;
  wire _2092_;
  wire _2093_;
  wire _2094_;
  wire _2095_;
  wire _2096_;
  wire _2097_;
  wire _2098_;
  wire _2099_;
  wire _2100_;
  wire _2101_;
  wire _2102_;
  wire _2103_;
  wire _2104_;
  wire _2105_;
  wire _2106_;
  wire _2107_;
  wire _2108_;
  wire _2109_;
  wire _2110_;
  wire _2111_;
  wire _2112_;
  wire _2113_;
  wire _2114_;
  wire _2115_;
  wire _2116_;
  wire _2117_;
  wire _2118_;
  wire _2119_;
  wire _2120_;
  wire _2121_;
  wire _2122_;
  wire _2123_;
  wire _2124_;
  wire _2125_;
  wire _2126_;
  wire _2127_;
  wire _2128_;
  wire _2129_;
  wire _2130_;
  wire _2131_;
  wire _2132_;
  wire _2133_;
  wire _2134_;
  wire _2135_;
  wire _2136_;
  wire _2137_;
  wire _2138_;
  wire _2139_;
  wire _2140_;
  wire _2141_;
  wire _2142_;
  wire _2143_;
  wire _2144_;
  wire _2145_;
  wire _2146_;
  wire _2147_;
  wire _2148_;
  wire _2149_;
  wire _2150_;
  wire _2151_;
  wire _2152_;
  wire _2153_;
  wire _2154_;
  wire _2155_;
  wire _2156_;
  wire _2157_;
  wire _2158_;
  wire _2159_;
  wire _2160_;
  wire _2161_;
  wire _2162_;
  wire _2163_;
  wire _2164_;
  wire _2165_;
  wire _2166_;
  wire _2167_;
  wire _2168_;
  wire _2169_;
  wire _2170_;
  wire _2171_;
  wire _2172_;
  wire _2173_;
  wire _2174_;
  wire _2175_;
  wire _2176_;
  wire _2177_;
  wire _2178_;
  wire _2179_;
  wire _2180_;
  wire _2181_;
  wire _2182_;
  wire _2183_;
  wire _2184_;
  wire _2185_;
  wire _2186_;
  wire _2187_;
  wire _2188_;
  wire _2189_;
  wire _2190_;
  wire _2191_;
  wire _2192_;
  wire _2193_;
  wire _2194_;
  wire _2195_;
  wire _2196_;
  wire _2197_;
  wire _2198_;
  wire _2199_;
  wire _2200_;
  wire _2201_;
  wire _2202_;
  wire _2203_;
  wire _2204_;
  wire _2205_;
  wire _2206_;
  wire _2207_;
  wire _2208_;
  wire _2209_;
  wire _2210_;
  wire _2211_;
  wire _2212_;
  wire _2213_;
  wire _2214_;
  wire _2215_;
  wire _2216_;
  wire _2217_;
  wire _2218_;
  wire _2219_;
  wire _2220_;
  wire _2221_;
  wire _2222_;
  wire _2223_;
  wire _2224_;
  wire _2225_;
  wire _2226_;
  wire _2227_;
  wire _2228_;
  wire _2229_;
  wire _2230_;
  wire _2231_;
  wire _2232_;
  wire _2233_;
  wire _2234_;
  wire _2235_;
  wire _2236_;
  wire _2237_;
  wire _2238_;
  wire _2239_;
  wire _2240_;
  wire _2241_;
  wire _2242_;
  wire _2243_;
  wire _2244_;
  wire _2245_;
  wire _2246_;
  wire _2247_;
  wire _2248_;
  wire _2249_;
  wire _2250_;
  wire _2251_;
  wire _2252_;
  wire _2253_;
  wire [15:0] _2254_;
  wire [15:0] _2255_;
  wire [15:0] _2256_;
  wire [15:0] _2257_;
  wire [15:0] _2258_;
  wire [15:0] _2259_;
  wire _2260_;
  wire _2261_;
  wire _2262_;
  wire _2263_;
  wire _2264_;
  wire _2265_;
  wire _2266_;
  wire _2267_;
  wire _2268_;
  wire _2269_;
  wire _2270_;
  wire _2271_;
  wire _2272_;
  wire _2273_;
  wire _2274_;
  wire _2275_;
  wire _2276_;
  wire _2277_;
  wire _2278_;
  wire _2279_;
  wire _2280_;
  wire _2281_;
  wire _2282_;
  wire _2283_;
  wire _2284_;
  wire _2285_;
  wire _2286_;
  wire _2287_;
  wire _2288_;
  wire _2289_;
  wire _2290_;
  wire _2291_;
  wire _2292_;
  wire _2293_;
  wire _2294_;
  wire _2295_;
  wire _2296_;
  wire _2297_;
  wire _2298_;
  wire _2299_;
  wire _2300_;
  wire _2301_;
  wire _2302_;
  wire _2303_;
  wire _2304_;
  wire _2305_;
  wire _2306_;
  wire _2307_;
  wire _2308_;
  wire _2309_;
  wire _2310_;
  wire _2311_;
  wire _2312_;
  wire _2313_;
  wire _2314_;
  wire _2315_;
  wire _2316_;
  wire _2317_;
  wire _2318_;
  wire _2319_;
  wire _2320_;
  wire _2321_;
  wire _2322_;
  wire _2323_;
  wire _2324_;
  wire _2325_;
  wire _2326_;
  wire _2327_;
  wire _2328_;
  wire _2329_;
  wire _2330_;
  wire _2331_;
  wire _2332_;
  wire _2333_;
  wire _2334_;
  wire _2335_;
  wire _2336_;
  wire _2337_;
  wire _2338_;
  wire _2339_;
  wire _2340_;
  wire _2341_;
  wire _2342_;
  wire _2343_;
  wire _2344_;
  wire _2345_;
  wire _2346_;
  wire _2347_;
  wire _2348_;
  wire _2349_;
  wire _2350_;
  wire _2351_;
  wire _2352_;
  wire _2353_;
  wire _2354_;
  wire _2355_;
  wire _2356_;
  wire _2357_;
  wire _2358_;
  wire _2359_;
  wire _2360_;
  wire _2361_;
  wire _2362_;
  wire _2363_;
  wire _2364_;
  wire _2365_;
  wire _2366_;
  wire _2367_;
  wire _2368_;
  wire _2369_;
  wire _2370_;
  wire _2371_;
  wire _2372_;
  wire _2373_;
  wire _2374_;
  wire _2375_;
  wire _2376_;
  wire _2377_;
  wire _2378_;
  wire _2379_;
  wire _2380_;
  wire _2381_;
  wire _2382_;
  wire _2383_;
  wire _2384_;
  wire _2385_;
  wire _2386_;
  wire _2387_;
  wire _2388_;
  wire _2389_;
  wire _2390_;
  wire _2391_;
  wire _2392_;
  wire _2393_;
  wire _2394_;
  wire _2395_;
  wire _2396_;
  wire _2397_;
  wire _2398_;
  wire _2399_;
  wire _2400_;
  wire _2401_;
  wire _2402_;
  wire _2403_;
  wire _2404_;
  wire _2405_;
  wire _2406_;
  wire _2407_;
  wire _2408_;
  wire _2409_;
  wire _2410_;
  wire _2411_;
  wire _2412_;
  wire _2413_;
  wire _2414_;
  wire _2415_;
  wire _2416_;
  wire _2417_;
  wire _2418_;
  wire _2419_;
  wire _2420_;
  wire _2421_;
  wire _2422_;
  wire _2423_;
  wire _2424_;
  wire _2425_;
  wire _2426_;
  wire _2427_;
  wire _2428_;
  wire _2429_;
  wire _2430_;
  wire _2431_;
  wire _2432_;
  wire _2433_;
  wire _2434_;
  wire _2435_;
  wire _2436_;
  wire _2437_;
  wire _2438_;
  wire _2439_;
  wire _2440_;
  wire _2441_;
  wire _2442_;
  wire _2443_;
  wire _2444_;
  wire _2445_;
  wire _2446_;
  wire _2447_;
  wire _2448_;
  wire _2449_;
  wire _2450_;
  wire _2451_;
  wire _2452_;
  wire _2453_;
  wire _2454_;
  wire _2455_;
  wire _2456_;
  wire _2457_;
  wire _2458_;
  wire _2459_;
  wire _2460_;
  wire _2461_;
  wire _2462_;
  wire _2463_;
  wire _2464_;
  wire _2465_;
  wire _2466_;
  wire _2467_;
  wire _2468_;
  wire _2469_;
  wire _2470_;
  wire _2471_;
  wire _2472_;
  wire _2473_;
  wire _2474_;
  wire _2475_;
  wire _2476_;
  wire _2477_;
  wire _2478_;
  wire _2479_;
  wire _2480_;
  wire _2481_;
  wire _2482_;
  wire _2483_;
  wire _2484_;
  wire _2485_;
  wire _2486_;
  wire _2487_;
  wire _2488_;
  wire _2489_;
  wire _2490_;
  wire _2491_;
  wire _2492_;
  wire _2493_;
  wire _2494_;
  wire _2495_;
  wire _2496_;
  wire _2497_;
  wire _2498_;
  wire _2499_;
  wire _2500_;
  wire _2501_;
  wire _2502_;
  wire _2503_;
  wire _2504_;
  wire _2505_;
  wire _2506_;
  wire _2507_;
  wire _2508_;
  wire _2509_;
  wire _2510_;
  wire _2511_;
  wire _2512_;
  wire _2513_;
  wire _2514_;
  wire _2515_;
  wire _2516_;
  wire [15:0] _2517_;
  wire [15:0] _2518_;
  wire [15:0] _2519_;
  wire [15:0] _2520_;
  wire [15:0] _2521_;
  wire [15:0] _2522_;
  wire _2523_;
  wire _2524_;
  wire _2525_;
  wire _2526_;
  wire _2527_;
  wire _2528_;
  wire _2529_;
  wire _2530_;
  wire _2531_;
  wire _2532_;
  wire _2533_;
  wire _2534_;
  wire _2535_;
  wire _2536_;
  wire _2537_;
  wire _2538_;
  wire _2539_;
  wire _2540_;
  wire _2541_;
  wire _2542_;
  wire _2543_;
  wire _2544_;
  wire _2545_;
  wire _2546_;
  wire _2547_;
  wire _2548_;
  wire _2549_;
  wire _2550_;
  wire _2551_;
  wire _2552_;
  wire _2553_;
  wire _2554_;
  wire _2555_;
  wire _2556_;
  wire _2557_;
  wire _2558_;
  wire _2559_;
  wire _2560_;
  wire _2561_;
  wire _2562_;
  wire _2563_;
  wire _2564_;
  wire _2565_;
  wire _2566_;
  wire _2567_;
  wire _2568_;
  wire _2569_;
  wire _2570_;
  wire _2571_;
  wire _2572_;
  wire _2573_;
  wire _2574_;
  wire _2575_;
  wire _2576_;
  wire _2577_;
  wire _2578_;
  wire _2579_;
  wire _2580_;
  wire _2581_;
  wire _2582_;
  wire _2583_;
  wire _2584_;
  wire _2585_;
  wire _2586_;
  wire _2587_;
  wire _2588_;
  wire _2589_;
  wire _2590_;
  wire _2591_;
  wire _2592_;
  wire _2593_;
  wire _2594_;
  wire _2595_;
  wire _2596_;
  wire _2597_;
  wire _2598_;
  wire _2599_;
  wire _2600_;
  wire _2601_;
  wire _2602_;
  wire _2603_;
  wire _2604_;
  wire _2605_;
  wire _2606_;
  wire _2607_;
  wire _2608_;
  wire _2609_;
  wire _2610_;
  wire _2611_;
  wire _2612_;
  wire _2613_;
  wire _2614_;
  wire _2615_;
  wire _2616_;
  wire _2617_;
  wire _2618_;
  wire _2619_;
  wire _2620_;
  wire _2621_;
  wire _2622_;
  wire _2623_;
  wire _2624_;
  wire _2625_;
  wire _2626_;
  wire _2627_;
  wire _2628_;
  wire _2629_;
  wire _2630_;
  wire _2631_;
  wire _2632_;
  wire _2633_;
  wire _2634_;
  wire _2635_;
  wire _2636_;
  wire _2637_;
  wire _2638_;
  wire _2639_;
  wire _2640_;
  wire _2641_;
  wire _2642_;
  wire _2643_;
  wire _2644_;
  wire _2645_;
  wire _2646_;
  wire _2647_;
  wire _2648_;
  wire _2649_;
  wire _2650_;
  wire _2651_;
  wire _2652_;
  wire _2653_;
  wire _2654_;
  wire _2655_;
  wire _2656_;
  wire _2657_;
  wire _2658_;
  wire _2659_;
  wire _2660_;
  wire _2661_;
  wire _2662_;
  wire _2663_;
  wire _2664_;
  wire _2665_;
  wire _2666_;
  wire _2667_;
  wire _2668_;
  wire _2669_;
  wire _2670_;
  wire _2671_;
  wire _2672_;
  wire _2673_;
  wire _2674_;
  wire _2675_;
  wire _2676_;
  wire _2677_;
  wire _2678_;
  wire _2679_;
  wire _2680_;
  wire _2681_;
  wire _2682_;
  wire _2683_;
  wire _2684_;
  wire _2685_;
  wire _2686_;
  wire _2687_;
  wire _2688_;
  wire _2689_;
  wire _2690_;
  wire _2691_;
  wire _2692_;
  wire _2693_;
  wire _2694_;
  wire _2695_;
  wire _2696_;
  wire _2697_;
  wire _2698_;
  wire _2699_;
  wire _2700_;
  wire _2701_;
  wire _2702_;
  wire _2703_;
  wire _2704_;
  wire _2705_;
  wire _2706_;
  wire _2707_;
  wire _2708_;
  wire _2709_;
  wire _2710_;
  wire _2711_;
  wire _2712_;
  wire _2713_;
  wire _2714_;
  wire _2715_;
  wire _2716_;
  wire _2717_;
  wire _2718_;
  wire _2719_;
  wire _2720_;
  wire _2721_;
  wire _2722_;
  wire _2723_;
  wire _2724_;
  wire _2725_;
  wire _2726_;
  wire _2727_;
  wire _2728_;
  wire _2729_;
  wire _2730_;
  wire _2731_;
  wire _2732_;
  wire _2733_;
  wire _2734_;
  wire _2735_;
  wire _2736_;
  wire _2737_;
  wire _2738_;
  wire _2739_;
  wire _2740_;
  wire _2741_;
  wire _2742_;
  wire _2743_;
  wire _2744_;
  wire _2745_;
  wire _2746_;
  wire _2747_;
  wire _2748_;
  wire _2749_;
  wire _2750_;
  wire _2751_;
  wire _2752_;
  wire _2753_;
  wire _2754_;
  wire _2755_;
  wire _2756_;
  wire _2757_;
  wire _2758_;
  wire _2759_;
  wire _2760_;
  wire _2761_;
  wire _2762_;
  wire _2763_;
  wire _2764_;
  wire _2765_;
  wire _2766_;
  wire _2767_;
  wire _2768_;
  wire _2769_;
  wire _2770_;
  wire _2771_;
  wire _2772_;
  wire _2773_;
  wire _2774_;
  wire _2775_;
  wire _2776_;
  wire _2777_;
  wire _2778_;
  wire _2779_;
  wire [15:0] _2780_;
  wire [15:0] _2781_;
  wire [15:0] _2782_;
  wire [15:0] _2783_;
  wire [15:0] _2784_;
  wire [15:0] _2785_;
  wire _2786_;
  wire _2787_;
  wire _2788_;
  wire _2789_;
  wire _2790_;
  wire _2791_;
  wire _2792_;
  wire _2793_;
  wire _2794_;
  wire _2795_;
  wire _2796_;
  wire _2797_;
  wire _2798_;
  wire _2799_;
  wire _2800_;
  wire _2801_;
  wire _2802_;
  wire _2803_;
  wire _2804_;
  wire _2805_;
  wire _2806_;
  wire _2807_;
  wire _2808_;
  wire _2809_;
  wire _2810_;
  wire _2811_;
  wire _2812_;
  wire _2813_;
  wire _2814_;
  wire _2815_;
  wire _2816_;
  wire _2817_;
  wire _2818_;
  wire _2819_;
  wire _2820_;
  wire _2821_;
  wire _2822_;
  wire _2823_;
  wire _2824_;
  wire _2825_;
  wire _2826_;
  wire _2827_;
  wire _2828_;
  wire _2829_;
  wire _2830_;
  wire _2831_;
  wire _2832_;
  wire _2833_;
  wire _2834_;
  wire _2835_;
  wire _2836_;
  wire _2837_;
  wire _2838_;
  wire _2839_;
  wire _2840_;
  wire _2841_;
  wire _2842_;
  wire _2843_;
  wire _2844_;
  wire _2845_;
  wire _2846_;
  wire _2847_;
  wire _2848_;
  wire _2849_;
  wire _2850_;
  wire [15:0] _2851_;
  wire [15:0] _2852_;
  wire [15:0] _2853_;
  wire [15:0] _2854_;
  wire [15:0] _2855_;
  wire [15:0] _2856_;
  wire _2857_;
  wire _2858_;
  wire _2859_;
  wire _2860_;
  wire _2861_;
  wire _2862_;
  wire _2863_;
  wire _2864_;
  wire _2865_;
  wire _2866_;
  wire _2867_;
  wire _2868_;
  wire _2869_;
  wire _2870_;
  wire _2871_;
  wire _2872_;
  wire _2873_;
  wire _2874_;
  wire _2875_;
  wire _2876_;
  wire _2877_;
  wire _2878_;
  wire _2879_;
  wire _2880_;
  wire _2881_;
  wire _2882_;
  wire _2883_;
  wire _2884_;
  wire _2885_;
  wire _2886_;
  wire _2887_;
  wire _2888_;
  wire _2889_;
  wire _2890_;
  wire _2891_;
  wire _2892_;
  wire _2893_;
  wire _2894_;
  wire _2895_;
  wire _2896_;
  wire _2897_;
  wire _2898_;
  wire _2899_;
  wire _2900_;
  wire _2901_;
  wire _2902_;
  wire _2903_;
  wire _2904_;
  wire _2905_;
  wire _2906_;
  wire _2907_;
  wire _2908_;
  wire _2909_;
  wire _2910_;
  wire _2911_;
  wire _2912_;
  wire _2913_;
  wire _2914_;
  wire _2915_;
  wire _2916_;
  wire _2917_;
  wire _2918_;
  wire _2919_;
  wire _2920_;
  wire _2921_;
  wire [15:0] _2922_;
  wire [15:0] _2923_;
  wire [15:0] _2924_;
  wire [15:0] _2925_;
  wire [15:0] _2926_;
  wire [15:0] _2927_;
  wire _2928_;
  wire _2929_;
  wire _2930_;
  wire _2931_;
  wire _2932_;
  wire _2933_;
  wire _2934_;
  wire _2935_;
  wire _2936_;
  wire _2937_;
  wire _2938_;
  wire _2939_;
  wire _2940_;
  wire _2941_;
  wire _2942_;
  wire _2943_;
  wire _2944_;
  wire _2945_;
  wire _2946_;
  wire _2947_;
  wire _2948_;
  wire _2949_;
  wire _2950_;
  wire _2951_;
  wire _2952_;
  wire _2953_;
  wire _2954_;
  wire _2955_;
  wire _2956_;
  wire _2957_;
  wire _2958_;
  wire _2959_;
  wire _2960_;
  wire _2961_;
  wire _2962_;
  wire _2963_;
  wire _2964_;
  wire _2965_;
  wire _2966_;
  wire _2967_;
  wire _2968_;
  wire _2969_;
  wire _2970_;
  wire _2971_;
  wire _2972_;
  wire _2973_;
  wire _2974_;
  wire _2975_;
  wire _2976_;
  wire _2977_;
  wire _2978_;
  wire _2979_;
  wire _2980_;
  wire _2981_;
  wire _2982_;
  wire _2983_;
  wire _2984_;
  wire _2985_;
  wire _2986_;
  wire _2987_;
  wire _2988_;
  wire _2989_;
  wire _2990_;
  wire _2991_;
  wire _2992_;
  wire [15:0] _2993_;
  wire [15:0] _2994_;
  wire [15:0] _2995_;
  wire [15:0] _2996_;
  wire [15:0] _2997_;
  wire [15:0] _2998_;
  wire _2999_;
  wire _3000_;
  wire _3001_;
  wire _3002_;
  wire _3003_;
  wire _3004_;
  wire _3005_;
  wire _3006_;
  wire _3007_;
  wire _3008_;
  wire _3009_;
  wire _3010_;
  wire _3011_;
  wire _3012_;
  wire _3013_;
  wire _3014_;
  wire _3015_;
  wire _3016_;
  wire _3017_;
  wire _3018_;
  wire _3019_;
  wire _3020_;
  wire _3021_;
  wire _3022_;
  wire _3023_;
  wire _3024_;
  wire _3025_;
  wire _3026_;
  wire _3027_;
  wire _3028_;
  wire _3029_;
  wire _3030_;
  wire _3031_;
  wire _3032_;
  wire _3033_;
  wire _3034_;
  wire _3035_;
  wire _3036_;
  wire _3037_;
  wire _3038_;
  wire _3039_;
  wire _3040_;
  wire _3041_;
  wire _3042_;
  wire _3043_;
  wire _3044_;
  wire _3045_;
  wire _3046_;
  wire _3047_;
  wire _3048_;
  wire _3049_;
  wire _3050_;
  wire _3051_;
  wire _3052_;
  wire _3053_;
  wire _3054_;
  wire _3055_;
  wire _3056_;
  wire _3057_;
  wire _3058_;
  wire _3059_;
  wire _3060_;
  wire _3061_;
  wire _3062_;
  wire _3063_;
  wire [15:0] _3064_;
  wire [15:0] _3065_;
  wire [15:0] _3066_;
  wire [15:0] _3067_;
  wire [15:0] _3068_;
  wire [15:0] _3069_;
  wire _3070_;
  wire _3071_;
  wire _3072_;
  wire _3073_;
  wire _3074_;
  wire _3075_;
  wire _3076_;
  wire _3077_;
  wire _3078_;
  wire _3079_;
  wire _3080_;
  wire _3081_;
  wire _3082_;
  wire _3083_;
  wire _3084_;
  wire _3085_;
  wire _3086_;
  wire _3087_;
  wire _3088_;
  wire _3089_;
  wire _3090_;
  wire _3091_;
  wire _3092_;
  wire _3093_;
  wire _3094_;
  wire _3095_;
  wire _3096_;
  wire _3097_;
  wire _3098_;
  wire _3099_;
  wire _3100_;
  wire _3101_;
  wire _3102_;
  wire _3103_;
  wire _3104_;
  wire _3105_;
  wire _3106_;
  wire _3107_;
  wire _3108_;
  wire _3109_;
  wire _3110_;
  wire _3111_;
  wire _3112_;
  wire _3113_;
  wire _3114_;
  wire _3115_;
  wire _3116_;
  wire _3117_;
  wire _3118_;
  wire _3119_;
  wire _3120_;
  wire _3121_;
  wire _3122_;
  wire _3123_;
  wire _3124_;
  wire _3125_;
  wire _3126_;
  wire _3127_;
  wire _3128_;
  wire _3129_;
  wire _3130_;
  wire _3131_;
  wire _3132_;
  wire _3133_;
  wire _3134_;
  wire [15:0] _3135_;
  wire [15:0] _3136_;
  wire [15:0] _3137_;
  wire [15:0] _3138_;
  wire [15:0] _3139_;
  wire [15:0] _3140_;
  wire _3141_;
  wire _3142_;
  wire _3143_;
  wire _3144_;
  wire _3145_;
  wire _3146_;
  wire _3147_;
  wire _3148_;
  wire _3149_;
  wire _3150_;
  wire _3151_;
  wire _3152_;
  wire _3153_;
  wire _3154_;
  wire _3155_;
  wire _3156_;
  wire _3157_;
  wire _3158_;
  wire _3159_;
  wire _3160_;
  wire _3161_;
  wire _3162_;
  wire _3163_;
  wire _3164_;
  wire _3165_;
  wire _3166_;
  wire _3167_;
  wire _3168_;
  wire _3169_;
  wire _3170_;
  wire _3171_;
  wire _3172_;
  wire _3173_;
  wire _3174_;
  wire _3175_;
  wire _3176_;
  wire _3177_;
  wire _3178_;
  wire _3179_;
  wire _3180_;
  wire _3181_;
  wire _3182_;
  wire _3183_;
  wire _3184_;
  wire _3185_;
  wire _3186_;
  wire _3187_;
  wire _3188_;
  wire _3189_;
  wire _3190_;
  wire _3191_;
  wire _3192_;
  wire _3193_;
  wire _3194_;
  wire _3195_;
  wire _3196_;
  wire _3197_;
  wire _3198_;
  wire _3199_;
  wire _3200_;
  wire _3201_;
  wire _3202_;
  wire _3203_;
  wire _3204_;
  wire _3205_;
  wire [15:0] _3206_;
  wire [15:0] _3207_;
  wire [15:0] _3208_;
  wire [15:0] _3209_;
  wire [15:0] _3210_;
  wire [15:0] _3211_;
  wire _3212_;
  wire _3213_;
  wire _3214_;
  wire _3215_;
  wire _3216_;
  wire _3217_;
  wire _3218_;
  wire _3219_;
  wire _3220_;
  wire _3221_;
  wire _3222_;
  wire _3223_;
  wire _3224_;
  wire _3225_;
  wire _3226_;
  wire _3227_;
  wire _3228_;
  wire _3229_;
  wire _3230_;
  wire _3231_;
  wire _3232_;
  wire _3233_;
  wire _3234_;
  wire _3235_;
  wire _3236_;
  wire _3237_;
  wire _3238_;
  wire _3239_;
  wire _3240_;
  wire _3241_;
  wire _3242_;
  wire _3243_;
  wire _3244_;
  wire _3245_;
  wire _3246_;
  wire _3247_;
  wire _3248_;
  wire _3249_;
  wire _3250_;
  wire _3251_;
  wire _3252_;
  wire _3253_;
  wire _3254_;
  wire _3255_;
  wire _3256_;
  wire _3257_;
  wire _3258_;
  wire _3259_;
  wire _3260_;
  wire _3261_;
  wire _3262_;
  wire _3263_;
  wire _3264_;
  wire _3265_;
  wire _3266_;
  wire _3267_;
  wire _3268_;
  wire _3269_;
  wire _3270_;
  wire _3271_;
  wire _3272_;
  wire _3273_;
  wire _3274_;
  wire _3275_;
  wire _3276_;
  wire [15:0] _3277_;
  wire [15:0] _3278_;
  wire [15:0] _3279_;
  wire [15:0] _3280_;
  wire [15:0] _3281_;
  wire [15:0] _3282_;
  wire _3283_;
  wire _3284_;
  wire _3285_;
  wire _3286_;
  wire _3287_;
  wire _3288_;
  wire _3289_;
  wire _3290_;
  wire _3291_;
  wire _3292_;
  wire _3293_;
  wire _3294_;
  wire _3295_;
  wire _3296_;
  wire _3297_;
  wire _3298_;
  wire _3299_;
  wire _3300_;
  wire _3301_;
  wire _3302_;
  wire _3303_;
  wire _3304_;
  wire _3305_;
  wire _3306_;
  wire _3307_;
  wire _3308_;
  wire _3309_;
  wire _3310_;
  wire _3311_;
  wire _3312_;
  wire _3313_;
  wire _3314_;
  wire _3315_;
  wire _3316_;
  wire _3317_;
  wire _3318_;
  wire _3319_;
  wire _3320_;
  wire _3321_;
  wire _3322_;
  wire _3323_;
  wire _3324_;
  wire _3325_;
  wire _3326_;
  wire _3327_;
  wire _3328_;
  wire _3329_;
  wire _3330_;
  wire _3331_;
  wire _3332_;
  wire _3333_;
  wire _3334_;
  wire _3335_;
  wire _3336_;
  wire _3337_;
  wire _3338_;
  wire _3339_;
  wire _3340_;
  wire _3341_;
  wire _3342_;
  wire _3343_;
  wire _3344_;
  wire _3345_;
  wire _3346_;
  wire _3347_;
  wire [15:0] _3348_;
  wire [15:0] _3349_;
  wire [15:0] _3350_;
  wire [15:0] _3351_;
  wire [15:0] _3352_;
  wire _3353_;
  wire _3354_;
  wire [1:0] _3355_;
  wire _3356_;
  wire [2:0] _3357_;
  wire _3358_;
  wire _3359_;
  wire _3360_;
  wire [1:0] _3361_;
  wire _3362_;
  wire [2:0] _3363_;
  wire _3364_;
  wire _3365_;
  wire _3366_;
  wire [1:0] _3367_;
  wire _3368_;
  wire [2:0] _3369_;
  wire _3370_;
  wire _3371_;
  wire _3372_;
  wire [1:0] _3373_;
  wire _3374_;
  wire [2:0] _3375_;
  wire _3376_;
  wire _3377_;
  wire _3378_;
  wire [1:0] _3379_;
  wire _3380_;
  wire [2:0] _3381_;
  wire _3382_;
  wire _3383_;
  wire _3384_;
  wire [1:0] _3385_;
  wire _3386_;
  wire [2:0] _3387_;
  wire _3388_;
  wire _3389_;
  wire _3390_;
  wire [1:0] _3391_;
  wire _3392_;
  wire [2:0] _3393_;
  wire _3394_;
  wire _3395_;
  wire _3396_;
  wire [1:0] _3397_;
  wire _3398_;
  wire [2:0] _3399_;
  wire _3400_;
  wire [1:0] _3401_;
  wire _3402_;
  wire [1:0] _3403_;
  wire _3404_;
  wire [1:0] _3405_;
  wire _3406_;
  wire [1:0] _3407_;
  wire _3408_;
  wire [1:0] _3409_;
  wire _3410_;
  wire [1:0] _3411_;
  wire _3412_;
  wire [1:0] _3413_;
  wire _3414_;
  wire [1:0] _3415_;
  wire _3416_;
  wire [15:0] _3417_;
  wire [15:0] _3418_;
  wire [15:0] _3419_;
  wire [15:0] _3420_;
  wire [15:0] _3421_;
  wire [15:0] _3422_;
  wire [15:0] _3423_;
  wire [15:0] _3424_;
  wire [15:0] _3425_;
  wire [15:0] _3426_;
  wire [15:0] _3427_;
  wire [15:0] _3428_;
  wire [15:0] _3429_;
  wire [15:0] _3430_;
  wire [15:0] _3431_;
  wire [15:0] _3432_;
  wire [15:0] _3433_;
  wire [15:0] _3434_;
  wire [15:0] _3435_;
  wire [15:0] _3436_;
  wire [15:0] _3437_;
  wire [15:0] _3438_;
  wire [15:0] _3439_;
  wire [15:0] _3440_;
  wire [15:0] _3441_;
  wire [15:0] _3442_;
  wire [15:0] _3443_;
  wire [15:0] _3444_;
  wire [15:0] _3445_;
  wire [15:0] _3446_;
  wire [15:0] _3447_;
  wire [15:0] _3448_;
  wire [15:0] _3449_;
  wire [15:0] _3450_;
  wire [15:0] _3451_;
  wire [15:0] _3452_;
  wire [15:0] _3453_;
  wire [15:0] _3454_;
  wire [15:0] _3455_;
  wire [15:0] _3456_;
  wire [15:0] _3457_;
  wire [15:0] _3458_;
  wire [15:0] _3459_;
  wire [15:0] _3460_;
  wire [15:0] _3461_;
  wire [15:0] _3462_;
  wire [15:0] _3463_;
  wire [15:0] _3464_;
  wire [15:0] _3465_;
  wire [15:0] _3466_;
  wire [15:0] _3467_;
  wire [15:0] _3468_;
  wire [15:0] _3469_;
  wire [15:0] _3470_;
  wire [15:0] _3471_;
  wire [15:0] _3472_;
  wire [15:0] _3473_;
  wire [15:0] _3474_;
  wire [15:0] _3475_;
  wire [15:0] _3476_;
  wire [15:0] _3477_;
  wire [15:0] _3478_;
  wire [15:0] _3479_;
  wire [15:0] _3480_;
  wire [15:0] _3481_;
  wire [15:0] _3482_;
  wire [15:0] _3483_;
  wire [15:0] _3484_;
  wire [15:0] _3485_;
  wire [15:0] _3486_;
  wire [15:0] _3487_;
  wire [15:0] _3488_;
  wire [15:0] _3489_;
  wire [15:0] _3490_;
  wire [15:0] _3491_;
  wire [15:0] _3492_;
  wire [15:0] _3493_;
  wire [15:0] _3494_;
  wire [15:0] _3495_;
  wire [15:0] _3496_;
  wire [15:0] _3497_;
  wire [15:0] _3498_;
  wire [15:0] _3499_;
  wire [15:0] _3500_;
  wire [15:0] _3501_;
  wire [15:0] _3502_;
  wire [15:0] _3503_;
  wire [15:0] _3504_;
  wire [15:0] _3505_;
  wire [15:0] _3506_;
  wire [15:0] _3507_;
  wire [15:0] _3508_;
  wire [15:0] _3509_;
  wire [15:0] _3510_;
  wire [15:0] _3511_;
  wire [15:0] _3512_;
  wire [15:0] _3513_;
  wire [15:0] _3514_;
  wire [15:0] _3515_;
  wire [15:0] _3516_;
  wire [15:0] _3517_;
  wire [15:0] _3518_;
  wire [15:0] _3519_;
  wire [15:0] _3520_;
  wire [15:0] _3521_;
  wire [15:0] _3522_;
  wire [15:0] _3523_;
  wire [15:0] _3524_;
  wire [15:0] _3525_;
  wire [15:0] _3526_;
  wire [15:0] _3527_;
  wire [15:0] _3528_;
  wire [15:0] _3529_;
  wire [15:0] _3530_;
  wire [15:0] _3531_;
  wire [15:0] _3532_;
  wire [15:0] _3533_;
  wire [15:0] _3534_;
  wire [15:0] _3535_;
  wire [15:0] _3536_;
  wire [15:0] _3537_;
  wire [15:0] _3538_;
  wire [15:0] _3539_;
  wire [15:0] _3540_;
  wire [15:0] _3541_;
  wire [15:0] _3542_;
  wire [15:0] _3543_;
  wire [15:0] _3544_;
  wire [15:0] _3545_;
  wire [15:0] _3546_;
  wire [15:0] _3547_;
  wire [15:0] _3548_;
  wire [15:0] _3549_;
  wire [15:0] _3550_;
  wire [15:0] _3551_;
  wire [15:0] _3552_;
  wire [15:0] _3553_;
  wire [15:0] _3554_;
  wire [15:0] _3555_;
  wire [15:0] _3556_;
  wire [15:0] _3557_;
  wire [15:0] _3558_;
  wire [15:0] _3559_;
  wire [15:0] _3560_;
  wire [15:0] _3561_;
  wire [15:0] _3562_;
  wire [15:0] _3563_;
  wire [15:0] _3564_;
  wire [15:0] _3565_;
  wire [15:0] _3566_;
  wire [15:0] _3567_;
  wire [15:0] _3568_;
  wire [15:0] _3569_;
  wire [15:0] _3570_;
  wire [15:0] _3571_;
  wire [15:0] _3572_;
  wire [15:0] _3573_;
  wire [15:0] _3574_;
  wire [15:0] _3575_;
  wire [15:0] _3576_;
  wire [15:0] _3577_;
  wire [15:0] _3578_;
  wire [15:0] _3579_;
  wire [15:0] _3580_;
  wire [15:0] _3581_;
  wire [15:0] _3582_;
  wire [15:0] _3583_;
  wire [15:0] _3584_;
  wire [15:0] _3585_;
  wire [15:0] _3586_;
  wire [15:0] _3587_;
  wire [15:0] _3588_;
  wire [15:0] _3589_;
  wire [15:0] _3590_;
  wire [15:0] _3591_;
  wire [15:0] _3592_;
  wire [15:0] _3593_;
  wire [15:0] _3594_;
  wire [15:0] _3595_;
  wire [15:0] _3596_;
  wire [15:0] _3597_;
  wire [15:0] _3598_;
  wire [15:0] _3599_;
  wire [15:0] _3600_;
  wire [15:0] _3601_;
  wire [15:0] _3602_;
  wire [15:0] _3603_;
  wire [15:0] _3604_;
  wire [15:0] _3605_;
  wire [15:0] _3606_;
  wire [15:0] _3607_;
  wire [15:0] _3608_;
  wire [15:0] _3609_;
  wire [15:0] _3610_;
  wire [15:0] _3611_;
  wire [15:0] _3612_;
  wire [15:0] _3613_;
  wire [15:0] _3614_;
  wire [15:0] _3615_;
  wire [15:0] _3616_;
  wire [15:0] _3617_;
  wire [15:0] _3618_;
  wire [15:0] _3619_;
  wire [15:0] _3620_;
  wire [15:0] _3621_;
  wire [15:0] _3622_;
  wire [15:0] _3623_;
  wire [15:0] _3624_;
  wire [15:0] _3625_;
  wire [15:0] _3626_;
  wire [15:0] _3627_;
  wire [15:0] _3628_;
  wire [15:0] _3629_;
  wire [15:0] _3630_;
  wire [15:0] _3631_;
  wire [15:0] _3632_;
  wire [15:0] _3633_;
  wire [15:0] _3634_;
  wire [15:0] _3635_;
  wire [15:0] _3636_;
  wire [15:0] _3637_;
  wire [15:0] _3638_;
  wire [15:0] _3639_;
  wire [15:0] _3640_;
  wire [15:0] _3641_;
  wire [15:0] _3642_;
  wire [15:0] _3643_;
  wire [15:0] _3644_;
  wire [15:0] _3645_;
  wire [15:0] _3646_;
  wire [15:0] _3647_;
  wire [15:0] _3648_;
  wire [15:0] _3649_;
  wire [15:0] _3650_;
  wire [15:0] _3651_;
  wire [15:0] _3652_;
  wire [15:0] _3653_;
  wire [15:0] _3654_;
  wire [15:0] _3655_;
  wire [15:0] _3656_;
  wire [15:0] _3657_;
  wire [15:0] _3658_;
  wire [15:0] _3659_;
  wire [15:0] _3660_;
  wire [15:0] _3661_;
  wire [15:0] _3662_;
  wire [15:0] _3663_;
  wire [15:0] _3664_;
  wire [15:0] _3665_;
  wire [15:0] _3666_;
  wire [15:0] _3667_;
  wire [15:0] _3668_;
  wire [15:0] _3669_;
  wire [15:0] _3670_;
  wire [15:0] _3671_;
  wire [15:0] _3672_;
  wire [15:0] _3673_;
  wire [15:0] _3674_;
  wire [15:0] _3675_;
  wire [15:0] _3676_;
  wire [15:0] _3677_;
  wire [15:0] _3678_;
  wire [15:0] _3679_;
  wire [15:0] _3680_;
  wire [15:0] _3681_;
  wire [15:0] _3682_;
  wire [15:0] _3683_;
  wire [15:0] _3684_;
  wire [15:0] _3685_;
  wire [15:0] _3686_;
  wire [15:0] _3687_;
  wire [15:0] _3688_;
  wire [15:0] _3689_;
  wire [15:0] _3690_;
  wire [15:0] _3691_;
  wire [15:0] _3692_;
  wire [15:0] _3693_;
  wire [15:0] _3694_;
  wire [15:0] _3695_;
  wire [15:0] _3696_;
  wire [15:0] _3697_;
  wire [15:0] _3698_;
  wire [15:0] _3699_;
  wire [15:0] _3700_;
  wire [15:0] _3701_;
  wire [15:0] _3702_;
  wire [15:0] _3703_;
  wire [15:0] _3704_;
  wire [15:0] _3705_;
  wire [15:0] _3706_;
  wire [15:0] _3707_;
  wire [15:0] _3708_;
  wire [15:0] _3709_;
  wire [15:0] _3710_;
  wire [15:0] _3711_;
  wire [15:0] _3712_;
  wire [15:0] _3713_;
  wire [15:0] _3714_;
  wire [15:0] _3715_;
  wire [15:0] _3716_;
  wire [15:0] _3717_;
  wire [15:0] _3718_;
  wire [15:0] _3719_;
  wire [15:0] _3720_;
  wire [15:0] _3721_;
  wire [15:0] _3722_;
  wire [15:0] _3723_;
  wire [15:0] _3724_;
  wire [15:0] _3725_;
  wire [15:0] _3726_;
  wire [15:0] _3727_;
  wire [15:0] _3728_;
  wire [15:0] _3729_;
  wire [15:0] _3730_;
  wire [15:0] _3731_;
  wire [15:0] _3732_;
  wire [15:0] _3733_;
  wire [15:0] _3734_;
  wire [15:0] _3735_;
  wire [15:0] _3736_;
  wire [15:0] _3737_;
  wire [15:0] _3738_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:16763" *)
  wire _3739_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:16764" *)
  wire _3740_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:16765" *)
  wire _3741_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:16766" *)
  wire _3742_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:16863" *)
  wire _3743_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:16864" *)
  wire _3744_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:16865" *)
  wire _3745_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:16866" *)
  wire _3746_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:16716" *)
  wire [15:0] _3747_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:16717" *)
  wire [15:0] _3748_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:16718" *)
  wire [15:0] _3749_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:16719" *)
  wire [15:0] _3750_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:16720" *)
  wire [15:0] _3751_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:16721" *)
  wire [15:0] _3752_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:16722" *)
  wire [15:0] _3753_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:16723" *)
  wire [15:0] _3754_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:16724" *)
  wire [15:0] _3755_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:16725" *)
  wire [15:0] _3756_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:16726" *)
  wire [15:0] _3757_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:16727" *)
  wire [15:0] _3758_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:16728" *)
  wire [15:0] _3759_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:16729" *)
  wire [15:0] _3760_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:16730" *)
  wire [15:0] _3761_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:16731" *)
  wire [15:0] _3762_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:16732" *)
  wire [15:0] _3763_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:16733" *)
  wire [15:0] _3764_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:16734" *)
  wire [15:0] _3765_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:16735" *)
  wire [15:0] _3766_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:16736" *)
  wire [15:0] _3767_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:16737" *)
  wire [15:0] _3768_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:16738" *)
  wire [15:0] _3769_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:16739" *)
  wire [15:0] _3770_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:593" *)
  wire [3:0] FMcvt_in_rdy;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:594" *)
  wire [3:0] FMcvt_in_vld;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:595" *)
  wire [3:0] FMcvt_out_rdy;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:596" *)
  wire [3:0] FMcvt_out_vld;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:597" *)
  wire both_hybrid_sel;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:598" *)
  wire both_of_sel;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:599" *)
  wire both_uf_sel;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:181" *)
  reg [15:0] density_out;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:182" *)
  reg [15:0] density_reg0;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:183" *)
  reg [15:0] density_reg1;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:184" *)
  reg [15:0] density_reg10;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:185" *)
  reg [15:0] density_reg100;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:186" *)
  reg [15:0] density_reg101;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:187" *)
  reg [15:0] density_reg102;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:188" *)
  reg [15:0] density_reg103;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:189" *)
  reg [15:0] density_reg104;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:190" *)
  reg [15:0] density_reg105;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:191" *)
  reg [15:0] density_reg106;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:192" *)
  reg [15:0] density_reg107;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:193" *)
  reg [15:0] density_reg108;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:194" *)
  reg [15:0] density_reg109;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:195" *)
  reg [15:0] density_reg11;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:196" *)
  reg [15:0] density_reg110;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:197" *)
  reg [15:0] density_reg111;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:198" *)
  reg [15:0] density_reg112;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:199" *)
  reg [15:0] density_reg113;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:200" *)
  reg [15:0] density_reg114;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:201" *)
  reg [15:0] density_reg115;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:202" *)
  reg [15:0] density_reg116;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:203" *)
  reg [15:0] density_reg117;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:204" *)
  reg [15:0] density_reg118;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:205" *)
  reg [15:0] density_reg119;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:206" *)
  reg [15:0] density_reg12;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:207" *)
  reg [15:0] density_reg120;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:208" *)
  reg [15:0] density_reg121;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:209" *)
  reg [15:0] density_reg122;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:210" *)
  reg [15:0] density_reg123;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:211" *)
  reg [15:0] density_reg124;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:212" *)
  reg [15:0] density_reg125;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:213" *)
  reg [15:0] density_reg126;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:214" *)
  reg [15:0] density_reg127;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:215" *)
  reg [15:0] density_reg128;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:216" *)
  reg [15:0] density_reg129;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:217" *)
  reg [15:0] density_reg13;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:218" *)
  reg [15:0] density_reg130;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:219" *)
  reg [15:0] density_reg131;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:220" *)
  reg [15:0] density_reg132;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:221" *)
  reg [15:0] density_reg133;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:222" *)
  reg [15:0] density_reg134;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:223" *)
  reg [15:0] density_reg135;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:224" *)
  reg [15:0] density_reg136;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:225" *)
  reg [15:0] density_reg137;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:226" *)
  reg [15:0] density_reg138;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:227" *)
  reg [15:0] density_reg139;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:228" *)
  reg [15:0] density_reg14;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:229" *)
  reg [15:0] density_reg140;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:230" *)
  reg [15:0] density_reg141;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:231" *)
  reg [15:0] density_reg142;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:232" *)
  reg [15:0] density_reg143;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:233" *)
  reg [15:0] density_reg144;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:234" *)
  reg [15:0] density_reg145;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:235" *)
  reg [15:0] density_reg146;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:236" *)
  reg [15:0] density_reg147;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:237" *)
  reg [15:0] density_reg148;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:238" *)
  reg [15:0] density_reg149;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:239" *)
  reg [15:0] density_reg15;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:240" *)
  reg [15:0] density_reg150;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:241" *)
  reg [15:0] density_reg151;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:242" *)
  reg [15:0] density_reg152;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:243" *)
  reg [15:0] density_reg153;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:244" *)
  reg [15:0] density_reg154;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:245" *)
  reg [15:0] density_reg155;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:246" *)
  reg [15:0] density_reg156;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:247" *)
  reg [15:0] density_reg157;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:248" *)
  reg [15:0] density_reg158;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:249" *)
  reg [15:0] density_reg159;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:250" *)
  reg [15:0] density_reg16;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:251" *)
  reg [15:0] density_reg160;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:252" *)
  reg [15:0] density_reg161;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:253" *)
  reg [15:0] density_reg162;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:254" *)
  reg [15:0] density_reg163;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:255" *)
  reg [15:0] density_reg164;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:256" *)
  reg [15:0] density_reg165;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:257" *)
  reg [15:0] density_reg166;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:258" *)
  reg [15:0] density_reg167;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:259" *)
  reg [15:0] density_reg168;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:260" *)
  reg [15:0] density_reg169;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:261" *)
  reg [15:0] density_reg17;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:262" *)
  reg [15:0] density_reg170;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:263" *)
  reg [15:0] density_reg171;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:264" *)
  reg [15:0] density_reg172;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:265" *)
  reg [15:0] density_reg173;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:266" *)
  reg [15:0] density_reg174;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:267" *)
  reg [15:0] density_reg175;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:268" *)
  reg [15:0] density_reg176;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:269" *)
  reg [15:0] density_reg177;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:270" *)
  reg [15:0] density_reg178;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:271" *)
  reg [15:0] density_reg179;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:272" *)
  reg [15:0] density_reg18;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:273" *)
  reg [15:0] density_reg180;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:274" *)
  reg [15:0] density_reg181;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:275" *)
  reg [15:0] density_reg182;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:276" *)
  reg [15:0] density_reg183;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:277" *)
  reg [15:0] density_reg184;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:278" *)
  reg [15:0] density_reg185;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:279" *)
  reg [15:0] density_reg186;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:280" *)
  reg [15:0] density_reg187;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:281" *)
  reg [15:0] density_reg188;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:282" *)
  reg [15:0] density_reg189;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:283" *)
  reg [15:0] density_reg19;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:284" *)
  reg [15:0] density_reg190;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:285" *)
  reg [15:0] density_reg191;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:286" *)
  reg [15:0] density_reg192;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:287" *)
  reg [15:0] density_reg193;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:288" *)
  reg [15:0] density_reg194;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:289" *)
  reg [15:0] density_reg195;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:290" *)
  reg [15:0] density_reg196;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:291" *)
  reg [15:0] density_reg197;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:292" *)
  reg [15:0] density_reg198;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:293" *)
  reg [15:0] density_reg199;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:294" *)
  reg [15:0] density_reg2;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:295" *)
  reg [15:0] density_reg20;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:296" *)
  reg [15:0] density_reg200;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:297" *)
  reg [15:0] density_reg201;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:298" *)
  reg [15:0] density_reg202;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:299" *)
  reg [15:0] density_reg203;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:300" *)
  reg [15:0] density_reg204;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:301" *)
  reg [15:0] density_reg205;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:302" *)
  reg [15:0] density_reg206;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:303" *)
  reg [15:0] density_reg207;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:304" *)
  reg [15:0] density_reg208;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:305" *)
  reg [15:0] density_reg209;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:306" *)
  reg [15:0] density_reg21;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:307" *)
  reg [15:0] density_reg210;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:308" *)
  reg [15:0] density_reg211;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:309" *)
  reg [15:0] density_reg212;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:310" *)
  reg [15:0] density_reg213;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:311" *)
  reg [15:0] density_reg214;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:312" *)
  reg [15:0] density_reg215;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:313" *)
  reg [15:0] density_reg216;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:314" *)
  reg [15:0] density_reg217;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:315" *)
  reg [15:0] density_reg218;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:316" *)
  reg [15:0] density_reg219;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:317" *)
  reg [15:0] density_reg22;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:318" *)
  reg [15:0] density_reg220;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:319" *)
  reg [15:0] density_reg221;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:320" *)
  reg [15:0] density_reg222;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:321" *)
  reg [15:0] density_reg223;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:322" *)
  reg [15:0] density_reg224;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:323" *)
  reg [15:0] density_reg225;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:324" *)
  reg [15:0] density_reg226;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:325" *)
  reg [15:0] density_reg227;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:326" *)
  reg [15:0] density_reg228;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:327" *)
  reg [15:0] density_reg229;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:328" *)
  reg [15:0] density_reg23;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:329" *)
  reg [15:0] density_reg230;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:330" *)
  reg [15:0] density_reg231;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:331" *)
  reg [15:0] density_reg232;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:332" *)
  reg [15:0] density_reg233;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:333" *)
  reg [15:0] density_reg234;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:334" *)
  reg [15:0] density_reg235;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:335" *)
  reg [15:0] density_reg236;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:336" *)
  reg [15:0] density_reg237;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:337" *)
  reg [15:0] density_reg238;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:338" *)
  reg [15:0] density_reg239;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:339" *)
  reg [15:0] density_reg24;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:340" *)
  reg [15:0] density_reg240;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:341" *)
  reg [15:0] density_reg241;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:342" *)
  reg [15:0] density_reg242;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:343" *)
  reg [15:0] density_reg243;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:344" *)
  reg [15:0] density_reg244;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:345" *)
  reg [15:0] density_reg245;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:346" *)
  reg [15:0] density_reg246;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:347" *)
  reg [15:0] density_reg247;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:348" *)
  reg [15:0] density_reg248;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:349" *)
  reg [15:0] density_reg249;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:350" *)
  reg [15:0] density_reg25;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:351" *)
  reg [15:0] density_reg250;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:352" *)
  reg [15:0] density_reg251;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:353" *)
  reg [15:0] density_reg252;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:354" *)
  reg [15:0] density_reg253;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:355" *)
  reg [15:0] density_reg254;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:356" *)
  reg [15:0] density_reg255;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:357" *)
  reg [15:0] density_reg256;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:358" *)
  reg [15:0] density_reg26;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:359" *)
  reg [15:0] density_reg27;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:360" *)
  reg [15:0] density_reg28;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:361" *)
  reg [15:0] density_reg29;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:362" *)
  reg [15:0] density_reg3;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:363" *)
  reg [15:0] density_reg30;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:364" *)
  reg [15:0] density_reg31;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:365" *)
  reg [15:0] density_reg32;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:366" *)
  reg [15:0] density_reg33;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:367" *)
  reg [15:0] density_reg34;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:368" *)
  reg [15:0] density_reg35;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:369" *)
  reg [15:0] density_reg36;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:370" *)
  reg [15:0] density_reg37;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:371" *)
  reg [15:0] density_reg38;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:372" *)
  reg [15:0] density_reg39;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:373" *)
  reg [15:0] density_reg4;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:374" *)
  reg [15:0] density_reg40;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:375" *)
  reg [15:0] density_reg41;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:376" *)
  reg [15:0] density_reg42;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:377" *)
  reg [15:0] density_reg43;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:378" *)
  reg [15:0] density_reg44;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:379" *)
  reg [15:0] density_reg45;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:380" *)
  reg [15:0] density_reg46;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:381" *)
  reg [15:0] density_reg47;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:382" *)
  reg [15:0] density_reg48;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:383" *)
  reg [15:0] density_reg49;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:384" *)
  reg [15:0] density_reg5;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:385" *)
  reg [15:0] density_reg50;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:386" *)
  reg [15:0] density_reg51;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:387" *)
  reg [15:0] density_reg52;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:388" *)
  reg [15:0] density_reg53;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:389" *)
  reg [15:0] density_reg54;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:390" *)
  reg [15:0] density_reg55;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:391" *)
  reg [15:0] density_reg56;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:392" *)
  reg [15:0] density_reg57;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:393" *)
  reg [15:0] density_reg58;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:394" *)
  reg [15:0] density_reg59;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:395" *)
  reg [15:0] density_reg6;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:396" *)
  reg [15:0] density_reg60;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:397" *)
  reg [15:0] density_reg61;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:398" *)
  reg [15:0] density_reg62;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:399" *)
  reg [15:0] density_reg63;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:400" *)
  reg [15:0] density_reg64;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:401" *)
  reg [15:0] density_reg65;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:402" *)
  reg [15:0] density_reg66;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:403" *)
  reg [15:0] density_reg67;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:404" *)
  reg [15:0] density_reg68;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:405" *)
  reg [15:0] density_reg69;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:406" *)
  reg [15:0] density_reg7;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:407" *)
  reg [15:0] density_reg70;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:408" *)
  reg [15:0] density_reg71;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:409" *)
  reg [15:0] density_reg72;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:410" *)
  reg [15:0] density_reg73;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:411" *)
  reg [15:0] density_reg74;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:412" *)
  reg [15:0] density_reg75;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:413" *)
  reg [15:0] density_reg76;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:414" *)
  reg [15:0] density_reg77;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:415" *)
  reg [15:0] density_reg78;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:416" *)
  reg [15:0] density_reg79;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:417" *)
  reg [15:0] density_reg8;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:418" *)
  reg [15:0] density_reg80;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:419" *)
  reg [15:0] density_reg81;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:420" *)
  reg [15:0] density_reg82;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:421" *)
  reg [15:0] density_reg83;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:422" *)
  reg [15:0] density_reg84;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:423" *)
  reg [15:0] density_reg85;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:424" *)
  reg [15:0] density_reg86;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:425" *)
  reg [15:0] density_reg87;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:426" *)
  reg [15:0] density_reg88;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:427" *)
  reg [15:0] density_reg89;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:428" *)
  reg [15:0] density_reg9;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:429" *)
  reg [15:0] density_reg90;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:430" *)
  reg [15:0] density_reg91;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:431" *)
  reg [15:0] density_reg92;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:432" *)
  reg [15:0] density_reg93;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:433" *)
  reg [15:0] density_reg94;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:434" *)
  reg [15:0] density_reg95;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:435" *)
  reg [15:0] density_reg96;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:436" *)
  reg [15:0] density_reg97;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:437" *)
  reg [15:0] density_reg98;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:438" *)
  reg [15:0] density_reg99;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:99" *)
  input [9:0] dp2lut_X_entry_0;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:100" *)
  input [9:0] dp2lut_X_entry_1;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:101" *)
  input [9:0] dp2lut_X_entry_2;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:102" *)
  input [9:0] dp2lut_X_entry_3;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:103" *)
  input [9:0] dp2lut_X_entry_4;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:104" *)
  input [9:0] dp2lut_X_entry_5;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:105" *)
  input [9:0] dp2lut_X_entry_6;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:106" *)
  input [9:0] dp2lut_X_entry_7;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:107" *)
  input [17:0] dp2lut_Xinfo_0;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:108" *)
  input [17:0] dp2lut_Xinfo_1;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:109" *)
  input [17:0] dp2lut_Xinfo_2;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:110" *)
  input [17:0] dp2lut_Xinfo_3;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:111" *)
  input [17:0] dp2lut_Xinfo_4;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:112" *)
  input [17:0] dp2lut_Xinfo_5;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:113" *)
  input [17:0] dp2lut_Xinfo_6;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:114" *)
  input [17:0] dp2lut_Xinfo_7;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:115" *)
  input [9:0] dp2lut_Y_entry_0;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:116" *)
  input [9:0] dp2lut_Y_entry_1;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:117" *)
  input [9:0] dp2lut_Y_entry_2;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:118" *)
  input [9:0] dp2lut_Y_entry_3;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:119" *)
  input [9:0] dp2lut_Y_entry_4;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:120" *)
  input [9:0] dp2lut_Y_entry_5;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:121" *)
  input [9:0] dp2lut_Y_entry_6;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:122" *)
  input [9:0] dp2lut_Y_entry_7;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:123" *)
  input [17:0] dp2lut_Yinfo_0;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:124" *)
  input [17:0] dp2lut_Yinfo_1;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:125" *)
  input [17:0] dp2lut_Yinfo_2;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:126" *)
  input [17:0] dp2lut_Yinfo_3;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:127" *)
  input [17:0] dp2lut_Yinfo_4;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:128" *)
  input [17:0] dp2lut_Yinfo_5;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:129" *)
  input [17:0] dp2lut_Yinfo_6;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:130" *)
  input [17:0] dp2lut_Yinfo_7;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:144" *)
  output dp2lut_prdy;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:600" *)
  wire dp2lut_prdy_f;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:131" *)
  input dp2lut_pvld;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:145" *)
  output [15:0] dp2reg_lut_data;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:439" *)
  reg fp16_en_f;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:601" *)
  wire fp_lut_prdy_f;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:602" *)
  wire fp_lut_pvld_f;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:603" *)
  wire fp_out_prdy;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:604" *)
  wire fp_out_vld;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:132" *)
  input int8_en;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:605" *)
  wire load_din;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:146" *)
  output [31:0] lut2intp_X_data_00;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:147" *)
  output [16:0] lut2intp_X_data_00_17b;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:148" *)
  output [31:0] lut2intp_X_data_01;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:149" *)
  output [31:0] lut2intp_X_data_10;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:150" *)
  output [16:0] lut2intp_X_data_10_17b;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:151" *)
  output [31:0] lut2intp_X_data_11;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:152" *)
  output [31:0] lut2intp_X_data_20;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:153" *)
  output [16:0] lut2intp_X_data_20_17b;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:154" *)
  output [31:0] lut2intp_X_data_21;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:155" *)
  output [31:0] lut2intp_X_data_30;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:156" *)
  output [16:0] lut2intp_X_data_30_17b;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:157" *)
  output [31:0] lut2intp_X_data_31;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:158" *)
  output [31:0] lut2intp_X_data_40;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:159" *)
  output [16:0] lut2intp_X_data_40_17b;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:160" *)
  output [31:0] lut2intp_X_data_41;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:161" *)
  output [31:0] lut2intp_X_data_50;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:162" *)
  output [16:0] lut2intp_X_data_50_17b;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:163" *)
  output [31:0] lut2intp_X_data_51;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:164" *)
  output [31:0] lut2intp_X_data_60;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:165" *)
  output [16:0] lut2intp_X_data_60_17b;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:166" *)
  output [31:0] lut2intp_X_data_61;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:167" *)
  output [31:0] lut2intp_X_data_70;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:168" *)
  output [16:0] lut2intp_X_data_70_17b;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:169" *)
  output [31:0] lut2intp_X_data_71;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:170" *)
  output [19:0] lut2intp_X_info_0;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:171" *)
  output [19:0] lut2intp_X_info_1;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:172" *)
  output [19:0] lut2intp_X_info_2;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:173" *)
  output [19:0] lut2intp_X_info_3;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:174" *)
  output [19:0] lut2intp_X_info_4;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:175" *)
  output [19:0] lut2intp_X_info_5;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:176" *)
  output [19:0] lut2intp_X_info_6;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:177" *)
  output [19:0] lut2intp_X_info_7;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:178" *)
  output [7:0] lut2intp_X_sel;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:179" *)
  output [7:0] lut2intp_Y_sel;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:133" *)
  input lut2intp_prdy;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:180" *)
  output lut2intp_pvld;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:606" *)
  wire [15:0] lutX_data_00;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:607" *)
  wire [15:0] lutX_data_01;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:608" *)
  wire [15:0] lutX_data_10;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:609" *)
  wire [15:0] lutX_data_11;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:610" *)
  wire [15:0] lutX_data_20;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:611" *)
  wire [15:0] lutX_data_21;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:612" *)
  wire [15:0] lutX_data_30;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:613" *)
  wire [15:0] lutX_data_31;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:614" *)
  wire [15:0] lutX_data_40;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:615" *)
  wire [15:0] lutX_data_41;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:616" *)
  wire [15:0] lutX_data_50;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:617" *)
  wire [15:0] lutX_data_51;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:618" *)
  wire [15:0] lutX_data_60;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:619" *)
  wire [15:0] lutX_data_61;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:620" *)
  wire [15:0] lutX_data_70;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:621" *)
  wire [15:0] lutX_data_71;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:622" *)
  wire [15:0] lutX_info_0;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:623" *)
  wire [15:0] lutX_info_1;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:624" *)
  wire [15:0] lutX_info_2;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:625" *)
  wire [15:0] lutX_info_3;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:626" *)
  wire [15:0] lutX_info_4;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:627" *)
  wire [15:0] lutX_info_5;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:628" *)
  wire [15:0] lutX_info_6;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:629" *)
  wire [15:0] lutX_info_7;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:474" *)
  reg [7:0] lutX_sel;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:630" *)
  wire [3:0] lutX_sel_o;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:475" *)
  reg [7:0] lutY_sel;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:631" *)
  wire [3:0] lutY_sel_o;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:632" *)
  wire [31:0] lut_X_dat_00;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:633" *)
  wire [16:0] lut_X_dat_00_fp17;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:634" *)
  wire [31:0] lut_X_dat_01;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:635" *)
  wire [31:0] lut_X_dat_10;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:636" *)
  wire [16:0] lut_X_dat_10_fp17;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:637" *)
  wire [31:0] lut_X_dat_11;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:638" *)
  wire [31:0] lut_X_dat_20;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:639" *)
  wire [16:0] lut_X_dat_20_fp17;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:640" *)
  wire [31:0] lut_X_dat_21;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:641" *)
  wire [31:0] lut_X_dat_30;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:642" *)
  wire [16:0] lut_X_dat_30_fp17;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:643" *)
  wire [31:0] lut_X_dat_31;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:476" *)
  reg [15:0] lut_X_data_00;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:477" *)
  reg [15:0] lut_X_data_01;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:478" *)
  reg [15:0] lut_X_data_10;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:479" *)
  reg [15:0] lut_X_data_11;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:480" *)
  reg [15:0] lut_X_data_20;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:481" *)
  reg [15:0] lut_X_data_21;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:482" *)
  reg [15:0] lut_X_data_30;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:483" *)
  reg [15:0] lut_X_data_31;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:484" *)
  reg [15:0] lut_X_data_40;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:485" *)
  reg [15:0] lut_X_data_41;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:486" *)
  reg [15:0] lut_X_data_50;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:487" *)
  reg [15:0] lut_X_data_51;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:488" *)
  reg [15:0] lut_X_data_60;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:489" *)
  reg [15:0] lut_X_data_61;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:490" *)
  reg [15:0] lut_X_data_70;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:491" *)
  reg [15:0] lut_X_data_71;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:644" *)
  (* unused_bits = "16" *)
  wire [20:0] lut_X_inf_0;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:645" *)
  (* unused_bits = "16" *)
  wire [20:0] lut_X_inf_1;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:646" *)
  (* unused_bits = "16" *)
  wire [20:0] lut_X_inf_2;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:647" *)
  (* unused_bits = "16" *)
  wire [20:0] lut_X_inf_3;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:492" *)
  reg [17:0] lut_X_info_0;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:493" *)
  reg [17:0] lut_X_info_1;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:494" *)
  reg [17:0] lut_X_info_2;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:495" *)
  reg [17:0] lut_X_info_3;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:496" *)
  reg [17:0] lut_X_info_4;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:497" *)
  reg [17:0] lut_X_info_5;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:498" *)
  reg [17:0] lut_X_info_6;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:499" *)
  reg [17:0] lut_X_info_7;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:500" *)
  wire [7:0] lut_X_sel;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:501" *)
  reg [15:0] lut_Y_data_00;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:502" *)
  reg [15:0] lut_Y_data_01;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:503" *)
  reg [15:0] lut_Y_data_10;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:504" *)
  reg [15:0] lut_Y_data_11;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:505" *)
  reg [15:0] lut_Y_data_20;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:506" *)
  reg [15:0] lut_Y_data_21;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:507" *)
  reg [15:0] lut_Y_data_30;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:508" *)
  reg [15:0] lut_Y_data_31;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:509" *)
  reg [15:0] lut_Y_data_40;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:510" *)
  reg [15:0] lut_Y_data_41;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:511" *)
  reg [15:0] lut_Y_data_50;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:512" *)
  reg [15:0] lut_Y_data_51;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:513" *)
  reg [15:0] lut_Y_data_60;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:514" *)
  reg [15:0] lut_Y_data_61;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:515" *)
  reg [15:0] lut_Y_data_70;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:516" *)
  reg [15:0] lut_Y_data_71;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:517" *)
  reg [17:0] lut_Y_info_0;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:518" *)
  reg [17:0] lut_Y_info_1;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:519" *)
  reg [17:0] lut_Y_info_2;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:520" *)
  reg [17:0] lut_Y_info_3;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:521" *)
  reg [17:0] lut_Y_info_4;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:522" *)
  reg [17:0] lut_Y_info_5;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:523" *)
  reg [17:0] lut_Y_info_6;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:524" *)
  reg [17:0] lut_Y_info_7;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:525" *)
  wire [7:0] lut_Y_sel;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:648" *)
  wire lut_prdy;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:526" *)
  reg lut_pvld_f;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:649" *)
  wire lut_wr_en;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:96" *)
  input nvdla_core_clk;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:97" *)
  input nvdla_core_clk_orig;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:98" *)
  input nvdla_core_rstn;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:134" *)
  input nvdla_op_gated_clk_fp16;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:527" *)
  reg [15:0] raw_out;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:528" *)
  reg [15:0] raw_reg0;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:529" *)
  reg [15:0] raw_reg1;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:530" *)
  reg [15:0] raw_reg10;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:531" *)
  reg [15:0] raw_reg11;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:532" *)
  reg [15:0] raw_reg12;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:533" *)
  reg [15:0] raw_reg13;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:534" *)
  reg [15:0] raw_reg14;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:535" *)
  reg [15:0] raw_reg15;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:536" *)
  reg [15:0] raw_reg16;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:537" *)
  reg [15:0] raw_reg17;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:538" *)
  reg [15:0] raw_reg18;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:539" *)
  reg [15:0] raw_reg19;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:540" *)
  reg [15:0] raw_reg2;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:541" *)
  reg [15:0] raw_reg20;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:542" *)
  reg [15:0] raw_reg21;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:543" *)
  reg [15:0] raw_reg22;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:544" *)
  reg [15:0] raw_reg23;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:545" *)
  reg [15:0] raw_reg24;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:546" *)
  reg [15:0] raw_reg25;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:547" *)
  reg [15:0] raw_reg26;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:548" *)
  reg [15:0] raw_reg27;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:549" *)
  reg [15:0] raw_reg28;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:550" *)
  reg [15:0] raw_reg29;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:551" *)
  reg [15:0] raw_reg3;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:552" *)
  reg [15:0] raw_reg30;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:553" *)
  reg [15:0] raw_reg31;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:554" *)
  reg [15:0] raw_reg32;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:555" *)
  reg [15:0] raw_reg33;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:556" *)
  reg [15:0] raw_reg34;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:557" *)
  reg [15:0] raw_reg35;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:558" *)
  reg [15:0] raw_reg36;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:559" *)
  reg [15:0] raw_reg37;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:560" *)
  reg [15:0] raw_reg38;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:561" *)
  reg [15:0] raw_reg39;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:562" *)
  reg [15:0] raw_reg4;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:563" *)
  reg [15:0] raw_reg40;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:564" *)
  reg [15:0] raw_reg41;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:565" *)
  reg [15:0] raw_reg42;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:566" *)
  reg [15:0] raw_reg43;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:567" *)
  reg [15:0] raw_reg44;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:568" *)
  reg [15:0] raw_reg45;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:569" *)
  reg [15:0] raw_reg46;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:570" *)
  reg [15:0] raw_reg47;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:571" *)
  reg [15:0] raw_reg48;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:572" *)
  reg [15:0] raw_reg49;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:573" *)
  reg [15:0] raw_reg5;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:574" *)
  reg [15:0] raw_reg50;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:575" *)
  reg [15:0] raw_reg51;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:576" *)
  reg [15:0] raw_reg52;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:577" *)
  reg [15:0] raw_reg53;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:578" *)
  reg [15:0] raw_reg54;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:579" *)
  reg [15:0] raw_reg55;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:580" *)
  reg [15:0] raw_reg56;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:581" *)
  reg [15:0] raw_reg57;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:582" *)
  reg [15:0] raw_reg58;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:583" *)
  reg [15:0] raw_reg59;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:584" *)
  reg [15:0] raw_reg6;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:585" *)
  reg [15:0] raw_reg60;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:586" *)
  reg [15:0] raw_reg61;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:587" *)
  reg [15:0] raw_reg62;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:588" *)
  reg [15:0] raw_reg63;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:589" *)
  reg [15:0] raw_reg64;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:590" *)
  reg [15:0] raw_reg7;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:591" *)
  reg [15:0] raw_reg8;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:592" *)
  reg [15:0] raw_reg9;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:650" *)
  wire raw_select;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:135" *)
  input [1:0] reg2dp_input_data_type;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:136" *)
  input reg2dp_lut_access_type;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:137" *)
  input [9:0] reg2dp_lut_addr;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:138" *)
  input [15:0] reg2dp_lut_data;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:139" *)
  input reg2dp_lut_data_trigger;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:140" *)
  input reg2dp_lut_hybrid_priority;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:141" *)
  input reg2dp_lut_oflow_priority;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:142" *)
  input reg2dp_lut_table_id;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:143" *)
  input reg2dp_lut_uflow_priority;
  assign _0384_ = lut_wr_en & (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1001" *) raw_select;
  assign _0385_ = load_din & (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10368" *) lut_Y_sel[3];
  assign _0386_ = load_din & (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11419" *) int8_en;
  assign _0387_ = _0386_ & (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11419" *) lut_Y_sel[4];
  assign _0388_ = _0386_ & (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12470" *) lut_Y_sel[5];
  assign _0389_ = lut_wr_en & (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1322" *) reg2dp_lut_table_id;
  assign _0390_ = _0386_ & (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13521" *) lut_Y_sel[6];
  assign _0391_ = _0386_ & (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14572" *) lut_Y_sel[7];
  assign FMcvt_in_vld[0] = fp_lut_pvld_f & (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:16763" *) _3739_;
  assign FMcvt_in_vld[1] = fp_lut_pvld_f & (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:16764" *) _3740_;
  assign FMcvt_in_vld[2] = fp_lut_pvld_f & (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:16765" *) _3741_;
  assign FMcvt_in_vld[3] = fp_lut_pvld_f & (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:16766" *) _3742_;
  assign FMcvt_out_rdy[0] = fp_out_prdy & (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:16863" *) _3743_;
  assign FMcvt_out_rdy[1] = fp_out_prdy & (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:16864" *) _3744_;
  assign FMcvt_out_rdy[2] = fp_out_prdy & (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:16865" *) _3745_;
  assign FMcvt_out_rdy[3] = fp_out_prdy & (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:16866" *) _3746_;
  assign load_din = dp2lut_pvld & (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4557" *) dp2lut_prdy_f;
  assign _0392_ = load_din & (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4950" *) lut_X_sel[0];
  assign _0393_ = load_din & (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5233" *) lut_X_sel[1];
  assign _0394_ = load_din & (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5516" *) lut_X_sel[2];
  assign _0395_ = load_din & (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5799" *) lut_X_sel[3];
  assign _0396_ = _0386_ & (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6082" *) lut_X_sel[4];
  assign _0397_ = _0386_ & (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6365" *) lut_X_sel[5];
  assign _0398_ = _0386_ & (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6648" *) lut_X_sel[6];
  assign _0399_ = _0386_ & (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6931" *) lut_X_sel[7];
  assign _0400_ = load_din & (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7215" *) lut_Y_sel[0];
  assign _0401_ = load_din & (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8266" *) lut_Y_sel[1];
  assign _0402_ = load_din & (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9317" *) lut_Y_sel[2];
  assign _0403_ = | { _0946_, _0945_ };
  assign _0404_ = | { _1998_, _1997_ };
  assign _0405_ = | { _2261_, _2260_ };
  assign _0406_ = | { _2524_, _2523_ };
  assign _0407_ = | { _1209_, _1208_ };
  assign _0408_ = | { _2787_, _2786_ };
  assign _0409_ = | { _2858_, _2857_ };
  assign _0410_ = | { _2929_, _2928_ };
  assign _0411_ = | { _3000_, _2999_ };
  assign _0412_ = | { _0683_, _0682_ };
  assign _0413_ = | { _3071_, _3070_ };
  assign _0414_ = | { _1472_, _1471_ };
  assign _0415_ = | { _3142_, _3141_ };
  assign _0416_ = | { _3213_, _3212_ };
  assign _0417_ = | { _3284_, _3283_ };
  assign _0418_ = | { _1734_, _1735_ };
  assign _0419_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1002" *) 6'b100001;
  assign _0420_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1012" *) 6'b100010;
  assign _0421_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1022" *) 6'b100011;
  assign _0422_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1032" *) 6'b100100;
  assign _0423_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1042" *) 6'b100101;
  assign _0424_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1052" *) 6'b100110;
  assign _0425_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1062" *) 6'b100111;
  assign _0426_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1072" *) 6'b101000;
  assign _0427_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1082" *) 6'b101001;
  assign _0428_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1092" *) 6'b101010;
  assign _0429_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1102" *) 6'b101011;
  assign _0430_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1112" *) 6'b101100;
  assign _0431_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1122" *) 6'b101101;
  assign _0432_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1132" *) 6'b101110;
  assign _0433_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1142" *) 6'b101111;
  assign _0434_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1152" *) 6'b110000;
  assign _0435_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1162" *) 6'b110001;
  assign _0436_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1172" *) 6'b110010;
  assign _0437_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1182" *) 6'b110011;
  assign _0438_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1192" *) 6'b110100;
  assign _0439_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1202" *) 6'b110101;
  assign _0440_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1212" *) 6'b110110;
  assign _0441_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1222" *) 6'b110111;
  assign _0442_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1232" *) 6'b111000;
  assign _0443_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1242" *) 6'b111001;
  assign _0444_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1252" *) 6'b111010;
  assign _0445_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1262" *) 6'b111011;
  assign _0446_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1272" *) 6'b111100;
  assign _0447_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1282" *) 6'b111101;
  assign _0448_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1292" *) 6'b111110;
  assign _0449_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1302" *) 6'b111111;
  assign _0450_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1312" *) 7'b1000000;
  assign _0451_ = ! (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1323" *) reg2dp_lut_addr;
  assign _0452_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1333" *) 1'b1;
  assign _0453_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1343" *) 2'b10;
  assign _0454_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1353" *) 2'b11;
  assign _0455_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1363" *) 3'b100;
  assign _0456_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1373" *) 3'b101;
  assign _0457_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1383" *) 3'b110;
  assign _0458_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1393" *) 3'b111;
  assign _0459_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1403" *) 4'b1000;
  assign _0460_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1413" *) 4'b1001;
  assign _0461_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1423" *) 4'b1010;
  assign _0462_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1433" *) 4'b1011;
  assign _0463_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1443" *) 4'b1100;
  assign _0464_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1453" *) 4'b1101;
  assign _0465_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1463" *) 4'b1110;
  assign _0466_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1473" *) 4'b1111;
  assign _0467_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1483" *) 5'b10000;
  assign _0468_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1493" *) 5'b10001;
  assign _0469_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1503" *) 5'b10010;
  assign _0470_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1513" *) 5'b10011;
  assign _0471_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1523" *) 5'b10100;
  assign _0472_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1533" *) 5'b10101;
  assign _0473_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1543" *) 5'b10110;
  assign _0474_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1553" *) 5'b10111;
  assign _0475_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1563" *) 5'b11000;
  assign _0476_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1573" *) 5'b11001;
  assign _0477_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1583" *) 5'b11010;
  assign _0478_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1593" *) 5'b11011;
  assign _0479_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1603" *) 5'b11100;
  assign _0480_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1613" *) 5'b11101;
  assign _0481_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1623" *) 5'b11110;
  assign _0482_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1633" *) 5'b11111;
  assign _0483_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1643" *) 6'b100000;
  assign _0258_ = reg2dp_input_data_type == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:16754" *) 2'b10;
  assign _0484_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1973" *) 7'b1000001;
  assign _0485_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1983" *) 7'b1000010;
  assign _0486_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1993" *) 7'b1000011;
  assign _0487_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2003" *) 7'b1000100;
  assign _0488_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2013" *) 7'b1000101;
  assign _0489_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2023" *) 7'b1000110;
  assign _0490_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2033" *) 7'b1000111;
  assign _0491_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2043" *) 7'b1001000;
  assign _0492_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2053" *) 7'b1001001;
  assign _0493_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2063" *) 7'b1001010;
  assign _0494_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2073" *) 7'b1001011;
  assign _0495_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2083" *) 7'b1001100;
  assign _0496_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2093" *) 7'b1001101;
  assign _0497_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2103" *) 7'b1001110;
  assign _0498_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2113" *) 7'b1001111;
  assign _0499_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2123" *) 7'b1010000;
  assign _0500_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2133" *) 7'b1010001;
  assign _0501_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2143" *) 7'b1010010;
  assign _0502_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2153" *) 7'b1010011;
  assign _0503_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2163" *) 7'b1010100;
  assign _0504_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2173" *) 7'b1010101;
  assign _0505_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2183" *) 7'b1010110;
  assign _0506_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2193" *) 7'b1010111;
  assign _0507_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2203" *) 7'b1011000;
  assign _0508_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2213" *) 7'b1011001;
  assign _0509_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2223" *) 7'b1011010;
  assign _0510_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2233" *) 7'b1011011;
  assign _0511_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2243" *) 7'b1011100;
  assign _0512_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2253" *) 7'b1011101;
  assign _0513_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2263" *) 7'b1011110;
  assign _0514_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2273" *) 7'b1011111;
  assign _0515_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2283" *) 7'b1100000;
  assign _0516_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2293" *) 7'b1100001;
  assign _0517_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2303" *) 7'b1100010;
  assign _0518_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2313" *) 7'b1100011;
  assign _0519_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2323" *) 7'b1100100;
  assign _0520_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2333" *) 7'b1100101;
  assign _0521_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2343" *) 7'b1100110;
  assign _0522_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2353" *) 7'b1100111;
  assign _0523_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2363" *) 7'b1101000;
  assign _0524_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2373" *) 7'b1101001;
  assign _0525_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2383" *) 7'b1101010;
  assign _0526_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2393" *) 7'b1101011;
  assign _0527_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2403" *) 7'b1101100;
  assign _0528_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2413" *) 7'b1101101;
  assign _0529_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2423" *) 7'b1101110;
  assign _0530_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2433" *) 7'b1101111;
  assign _0531_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2443" *) 7'b1110000;
  assign _0532_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2453" *) 7'b1110001;
  assign _0533_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2463" *) 7'b1110010;
  assign _0534_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2473" *) 7'b1110011;
  assign _0535_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2483" *) 7'b1110100;
  assign _0536_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2493" *) 7'b1110101;
  assign _0537_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2503" *) 7'b1110110;
  assign _0538_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2513" *) 7'b1110111;
  assign _0539_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2523" *) 7'b1111000;
  assign _0540_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2533" *) 7'b1111001;
  assign _0541_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2543" *) 7'b1111010;
  assign _0542_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2553" *) 7'b1111011;
  assign _0543_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2563" *) 7'b1111100;
  assign _0544_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2573" *) 7'b1111101;
  assign _0545_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2583" *) 7'b1111110;
  assign _0546_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2593" *) 7'b1111111;
  assign _0547_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2603" *) 8'b10000000;
  assign _0548_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2613" *) 8'b10000001;
  assign _0549_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2623" *) 8'b10000010;
  assign _0550_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2633" *) 8'b10000011;
  assign _0551_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2643" *) 8'b10000100;
  assign _0552_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2653" *) 8'b10000101;
  assign _0553_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2663" *) 8'b10000110;
  assign _0554_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2673" *) 8'b10000111;
  assign _0555_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2683" *) 8'b10001000;
  assign _0556_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2693" *) 8'b10001001;
  assign _0557_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2703" *) 8'b10001010;
  assign _0558_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2713" *) 8'b10001011;
  assign _0559_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2723" *) 8'b10001100;
  assign _0560_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2733" *) 8'b10001101;
  assign _0561_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2743" *) 8'b10001110;
  assign _0562_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2753" *) 8'b10001111;
  assign _0563_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2763" *) 8'b10010000;
  assign _0564_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2773" *) 8'b10010001;
  assign _0565_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2783" *) 8'b10010010;
  assign _0566_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2793" *) 8'b10010011;
  assign _0567_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2803" *) 8'b10010100;
  assign _0568_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2813" *) 8'b10010101;
  assign _0569_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2823" *) 8'b10010110;
  assign _0570_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2833" *) 8'b10010111;
  assign _0571_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2843" *) 8'b10011000;
  assign _0572_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2853" *) 8'b10011001;
  assign _0573_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2863" *) 8'b10011010;
  assign _0574_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2873" *) 8'b10011011;
  assign _0575_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2883" *) 8'b10011100;
  assign _0576_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2893" *) 8'b10011101;
  assign _0577_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2903" *) 8'b10011110;
  assign _0578_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2913" *) 8'b10011111;
  assign _0579_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2923" *) 8'b10100000;
  assign _0580_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2933" *) 8'b10100001;
  assign _0581_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2943" *) 8'b10100010;
  assign _0582_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2953" *) 8'b10100011;
  assign _0583_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2963" *) 8'b10100100;
  assign _0584_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2973" *) 8'b10100101;
  assign _0585_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2983" *) 8'b10100110;
  assign _0586_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2993" *) 8'b10100111;
  assign _0587_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3003" *) 8'b10101000;
  assign _0588_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3013" *) 8'b10101001;
  assign _0589_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3023" *) 8'b10101010;
  assign _0590_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3033" *) 8'b10101011;
  assign _0591_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3043" *) 8'b10101100;
  assign _0592_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3053" *) 8'b10101101;
  assign _0593_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3063" *) 8'b10101110;
  assign _0594_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3073" *) 8'b10101111;
  assign _0595_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3083" *) 8'b10110000;
  assign _0596_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3093" *) 8'b10110001;
  assign _0597_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3103" *) 8'b10110010;
  assign _0598_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3113" *) 8'b10110011;
  assign _0599_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3123" *) 8'b10110100;
  assign _0600_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3133" *) 8'b10110101;
  assign _0601_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3143" *) 8'b10110110;
  assign _0602_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3153" *) 8'b10110111;
  assign _0603_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3163" *) 8'b10111000;
  assign _0604_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3173" *) 8'b10111001;
  assign _0605_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3183" *) 8'b10111010;
  assign _0606_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3193" *) 8'b10111011;
  assign _0607_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3203" *) 8'b10111100;
  assign _0608_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3213" *) 8'b10111101;
  assign _0609_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3223" *) 8'b10111110;
  assign _0610_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3233" *) 8'b10111111;
  assign _0611_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3243" *) 8'b11000000;
  assign _0612_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3253" *) 8'b11000001;
  assign _0613_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3263" *) 8'b11000010;
  assign _0614_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3273" *) 8'b11000011;
  assign _0615_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3283" *) 8'b11000100;
  assign _0616_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3293" *) 8'b11000101;
  assign _0617_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3303" *) 8'b11000110;
  assign _0618_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3313" *) 8'b11000111;
  assign _0619_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3323" *) 8'b11001000;
  assign _0620_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3333" *) 8'b11001001;
  assign _0621_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3343" *) 8'b11001010;
  assign _0622_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3353" *) 8'b11001011;
  assign _0623_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3363" *) 8'b11001100;
  assign _0624_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3373" *) 8'b11001101;
  assign _0625_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3383" *) 8'b11001110;
  assign _0626_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3393" *) 8'b11001111;
  assign _0627_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3403" *) 8'b11010000;
  assign _0628_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3413" *) 8'b11010001;
  assign _0629_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3423" *) 8'b11010010;
  assign _0630_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3433" *) 8'b11010011;
  assign _0631_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3443" *) 8'b11010100;
  assign _0632_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3453" *) 8'b11010101;
  assign _0633_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3463" *) 8'b11010110;
  assign _0634_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3473" *) 8'b11010111;
  assign _0635_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3483" *) 8'b11011000;
  assign _0636_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3493" *) 8'b11011001;
  assign _0637_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3503" *) 8'b11011010;
  assign _0638_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3513" *) 8'b11011011;
  assign _0639_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3523" *) 8'b11011100;
  assign _0640_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3533" *) 8'b11011101;
  assign _0641_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3543" *) 8'b11011110;
  assign _0642_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3553" *) 8'b11011111;
  assign _0643_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3563" *) 8'b11100000;
  assign _0644_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3573" *) 8'b11100001;
  assign _0645_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3583" *) 8'b11100010;
  assign _0646_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3593" *) 8'b11100011;
  assign _0647_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3603" *) 8'b11100100;
  assign _0648_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3613" *) 8'b11100101;
  assign _0649_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3623" *) 8'b11100110;
  assign _0650_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3633" *) 8'b11100111;
  assign _0651_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3643" *) 8'b11101000;
  assign _0652_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3653" *) 8'b11101001;
  assign _0653_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3663" *) 8'b11101010;
  assign _0654_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3673" *) 8'b11101011;
  assign _0655_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3683" *) 8'b11101100;
  assign _0656_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3693" *) 8'b11101101;
  assign _0657_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3703" *) 8'b11101110;
  assign _0658_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3713" *) 8'b11101111;
  assign _0659_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3723" *) 8'b11110000;
  assign _0660_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3733" *) 8'b11110001;
  assign _0661_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3743" *) 8'b11110010;
  assign _0662_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3753" *) 8'b11110011;
  assign _0663_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3763" *) 8'b11110100;
  assign _0664_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3773" *) 8'b11110101;
  assign _0665_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3783" *) 8'b11110110;
  assign _0666_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3793" *) 8'b11110111;
  assign _0667_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3803" *) 8'b11111000;
  assign _0668_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3813" *) 8'b11111001;
  assign _0669_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3823" *) 8'b11111010;
  assign _0670_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3833" *) 8'b11111011;
  assign _0671_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3843" *) 8'b11111100;
  assign _0672_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3853" *) 8'b11111101;
  assign _0673_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3863" *) 8'b11111110;
  assign _0674_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3873" *) 8'b11111111;
  assign _0675_ = reg2dp_lut_addr == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3883" *) 9'b100000000;
  assign raw_select = ~ (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:663" *) reg2dp_lut_table_id;
  assign lut_wr_en = reg2dp_lut_access_type && (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:662" *) reg2dp_lut_data_trigger;
  assign _0676_ = ~ (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4558" *) lut_pvld_f;
  assign _0677_ = ~ (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4574" *) reg2dp_lut_hybrid_priority;
  assign _0678_ = ~ (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4577" *) reg2dp_lut_uflow_priority;
  assign _0679_ = ~ (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4578" *) reg2dp_lut_oflow_priority;
  assign dp2lut_prdy_f = _0676_ | (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4558" *) lut_prdy;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      fp16_en_f <= 1'b0;
    else
      fp16_en_f <= _0258_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_pvld_f <= 1'b0;
    else
      lut_pvld_f <= _0309_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lutY_sel <= 8'b00000000;
    else
      lutY_sel <= _0260_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_Y_info_7 <= 18'b000000000000000000;
    else
      lut_Y_info_7 <= _0308_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_Y_info_6 <= 18'b000000000000000000;
    else
      lut_Y_info_6 <= _0307_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_Y_info_5 <= 18'b000000000000000000;
    else
      lut_Y_info_5 <= _0306_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_Y_info_4 <= 18'b000000000000000000;
    else
      lut_Y_info_4 <= _0305_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_Y_info_3 <= 18'b000000000000000000;
    else
      lut_Y_info_3 <= _0304_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_Y_info_2 <= 18'b000000000000000000;
    else
      lut_Y_info_2 <= _0303_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_Y_info_1 <= 18'b000000000000000000;
    else
      lut_Y_info_1 <= _0302_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_Y_info_0 <= 18'b000000000000000000;
    else
      lut_Y_info_0 <= _0301_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lutX_sel <= 8'b00000000;
    else
      lutX_sel <= _0259_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_X_info_7 <= 18'b000000000000000000;
    else
      lut_X_info_7 <= _0284_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_X_info_6 <= 18'b000000000000000000;
    else
      lut_X_info_6 <= _0283_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_X_info_5 <= 18'b000000000000000000;
    else
      lut_X_info_5 <= _0282_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_X_info_4 <= 18'b000000000000000000;
    else
      lut_X_info_4 <= _0281_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_X_info_3 <= 18'b000000000000000000;
    else
      lut_X_info_3 <= _0280_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_X_info_2 <= 18'b000000000000000000;
    else
      lut_X_info_2 <= _0279_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_X_info_1 <= 18'b000000000000000000;
    else
      lut_X_info_1 <= _0278_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_X_info_0 <= 18'b000000000000000000;
    else
      lut_X_info_0 <= _0277_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_Y_data_70 <= 16'b0000000000000000;
    else
      lut_Y_data_70 <= _0299_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_Y_data_71 <= 16'b0000000000000000;
    else
      lut_Y_data_71 <= _0300_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_Y_data_60 <= 16'b0000000000000000;
    else
      lut_Y_data_60 <= _0297_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_Y_data_61 <= 16'b0000000000000000;
    else
      lut_Y_data_61 <= _0298_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_Y_data_50 <= 16'b0000000000000000;
    else
      lut_Y_data_50 <= _0295_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_Y_data_51 <= 16'b0000000000000000;
    else
      lut_Y_data_51 <= _0296_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_Y_data_40 <= 16'b0000000000000000;
    else
      lut_Y_data_40 <= _0293_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_Y_data_41 <= 16'b0000000000000000;
    else
      lut_Y_data_41 <= _0294_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_Y_data_30 <= 16'b0000000000000000;
    else
      lut_Y_data_30 <= _0291_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_Y_data_31 <= 16'b0000000000000000;
    else
      lut_Y_data_31 <= _0292_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_Y_data_20 <= 16'b0000000000000000;
    else
      lut_Y_data_20 <= _0289_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_Y_data_21 <= 16'b0000000000000000;
    else
      lut_Y_data_21 <= _0290_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_Y_data_10 <= 16'b0000000000000000;
    else
      lut_Y_data_10 <= _0287_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_Y_data_11 <= 16'b0000000000000000;
    else
      lut_Y_data_11 <= _0288_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_Y_data_00 <= 16'b0000000000000000;
    else
      lut_Y_data_00 <= _0285_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_Y_data_01 <= 16'b0000000000000000;
    else
      lut_Y_data_01 <= _0286_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_X_data_70 <= 16'b0000000000000000;
    else
      lut_X_data_70 <= _0275_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_X_data_71 <= 16'b0000000000000000;
    else
      lut_X_data_71 <= _0276_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_X_data_60 <= 16'b0000000000000000;
    else
      lut_X_data_60 <= _0273_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_X_data_61 <= 16'b0000000000000000;
    else
      lut_X_data_61 <= _0274_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_X_data_50 <= 16'b0000000000000000;
    else
      lut_X_data_50 <= _0271_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_X_data_51 <= 16'b0000000000000000;
    else
      lut_X_data_51 <= _0272_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_X_data_40 <= 16'b0000000000000000;
    else
      lut_X_data_40 <= _0269_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_X_data_41 <= 16'b0000000000000000;
    else
      lut_X_data_41 <= _0270_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_X_data_30 <= 16'b0000000000000000;
    else
      lut_X_data_30 <= _0267_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_X_data_31 <= 16'b0000000000000000;
    else
      lut_X_data_31 <= _0268_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_X_data_20 <= 16'b0000000000000000;
    else
      lut_X_data_20 <= _0265_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_X_data_21 <= 16'b0000000000000000;
    else
      lut_X_data_21 <= _0266_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_X_data_10 <= 16'b0000000000000000;
    else
      lut_X_data_10 <= _0263_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_X_data_11 <= 16'b0000000000000000;
    else
      lut_X_data_11 <= _0264_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_X_data_00 <= 16'b0000000000000000;
    else
      lut_X_data_00 <= _0261_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_X_data_01 <= 16'b0000000000000000;
    else
      lut_X_data_01 <= _0262_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_out <= 16'b0000000000000000;
    else
      density_out <= _0000_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      raw_out <= 16'b0000000000000000;
    else
      raw_out <= _0310_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg256 <= 16'b0000000000000000;
    else
      density_reg256 <= _0174_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg255 <= 16'b0000000000000000;
    else
      density_reg255 <= _0173_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg254 <= 16'b0000000000000000;
    else
      density_reg254 <= _0172_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg253 <= 16'b0000000000000000;
    else
      density_reg253 <= _0171_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg252 <= 16'b0000000000000000;
    else
      density_reg252 <= _0170_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg251 <= 16'b0000000000000000;
    else
      density_reg251 <= _0169_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg250 <= 16'b0000000000000000;
    else
      density_reg250 <= _0168_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg249 <= 16'b0000000000000000;
    else
      density_reg249 <= _0166_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg248 <= 16'b0000000000000000;
    else
      density_reg248 <= _0165_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg247 <= 16'b0000000000000000;
    else
      density_reg247 <= _0164_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg246 <= 16'b0000000000000000;
    else
      density_reg246 <= _0163_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg245 <= 16'b0000000000000000;
    else
      density_reg245 <= _0162_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg244 <= 16'b0000000000000000;
    else
      density_reg244 <= _0161_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg243 <= 16'b0000000000000000;
    else
      density_reg243 <= _0160_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg242 <= 16'b0000000000000000;
    else
      density_reg242 <= _0159_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg241 <= 16'b0000000000000000;
    else
      density_reg241 <= _0158_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg240 <= 16'b0000000000000000;
    else
      density_reg240 <= _0157_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg239 <= 16'b0000000000000000;
    else
      density_reg239 <= _0155_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg238 <= 16'b0000000000000000;
    else
      density_reg238 <= _0154_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg237 <= 16'b0000000000000000;
    else
      density_reg237 <= _0153_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg236 <= 16'b0000000000000000;
    else
      density_reg236 <= _0152_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg235 <= 16'b0000000000000000;
    else
      density_reg235 <= _0151_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg234 <= 16'b0000000000000000;
    else
      density_reg234 <= _0150_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg233 <= 16'b0000000000000000;
    else
      density_reg233 <= _0149_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg232 <= 16'b0000000000000000;
    else
      density_reg232 <= _0148_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg231 <= 16'b0000000000000000;
    else
      density_reg231 <= _0147_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg230 <= 16'b0000000000000000;
    else
      density_reg230 <= _0146_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg229 <= 16'b0000000000000000;
    else
      density_reg229 <= _0144_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg228 <= 16'b0000000000000000;
    else
      density_reg228 <= _0143_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg227 <= 16'b0000000000000000;
    else
      density_reg227 <= _0142_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg226 <= 16'b0000000000000000;
    else
      density_reg226 <= _0141_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg225 <= 16'b0000000000000000;
    else
      density_reg225 <= _0140_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg224 <= 16'b0000000000000000;
    else
      density_reg224 <= _0139_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg223 <= 16'b0000000000000000;
    else
      density_reg223 <= _0138_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg222 <= 16'b0000000000000000;
    else
      density_reg222 <= _0137_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg221 <= 16'b0000000000000000;
    else
      density_reg221 <= _0136_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg220 <= 16'b0000000000000000;
    else
      density_reg220 <= _0135_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg219 <= 16'b0000000000000000;
    else
      density_reg219 <= _0133_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg218 <= 16'b0000000000000000;
    else
      density_reg218 <= _0132_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg217 <= 16'b0000000000000000;
    else
      density_reg217 <= _0131_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg216 <= 16'b0000000000000000;
    else
      density_reg216 <= _0130_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg215 <= 16'b0000000000000000;
    else
      density_reg215 <= _0129_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg214 <= 16'b0000000000000000;
    else
      density_reg214 <= _0128_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg213 <= 16'b0000000000000000;
    else
      density_reg213 <= _0127_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg212 <= 16'b0000000000000000;
    else
      density_reg212 <= _0126_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg211 <= 16'b0000000000000000;
    else
      density_reg211 <= _0125_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg210 <= 16'b0000000000000000;
    else
      density_reg210 <= _0124_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg209 <= 16'b0000000000000000;
    else
      density_reg209 <= _0122_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg208 <= 16'b0000000000000000;
    else
      density_reg208 <= _0121_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg207 <= 16'b0000000000000000;
    else
      density_reg207 <= _0120_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg206 <= 16'b0000000000000000;
    else
      density_reg206 <= _0119_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg205 <= 16'b0000000000000000;
    else
      density_reg205 <= _0118_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg204 <= 16'b0000000000000000;
    else
      density_reg204 <= _0117_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg203 <= 16'b0000000000000000;
    else
      density_reg203 <= _0116_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg202 <= 16'b0000000000000000;
    else
      density_reg202 <= _0115_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg201 <= 16'b0000000000000000;
    else
      density_reg201 <= _0114_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg200 <= 16'b0000000000000000;
    else
      density_reg200 <= _0113_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg199 <= 16'b0000000000000000;
    else
      density_reg199 <= _0110_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg198 <= 16'b0000000000000000;
    else
      density_reg198 <= _0109_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg197 <= 16'b0000000000000000;
    else
      density_reg197 <= _0108_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg196 <= 16'b0000000000000000;
    else
      density_reg196 <= _0107_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg195 <= 16'b0000000000000000;
    else
      density_reg195 <= _0106_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg194 <= 16'b0000000000000000;
    else
      density_reg194 <= _0105_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg193 <= 16'b0000000000000000;
    else
      density_reg193 <= _0104_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg192 <= 16'b0000000000000000;
    else
      density_reg192 <= _0103_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg191 <= 16'b0000000000000000;
    else
      density_reg191 <= _0102_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg190 <= 16'b0000000000000000;
    else
      density_reg190 <= _0101_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg189 <= 16'b0000000000000000;
    else
      density_reg189 <= _0099_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg188 <= 16'b0000000000000000;
    else
      density_reg188 <= _0098_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg187 <= 16'b0000000000000000;
    else
      density_reg187 <= _0097_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg186 <= 16'b0000000000000000;
    else
      density_reg186 <= _0096_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg185 <= 16'b0000000000000000;
    else
      density_reg185 <= _0095_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg184 <= 16'b0000000000000000;
    else
      density_reg184 <= _0094_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg183 <= 16'b0000000000000000;
    else
      density_reg183 <= _0093_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg182 <= 16'b0000000000000000;
    else
      density_reg182 <= _0092_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg181 <= 16'b0000000000000000;
    else
      density_reg181 <= _0091_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg180 <= 16'b0000000000000000;
    else
      density_reg180 <= _0090_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg179 <= 16'b0000000000000000;
    else
      density_reg179 <= _0088_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg178 <= 16'b0000000000000000;
    else
      density_reg178 <= _0087_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg177 <= 16'b0000000000000000;
    else
      density_reg177 <= _0086_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg176 <= 16'b0000000000000000;
    else
      density_reg176 <= _0085_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg175 <= 16'b0000000000000000;
    else
      density_reg175 <= _0084_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg174 <= 16'b0000000000000000;
    else
      density_reg174 <= _0083_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg173 <= 16'b0000000000000000;
    else
      density_reg173 <= _0082_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg172 <= 16'b0000000000000000;
    else
      density_reg172 <= _0081_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg171 <= 16'b0000000000000000;
    else
      density_reg171 <= _0080_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg170 <= 16'b0000000000000000;
    else
      density_reg170 <= _0079_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg169 <= 16'b0000000000000000;
    else
      density_reg169 <= _0077_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg168 <= 16'b0000000000000000;
    else
      density_reg168 <= _0076_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg167 <= 16'b0000000000000000;
    else
      density_reg167 <= _0075_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg166 <= 16'b0000000000000000;
    else
      density_reg166 <= _0074_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg165 <= 16'b0000000000000000;
    else
      density_reg165 <= _0073_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg164 <= 16'b0000000000000000;
    else
      density_reg164 <= _0072_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg163 <= 16'b0000000000000000;
    else
      density_reg163 <= _0071_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg162 <= 16'b0000000000000000;
    else
      density_reg162 <= _0070_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg161 <= 16'b0000000000000000;
    else
      density_reg161 <= _0069_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg160 <= 16'b0000000000000000;
    else
      density_reg160 <= _0068_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg159 <= 16'b0000000000000000;
    else
      density_reg159 <= _0066_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg158 <= 16'b0000000000000000;
    else
      density_reg158 <= _0065_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg157 <= 16'b0000000000000000;
    else
      density_reg157 <= _0064_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg156 <= 16'b0000000000000000;
    else
      density_reg156 <= _0063_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg155 <= 16'b0000000000000000;
    else
      density_reg155 <= _0062_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg154 <= 16'b0000000000000000;
    else
      density_reg154 <= _0061_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg153 <= 16'b0000000000000000;
    else
      density_reg153 <= _0060_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg152 <= 16'b0000000000000000;
    else
      density_reg152 <= _0059_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg151 <= 16'b0000000000000000;
    else
      density_reg151 <= _0058_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg150 <= 16'b0000000000000000;
    else
      density_reg150 <= _0057_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg149 <= 16'b0000000000000000;
    else
      density_reg149 <= _0055_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg148 <= 16'b0000000000000000;
    else
      density_reg148 <= _0054_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg147 <= 16'b0000000000000000;
    else
      density_reg147 <= _0053_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg146 <= 16'b0000000000000000;
    else
      density_reg146 <= _0052_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg145 <= 16'b0000000000000000;
    else
      density_reg145 <= _0051_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg144 <= 16'b0000000000000000;
    else
      density_reg144 <= _0050_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg143 <= 16'b0000000000000000;
    else
      density_reg143 <= _0049_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg142 <= 16'b0000000000000000;
    else
      density_reg142 <= _0048_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg141 <= 16'b0000000000000000;
    else
      density_reg141 <= _0047_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg140 <= 16'b0000000000000000;
    else
      density_reg140 <= _0046_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg139 <= 16'b0000000000000000;
    else
      density_reg139 <= _0044_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg138 <= 16'b0000000000000000;
    else
      density_reg138 <= _0043_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg137 <= 16'b0000000000000000;
    else
      density_reg137 <= _0042_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg136 <= 16'b0000000000000000;
    else
      density_reg136 <= _0041_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg135 <= 16'b0000000000000000;
    else
      density_reg135 <= _0040_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg134 <= 16'b0000000000000000;
    else
      density_reg134 <= _0039_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg133 <= 16'b0000000000000000;
    else
      density_reg133 <= _0038_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg132 <= 16'b0000000000000000;
    else
      density_reg132 <= _0037_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg131 <= 16'b0000000000000000;
    else
      density_reg131 <= _0036_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg130 <= 16'b0000000000000000;
    else
      density_reg130 <= _0035_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg129 <= 16'b0000000000000000;
    else
      density_reg129 <= _0033_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg128 <= 16'b0000000000000000;
    else
      density_reg128 <= _0032_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg127 <= 16'b0000000000000000;
    else
      density_reg127 <= _0031_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg126 <= 16'b0000000000000000;
    else
      density_reg126 <= _0030_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg125 <= 16'b0000000000000000;
    else
      density_reg125 <= _0029_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg124 <= 16'b0000000000000000;
    else
      density_reg124 <= _0028_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg123 <= 16'b0000000000000000;
    else
      density_reg123 <= _0027_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg122 <= 16'b0000000000000000;
    else
      density_reg122 <= _0026_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg121 <= 16'b0000000000000000;
    else
      density_reg121 <= _0025_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg120 <= 16'b0000000000000000;
    else
      density_reg120 <= _0024_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg119 <= 16'b0000000000000000;
    else
      density_reg119 <= _0022_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg118 <= 16'b0000000000000000;
    else
      density_reg118 <= _0021_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg117 <= 16'b0000000000000000;
    else
      density_reg117 <= _0020_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg116 <= 16'b0000000000000000;
    else
      density_reg116 <= _0019_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg115 <= 16'b0000000000000000;
    else
      density_reg115 <= _0018_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg114 <= 16'b0000000000000000;
    else
      density_reg114 <= _0017_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg113 <= 16'b0000000000000000;
    else
      density_reg113 <= _0016_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg112 <= 16'b0000000000000000;
    else
      density_reg112 <= _0015_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg111 <= 16'b0000000000000000;
    else
      density_reg111 <= _0014_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg110 <= 16'b0000000000000000;
    else
      density_reg110 <= _0013_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg109 <= 16'b0000000000000000;
    else
      density_reg109 <= _0011_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg108 <= 16'b0000000000000000;
    else
      density_reg108 <= _0010_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg107 <= 16'b0000000000000000;
    else
      density_reg107 <= _0009_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg106 <= 16'b0000000000000000;
    else
      density_reg106 <= _0008_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg105 <= 16'b0000000000000000;
    else
      density_reg105 <= _0007_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg104 <= 16'b0000000000000000;
    else
      density_reg104 <= _0006_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg103 <= 16'b0000000000000000;
    else
      density_reg103 <= _0005_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg102 <= 16'b0000000000000000;
    else
      density_reg102 <= _0004_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg101 <= 16'b0000000000000000;
    else
      density_reg101 <= _0003_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg100 <= 16'b0000000000000000;
    else
      density_reg100 <= _0002_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg99 <= 16'b0000000000000000;
    else
      density_reg99 <= _0256_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg98 <= 16'b0000000000000000;
    else
      density_reg98 <= _0255_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg97 <= 16'b0000000000000000;
    else
      density_reg97 <= _0254_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg96 <= 16'b0000000000000000;
    else
      density_reg96 <= _0253_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg95 <= 16'b0000000000000000;
    else
      density_reg95 <= _0252_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg94 <= 16'b0000000000000000;
    else
      density_reg94 <= _0251_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg93 <= 16'b0000000000000000;
    else
      density_reg93 <= _0250_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg92 <= 16'b0000000000000000;
    else
      density_reg92 <= _0249_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg91 <= 16'b0000000000000000;
    else
      density_reg91 <= _0248_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg90 <= 16'b0000000000000000;
    else
      density_reg90 <= _0247_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg89 <= 16'b0000000000000000;
    else
      density_reg89 <= _0245_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg88 <= 16'b0000000000000000;
    else
      density_reg88 <= _0244_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg87 <= 16'b0000000000000000;
    else
      density_reg87 <= _0243_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg86 <= 16'b0000000000000000;
    else
      density_reg86 <= _0242_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg85 <= 16'b0000000000000000;
    else
      density_reg85 <= _0241_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg84 <= 16'b0000000000000000;
    else
      density_reg84 <= _0240_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg83 <= 16'b0000000000000000;
    else
      density_reg83 <= _0239_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg82 <= 16'b0000000000000000;
    else
      density_reg82 <= _0238_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg81 <= 16'b0000000000000000;
    else
      density_reg81 <= _0237_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg80 <= 16'b0000000000000000;
    else
      density_reg80 <= _0236_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg79 <= 16'b0000000000000000;
    else
      density_reg79 <= _0234_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg78 <= 16'b0000000000000000;
    else
      density_reg78 <= _0233_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg77 <= 16'b0000000000000000;
    else
      density_reg77 <= _0232_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg76 <= 16'b0000000000000000;
    else
      density_reg76 <= _0231_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg75 <= 16'b0000000000000000;
    else
      density_reg75 <= _0230_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg74 <= 16'b0000000000000000;
    else
      density_reg74 <= _0229_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg73 <= 16'b0000000000000000;
    else
      density_reg73 <= _0228_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg72 <= 16'b0000000000000000;
    else
      density_reg72 <= _0227_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg71 <= 16'b0000000000000000;
    else
      density_reg71 <= _0226_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg70 <= 16'b0000000000000000;
    else
      density_reg70 <= _0225_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg69 <= 16'b0000000000000000;
    else
      density_reg69 <= _0223_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg68 <= 16'b0000000000000000;
    else
      density_reg68 <= _0222_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg67 <= 16'b0000000000000000;
    else
      density_reg67 <= _0221_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg66 <= 16'b0000000000000000;
    else
      density_reg66 <= _0220_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg65 <= 16'b0000000000000000;
    else
      density_reg65 <= _0219_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg64 <= 16'b0000000000000000;
    else
      density_reg64 <= _0218_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg63 <= 16'b0000000000000000;
    else
      density_reg63 <= _0217_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg62 <= 16'b0000000000000000;
    else
      density_reg62 <= _0216_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg61 <= 16'b0000000000000000;
    else
      density_reg61 <= _0215_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg60 <= 16'b0000000000000000;
    else
      density_reg60 <= _0214_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg59 <= 16'b0000000000000000;
    else
      density_reg59 <= _0212_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg58 <= 16'b0000000000000000;
    else
      density_reg58 <= _0211_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg57 <= 16'b0000000000000000;
    else
      density_reg57 <= _0210_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg56 <= 16'b0000000000000000;
    else
      density_reg56 <= _0209_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg55 <= 16'b0000000000000000;
    else
      density_reg55 <= _0208_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg54 <= 16'b0000000000000000;
    else
      density_reg54 <= _0207_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg53 <= 16'b0000000000000000;
    else
      density_reg53 <= _0206_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg52 <= 16'b0000000000000000;
    else
      density_reg52 <= _0205_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg51 <= 16'b0000000000000000;
    else
      density_reg51 <= _0204_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg50 <= 16'b0000000000000000;
    else
      density_reg50 <= _0203_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg49 <= 16'b0000000000000000;
    else
      density_reg49 <= _0201_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg48 <= 16'b0000000000000000;
    else
      density_reg48 <= _0200_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg47 <= 16'b0000000000000000;
    else
      density_reg47 <= _0199_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg46 <= 16'b0000000000000000;
    else
      density_reg46 <= _0198_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg45 <= 16'b0000000000000000;
    else
      density_reg45 <= _0197_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg44 <= 16'b0000000000000000;
    else
      density_reg44 <= _0196_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg43 <= 16'b0000000000000000;
    else
      density_reg43 <= _0195_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg42 <= 16'b0000000000000000;
    else
      density_reg42 <= _0194_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg41 <= 16'b0000000000000000;
    else
      density_reg41 <= _0193_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg40 <= 16'b0000000000000000;
    else
      density_reg40 <= _0192_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg39 <= 16'b0000000000000000;
    else
      density_reg39 <= _0190_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg38 <= 16'b0000000000000000;
    else
      density_reg38 <= _0189_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg37 <= 16'b0000000000000000;
    else
      density_reg37 <= _0188_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg36 <= 16'b0000000000000000;
    else
      density_reg36 <= _0187_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg35 <= 16'b0000000000000000;
    else
      density_reg35 <= _0186_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg34 <= 16'b0000000000000000;
    else
      density_reg34 <= _0185_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg33 <= 16'b0000000000000000;
    else
      density_reg33 <= _0184_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg32 <= 16'b0000000000000000;
    else
      density_reg32 <= _0183_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg31 <= 16'b0000000000000000;
    else
      density_reg31 <= _0182_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg30 <= 16'b0000000000000000;
    else
      density_reg30 <= _0181_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg29 <= 16'b0000000000000000;
    else
      density_reg29 <= _0179_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg28 <= 16'b0000000000000000;
    else
      density_reg28 <= _0178_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg27 <= 16'b0000000000000000;
    else
      density_reg27 <= _0177_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg26 <= 16'b0000000000000000;
    else
      density_reg26 <= _0176_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg25 <= 16'b0000000000000000;
    else
      density_reg25 <= _0175_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg24 <= 16'b0000000000000000;
    else
      density_reg24 <= _0167_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg23 <= 16'b0000000000000000;
    else
      density_reg23 <= _0156_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg22 <= 16'b0000000000000000;
    else
      density_reg22 <= _0145_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg21 <= 16'b0000000000000000;
    else
      density_reg21 <= _0134_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg20 <= 16'b0000000000000000;
    else
      density_reg20 <= _0123_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg19 <= 16'b0000000000000000;
    else
      density_reg19 <= _0111_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg18 <= 16'b0000000000000000;
    else
      density_reg18 <= _0100_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg17 <= 16'b0000000000000000;
    else
      density_reg17 <= _0089_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg16 <= 16'b0000000000000000;
    else
      density_reg16 <= _0078_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg15 <= 16'b0000000000000000;
    else
      density_reg15 <= _0067_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg14 <= 16'b0000000000000000;
    else
      density_reg14 <= _0056_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg13 <= 16'b0000000000000000;
    else
      density_reg13 <= _0045_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg12 <= 16'b0000000000000000;
    else
      density_reg12 <= _0034_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg11 <= 16'b0000000000000000;
    else
      density_reg11 <= _0023_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg10 <= 16'b0000000000000000;
    else
      density_reg10 <= _0012_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg9 <= 16'b0000000000000000;
    else
      density_reg9 <= _0257_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg8 <= 16'b0000000000000000;
    else
      density_reg8 <= _0246_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg7 <= 16'b0000000000000000;
    else
      density_reg7 <= _0235_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg6 <= 16'b0000000000000000;
    else
      density_reg6 <= _0224_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg5 <= 16'b0000000000000000;
    else
      density_reg5 <= _0213_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg4 <= 16'b0000000000000000;
    else
      density_reg4 <= _0202_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg3 <= 16'b0000000000000000;
    else
      density_reg3 <= _0191_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg2 <= 16'b0000000000000000;
    else
      density_reg2 <= _0180_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg1 <= 16'b0000000000000000;
    else
      density_reg1 <= _0112_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      density_reg0 <= 16'b0000000000000000;
    else
      density_reg0 <= _0001_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      raw_reg64 <= 16'b0000000000000000;
    else
      raw_reg64 <= _0371_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      raw_reg63 <= 16'b0000000000000000;
    else
      raw_reg63 <= _0370_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      raw_reg62 <= 16'b0000000000000000;
    else
      raw_reg62 <= _0369_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      raw_reg61 <= 16'b0000000000000000;
    else
      raw_reg61 <= _0368_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      raw_reg60 <= 16'b0000000000000000;
    else
      raw_reg60 <= _0367_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      raw_reg59 <= 16'b0000000000000000;
    else
      raw_reg59 <= _0365_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      raw_reg58 <= 16'b0000000000000000;
    else
      raw_reg58 <= _0364_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      raw_reg57 <= 16'b0000000000000000;
    else
      raw_reg57 <= _0363_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      raw_reg56 <= 16'b0000000000000000;
    else
      raw_reg56 <= _0362_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      raw_reg55 <= 16'b0000000000000000;
    else
      raw_reg55 <= _0361_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      raw_reg54 <= 16'b0000000000000000;
    else
      raw_reg54 <= _0360_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      raw_reg53 <= 16'b0000000000000000;
    else
      raw_reg53 <= _0359_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      raw_reg52 <= 16'b0000000000000000;
    else
      raw_reg52 <= _0358_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      raw_reg51 <= 16'b0000000000000000;
    else
      raw_reg51 <= _0357_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      raw_reg50 <= 16'b0000000000000000;
    else
      raw_reg50 <= _0356_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      raw_reg49 <= 16'b0000000000000000;
    else
      raw_reg49 <= _0354_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      raw_reg48 <= 16'b0000000000000000;
    else
      raw_reg48 <= _0353_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      raw_reg47 <= 16'b0000000000000000;
    else
      raw_reg47 <= _0352_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      raw_reg46 <= 16'b0000000000000000;
    else
      raw_reg46 <= _0351_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      raw_reg45 <= 16'b0000000000000000;
    else
      raw_reg45 <= _0350_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      raw_reg44 <= 16'b0000000000000000;
    else
      raw_reg44 <= _0349_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      raw_reg43 <= 16'b0000000000000000;
    else
      raw_reg43 <= _0348_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      raw_reg42 <= 16'b0000000000000000;
    else
      raw_reg42 <= _0347_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      raw_reg41 <= 16'b0000000000000000;
    else
      raw_reg41 <= _0346_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      raw_reg40 <= 16'b0000000000000000;
    else
      raw_reg40 <= _0345_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      raw_reg39 <= 16'b0000000000000000;
    else
      raw_reg39 <= _0343_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      raw_reg38 <= 16'b0000000000000000;
    else
      raw_reg38 <= _0342_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      raw_reg37 <= 16'b0000000000000000;
    else
      raw_reg37 <= _0341_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      raw_reg36 <= 16'b0000000000000000;
    else
      raw_reg36 <= _0340_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      raw_reg35 <= 16'b0000000000000000;
    else
      raw_reg35 <= _0339_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      raw_reg34 <= 16'b0000000000000000;
    else
      raw_reg34 <= _0338_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      raw_reg33 <= 16'b0000000000000000;
    else
      raw_reg33 <= _0337_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      raw_reg32 <= 16'b0000000000000000;
    else
      raw_reg32 <= _0336_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      raw_reg31 <= 16'b0000000000000000;
    else
      raw_reg31 <= _0335_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      raw_reg30 <= 16'b0000000000000000;
    else
      raw_reg30 <= _0334_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      raw_reg29 <= 16'b0000000000000000;
    else
      raw_reg29 <= _0332_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      raw_reg28 <= 16'b0000000000000000;
    else
      raw_reg28 <= _0331_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      raw_reg27 <= 16'b0000000000000000;
    else
      raw_reg27 <= _0330_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      raw_reg26 <= 16'b0000000000000000;
    else
      raw_reg26 <= _0329_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      raw_reg25 <= 16'b0000000000000000;
    else
      raw_reg25 <= _0328_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      raw_reg24 <= 16'b0000000000000000;
    else
      raw_reg24 <= _0327_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      raw_reg23 <= 16'b0000000000000000;
    else
      raw_reg23 <= _0326_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      raw_reg22 <= 16'b0000000000000000;
    else
      raw_reg22 <= _0325_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      raw_reg21 <= 16'b0000000000000000;
    else
      raw_reg21 <= _0324_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      raw_reg20 <= 16'b0000000000000000;
    else
      raw_reg20 <= _0323_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      raw_reg19 <= 16'b0000000000000000;
    else
      raw_reg19 <= _0321_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      raw_reg18 <= 16'b0000000000000000;
    else
      raw_reg18 <= _0320_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      raw_reg17 <= 16'b0000000000000000;
    else
      raw_reg17 <= _0319_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      raw_reg16 <= 16'b0000000000000000;
    else
      raw_reg16 <= _0318_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      raw_reg15 <= 16'b0000000000000000;
    else
      raw_reg15 <= _0317_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      raw_reg14 <= 16'b0000000000000000;
    else
      raw_reg14 <= _0316_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      raw_reg13 <= 16'b0000000000000000;
    else
      raw_reg13 <= _0315_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      raw_reg12 <= 16'b0000000000000000;
    else
      raw_reg12 <= _0314_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      raw_reg11 <= 16'b0000000000000000;
    else
      raw_reg11 <= _0313_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      raw_reg10 <= 16'b0000000000000000;
    else
      raw_reg10 <= _0312_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      raw_reg9 <= 16'b0000000000000000;
    else
      raw_reg9 <= _0375_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      raw_reg8 <= 16'b0000000000000000;
    else
      raw_reg8 <= _0374_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      raw_reg7 <= 16'b0000000000000000;
    else
      raw_reg7 <= _0373_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      raw_reg6 <= 16'b0000000000000000;
    else
      raw_reg6 <= _0372_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      raw_reg5 <= 16'b0000000000000000;
    else
      raw_reg5 <= _0366_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      raw_reg4 <= 16'b0000000000000000;
    else
      raw_reg4 <= _0355_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      raw_reg3 <= 16'b0000000000000000;
    else
      raw_reg3 <= _0344_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      raw_reg2 <= 16'b0000000000000000;
    else
      raw_reg2 <= _0333_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      raw_reg1 <= 16'b0000000000000000;
    else
      raw_reg1 <= _0322_;
  always @(posedge nvdla_core_clk_orig or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      raw_reg0 <= 16'b0000000000000000;
    else
      raw_reg0 <= _0311_;
  assign lut2intp_Y_sel[7] = fp16_en_f ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:16993" *) 1'b0 : lutY_sel[7];
  assign lut2intp_X_sel[7] = fp16_en_f ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:16993" *) 1'b0 : lutX_sel[7];
  assign lut2intp_X_info_7 = fp16_en_f ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:16993" *) 20'b00000000000000000000 : { lut_Y_info_7[17:16], lut_X_info_7[17:16], lutX_info_7 };
  assign lut2intp_X_data_70_17b = fp16_en_f ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:16993" *) 17'b00000000000000000 : { lutX_data_70[15], lutX_data_70 };
  assign lut2intp_X_data_71 = fp16_en_f ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:16993" *) 32'd0 : { lutX_data_71[15], lutX_data_71[15], lutX_data_71[15], lutX_data_71[15], lutX_data_71[15], lutX_data_71[15], lutX_data_71[15], lutX_data_71[15], lutX_data_71[15], lutX_data_71[15], lutX_data_71[15], lutX_data_71[15], lutX_data_71[15], lutX_data_71[15], lutX_data_71[15], lutX_data_71[15], lutX_data_71 };
  assign lut2intp_X_data_70 = fp16_en_f ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:16993" *) 32'd0 : { lutX_data_70[15], lutX_data_70[15], lutX_data_70[15], lutX_data_70[15], lutX_data_70[15], lutX_data_70[15], lutX_data_70[15], lutX_data_70[15], lutX_data_70[15], lutX_data_70[15], lutX_data_70[15], lutX_data_70[15], lutX_data_70[15], lutX_data_70[15], lutX_data_70[15], lutX_data_70[15], lutX_data_70 };
  assign lut2intp_Y_sel[6] = fp16_en_f ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:16993" *) 1'b0 : lutY_sel[6];
  assign lut2intp_X_sel[6] = fp16_en_f ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:16993" *) 1'b0 : lutX_sel[6];
  assign lut2intp_X_info_6 = fp16_en_f ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:16993" *) 20'b00000000000000000000 : { lut_Y_info_6[17:16], lut_X_info_6[17:16], lutX_info_6 };
  assign lut2intp_X_data_60_17b = fp16_en_f ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:16993" *) 17'b00000000000000000 : { lutX_data_60[15], lutX_data_60 };
  assign lut2intp_X_data_61 = fp16_en_f ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:16993" *) 32'd0 : { lutX_data_61[15], lutX_data_61[15], lutX_data_61[15], lutX_data_61[15], lutX_data_61[15], lutX_data_61[15], lutX_data_61[15], lutX_data_61[15], lutX_data_61[15], lutX_data_61[15], lutX_data_61[15], lutX_data_61[15], lutX_data_61[15], lutX_data_61[15], lutX_data_61[15], lutX_data_61[15], lutX_data_61 };
  assign lut2intp_X_data_60 = fp16_en_f ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:16993" *) 32'd0 : { lutX_data_60[15], lutX_data_60[15], lutX_data_60[15], lutX_data_60[15], lutX_data_60[15], lutX_data_60[15], lutX_data_60[15], lutX_data_60[15], lutX_data_60[15], lutX_data_60[15], lutX_data_60[15], lutX_data_60[15], lutX_data_60[15], lutX_data_60[15], lutX_data_60[15], lutX_data_60[15], lutX_data_60 };
  assign lut2intp_Y_sel[5] = fp16_en_f ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:16993" *) 1'b0 : lutY_sel[5];
  assign lut2intp_X_sel[5] = fp16_en_f ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:16993" *) 1'b0 : lutX_sel[5];
  assign lut2intp_X_info_5 = fp16_en_f ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:16993" *) 20'b00000000000000000000 : { lut_Y_info_5[17:16], lut_X_info_5[17:16], lutX_info_5 };
  assign lut2intp_X_data_50_17b = fp16_en_f ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:16993" *) 17'b00000000000000000 : { lutX_data_50[15], lutX_data_50 };
  assign lut2intp_X_data_51 = fp16_en_f ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:16993" *) 32'd0 : { lutX_data_51[15], lutX_data_51[15], lutX_data_51[15], lutX_data_51[15], lutX_data_51[15], lutX_data_51[15], lutX_data_51[15], lutX_data_51[15], lutX_data_51[15], lutX_data_51[15], lutX_data_51[15], lutX_data_51[15], lutX_data_51[15], lutX_data_51[15], lutX_data_51[15], lutX_data_51[15], lutX_data_51 };
  assign lut2intp_X_data_50 = fp16_en_f ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:16993" *) 32'd0 : { lutX_data_50[15], lutX_data_50[15], lutX_data_50[15], lutX_data_50[15], lutX_data_50[15], lutX_data_50[15], lutX_data_50[15], lutX_data_50[15], lutX_data_50[15], lutX_data_50[15], lutX_data_50[15], lutX_data_50[15], lutX_data_50[15], lutX_data_50[15], lutX_data_50[15], lutX_data_50[15], lutX_data_50 };
  assign lut2intp_Y_sel[4] = fp16_en_f ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:16993" *) 1'b0 : lutY_sel[4];
  assign lut2intp_X_sel[4] = fp16_en_f ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:16993" *) 1'b0 : lutX_sel[4];
  assign lut2intp_X_info_4 = fp16_en_f ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:16993" *) 20'b00000000000000000000 : { lut_Y_info_4[17:16], lut_X_info_4[17:16], lutX_info_4 };
  assign lut2intp_X_data_40_17b = fp16_en_f ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:16993" *) 17'b00000000000000000 : { lutX_data_40[15], lutX_data_40 };
  assign lut2intp_X_data_41 = fp16_en_f ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:16993" *) 32'd0 : { lutX_data_41[15], lutX_data_41[15], lutX_data_41[15], lutX_data_41[15], lutX_data_41[15], lutX_data_41[15], lutX_data_41[15], lutX_data_41[15], lutX_data_41[15], lutX_data_41[15], lutX_data_41[15], lutX_data_41[15], lutX_data_41[15], lutX_data_41[15], lutX_data_41[15], lutX_data_41[15], lutX_data_41 };
  assign lut2intp_X_data_40 = fp16_en_f ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:16993" *) 32'd0 : { lutX_data_40[15], lutX_data_40[15], lutX_data_40[15], lutX_data_40[15], lutX_data_40[15], lutX_data_40[15], lutX_data_40[15], lutX_data_40[15], lutX_data_40[15], lutX_data_40[15], lutX_data_40[15], lutX_data_40[15], lutX_data_40[15], lutX_data_40[15], lutX_data_40[15], lutX_data_40[15], lutX_data_40 };
  assign lut2intp_Y_sel[3] = fp16_en_f ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:16916" *) lutY_sel_o[3] : lutY_sel[3];
  assign lut2intp_X_sel[3] = fp16_en_f ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:16916" *) lutX_sel_o[3] : lutX_sel[3];
  assign lut2intp_X_info_3 = fp16_en_f ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:16916" *) { lut_X_inf_3[20:17], lut_X_inf_3[15:0] } : { lut_Y_info_3[17:16], lut_X_info_3[17:16], lutX_info_3 };
  assign lut2intp_X_data_30_17b = fp16_en_f ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:16916" *) lut_X_dat_30_fp17 : { lutX_data_30[15], lutX_data_30 };
  assign lut2intp_X_data_31 = fp16_en_f ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:16916" *) lut_X_dat_31 : { lutX_data_31[15], lutX_data_31[15], lutX_data_31[15], lutX_data_31[15], lutX_data_31[15], lutX_data_31[15], lutX_data_31[15], lutX_data_31[15], lutX_data_31[15], lutX_data_31[15], lutX_data_31[15], lutX_data_31[15], lutX_data_31[15], lutX_data_31[15], lutX_data_31[15], lutX_data_31[15], lutX_data_31 };
  assign lut2intp_X_data_30 = fp16_en_f ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:16916" *) lut_X_dat_30 : { lutX_data_30[15], lutX_data_30[15], lutX_data_30[15], lutX_data_30[15], lutX_data_30[15], lutX_data_30[15], lutX_data_30[15], lutX_data_30[15], lutX_data_30[15], lutX_data_30[15], lutX_data_30[15], lutX_data_30[15], lutX_data_30[15], lutX_data_30[15], lutX_data_30[15], lutX_data_30[15], lutX_data_30 };
  assign lut2intp_Y_sel[2] = fp16_en_f ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:16916" *) lutY_sel_o[2] : lutY_sel[2];
  assign lut2intp_X_sel[2] = fp16_en_f ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:16916" *) lutX_sel_o[2] : lutX_sel[2];
  assign lut2intp_X_info_2 = fp16_en_f ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:16916" *) { lut_X_inf_2[20:17], lut_X_inf_2[15:0] } : { lut_Y_info_2[17:16], lut_X_info_2[17:16], lutX_info_2 };
  assign lut2intp_X_data_20_17b = fp16_en_f ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:16916" *) lut_X_dat_20_fp17 : { lutX_data_20[15], lutX_data_20 };
  assign lut2intp_X_data_21 = fp16_en_f ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:16916" *) lut_X_dat_21 : { lutX_data_21[15], lutX_data_21[15], lutX_data_21[15], lutX_data_21[15], lutX_data_21[15], lutX_data_21[15], lutX_data_21[15], lutX_data_21[15], lutX_data_21[15], lutX_data_21[15], lutX_data_21[15], lutX_data_21[15], lutX_data_21[15], lutX_data_21[15], lutX_data_21[15], lutX_data_21[15], lutX_data_21 };
  assign lut2intp_X_data_20 = fp16_en_f ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:16916" *) lut_X_dat_20 : { lutX_data_20[15], lutX_data_20[15], lutX_data_20[15], lutX_data_20[15], lutX_data_20[15], lutX_data_20[15], lutX_data_20[15], lutX_data_20[15], lutX_data_20[15], lutX_data_20[15], lutX_data_20[15], lutX_data_20[15], lutX_data_20[15], lutX_data_20[15], lutX_data_20[15], lutX_data_20[15], lutX_data_20 };
  assign lut2intp_Y_sel[1] = fp16_en_f ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:16916" *) lutY_sel_o[1] : lutY_sel[1];
  assign lut2intp_X_sel[1] = fp16_en_f ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:16916" *) lutX_sel_o[1] : lutX_sel[1];
  assign lut2intp_X_info_1 = fp16_en_f ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:16916" *) { lut_X_inf_1[20:17], lut_X_inf_1[15:0] } : { lut_Y_info_1[17:16], lut_X_info_1[17:16], lutX_info_1 };
  assign lut2intp_X_data_10_17b = fp16_en_f ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:16916" *) lut_X_dat_10_fp17 : { lutX_data_10[15], lutX_data_10 };
  assign lut2intp_X_data_11 = fp16_en_f ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:16916" *) lut_X_dat_11 : { lutX_data_11[15], lutX_data_11[15], lutX_data_11[15], lutX_data_11[15], lutX_data_11[15], lutX_data_11[15], lutX_data_11[15], lutX_data_11[15], lutX_data_11[15], lutX_data_11[15], lutX_data_11[15], lutX_data_11[15], lutX_data_11[15], lutX_data_11[15], lutX_data_11[15], lutX_data_11[15], lutX_data_11 };
  assign lut2intp_X_data_10 = fp16_en_f ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:16916" *) lut_X_dat_10 : { lutX_data_10[15], lutX_data_10[15], lutX_data_10[15], lutX_data_10[15], lutX_data_10[15], lutX_data_10[15], lutX_data_10[15], lutX_data_10[15], lutX_data_10[15], lutX_data_10[15], lutX_data_10[15], lutX_data_10[15], lutX_data_10[15], lutX_data_10[15], lutX_data_10[15], lutX_data_10[15], lutX_data_10 };
  assign lut2intp_Y_sel[0] = fp16_en_f ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:16916" *) lutY_sel_o[0] : lutY_sel[0];
  assign lut2intp_X_sel[0] = fp16_en_f ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:16916" *) lutX_sel_o[0] : lutX_sel[0];
  assign lut2intp_X_info_0 = fp16_en_f ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:16916" *) { lut_X_inf_0[20:17], lut_X_inf_0[15:0] } : { lut_Y_info_0[17:16], lut_X_info_0[17:16], lutX_info_0 };
  assign lut2intp_X_data_00_17b = fp16_en_f ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:16916" *) lut_X_dat_00_fp17 : { lutX_data_00[15], lutX_data_00 };
  assign lut2intp_X_data_01 = fp16_en_f ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:16916" *) lut_X_dat_01 : { lutX_data_01[15], lutX_data_01[15], lutX_data_01[15], lutX_data_01[15], lutX_data_01[15], lutX_data_01[15], lutX_data_01[15], lutX_data_01[15], lutX_data_01[15], lutX_data_01[15], lutX_data_01[15], lutX_data_01[15], lutX_data_01[15], lutX_data_01[15], lutX_data_01[15], lutX_data_01[15], lutX_data_01 };
  assign lut2intp_X_data_00 = fp16_en_f ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:16916" *) lut_X_dat_00 : { lutX_data_00[15], lutX_data_00[15], lutX_data_00[15], lutX_data_00[15], lutX_data_00[15], lutX_data_00[15], lutX_data_00[15], lutX_data_00[15], lutX_data_00[15], lutX_data_00[15], lutX_data_00[15], lutX_data_00[15], lutX_data_00[15], lutX_data_00[15], lutX_data_00[15], lutX_data_00[15], lutX_data_00 };
  assign _0680_ = lut_prdy ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:16746" *) 1'b0 : lut_pvld_f;
  assign _0309_ = dp2lut_pvld ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:16744" *) 1'b1 : _0680_;
  assign _0260_ = load_din ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:16659" *) lut_Y_sel : lutY_sel;
  assign _0308_ = _0386_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:16598" *) dp2lut_Yinfo_7 : lut_Y_info_7;
  assign _0307_ = _0386_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:16537" *) dp2lut_Yinfo_6 : lut_Y_info_6;
  assign _0306_ = _0386_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:16476" *) dp2lut_Yinfo_5 : lut_Y_info_5;
  assign _0305_ = _0386_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:16415" *) dp2lut_Yinfo_4 : lut_Y_info_4;
  assign _0304_ = load_din ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:16354" *) dp2lut_Yinfo_3 : lut_Y_info_3;
  assign _0303_ = load_din ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:16293" *) dp2lut_Yinfo_2 : lut_Y_info_2;
  assign _0302_ = load_din ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:16232" *) dp2lut_Yinfo_1 : lut_Y_info_1;
  assign _0301_ = load_din ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:16171" *) dp2lut_Yinfo_0 : lut_Y_info_0;
  assign _0259_ = load_din ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:16110" *) lut_X_sel : lutX_sel;
  assign _0284_ = _0386_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:16049" *) dp2lut_Xinfo_7 : lut_X_info_7;
  assign _0283_ = _0386_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:15988" *) dp2lut_Xinfo_6 : lut_X_info_6;
  assign _0282_ = _0386_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:15927" *) dp2lut_Xinfo_5 : lut_X_info_5;
  assign _0281_ = _0386_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:15866" *) dp2lut_Xinfo_4 : lut_X_info_4;
  assign _0280_ = load_din ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:15805" *) dp2lut_Xinfo_3 : lut_X_info_3;
  assign _0279_ = load_din ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:15744" *) dp2lut_Xinfo_2 : lut_X_info_2;
  assign _0278_ = load_din ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:15683" *) dp2lut_Xinfo_1 : lut_X_info_1;
  assign _0277_ = load_din ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:15622" *) dp2lut_Xinfo_0 : lut_X_info_0;
  function [15:0] _4524_;
    input [15:0] a;
    input [4095:0] b;
    input [255:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:15605|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *)
    (* parallel_case *)
    casez (s)
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1:
        _4524_ = b[15:0];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?:
        _4524_ = b[31:16];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??:
        _4524_ = b[47:32];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???:
        _4524_ = b[63:48];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????:
        _4524_ = b[79:64];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????:
        _4524_ = b[95:80];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????:
        _4524_ = b[111:96];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????:
        _4524_ = b[127:112];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????:
        _4524_ = b[143:128];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????:
        _4524_ = b[159:144];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????:
        _4524_ = b[175:160];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????:
        _4524_ = b[191:176];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????:
        _4524_ = b[207:192];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????:
        _4524_ = b[223:208];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????:
        _4524_ = b[239:224];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????:
        _4524_ = b[255:240];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????:
        _4524_ = b[271:256];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????:
        _4524_ = b[287:272];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????:
        _4524_ = b[303:288];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????:
        _4524_ = b[319:304];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????:
        _4524_ = b[335:320];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????:
        _4524_ = b[351:336];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????:
        _4524_ = b[367:352];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????:
        _4524_ = b[383:368];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????:
        _4524_ = b[399:384];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????:
        _4524_ = b[415:400];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????:
        _4524_ = b[431:416];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????:
        _4524_ = b[447:432];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????:
        _4524_ = b[463:448];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????:
        _4524_ = b[479:464];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????:
        _4524_ = b[495:480];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????:
        _4524_ = b[511:496];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????:
        _4524_ = b[527:512];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????:
        _4524_ = b[543:528];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????:
        _4524_ = b[559:544];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????:
        _4524_ = b[575:560];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????:
        _4524_ = b[591:576];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????:
        _4524_ = b[607:592];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????:
        _4524_ = b[623:608];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????:
        _4524_ = b[639:624];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????:
        _4524_ = b[655:640];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????:
        _4524_ = b[671:656];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????:
        _4524_ = b[687:672];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????:
        _4524_ = b[703:688];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????:
        _4524_ = b[719:704];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????:
        _4524_ = b[735:720];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????:
        _4524_ = b[751:736];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????:
        _4524_ = b[767:752];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????:
        _4524_ = b[783:768];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????:
        _4524_ = b[799:784];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????:
        _4524_ = b[815:800];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????:
        _4524_ = b[831:816];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????:
        _4524_ = b[847:832];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????:
        _4524_ = b[863:848];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????:
        _4524_ = b[879:864];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????:
        _4524_ = b[895:880];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????:
        _4524_ = b[911:896];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????:
        _4524_ = b[927:912];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????:
        _4524_ = b[943:928];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????:
        _4524_ = b[959:944];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????:
        _4524_ = b[975:960];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????:
        _4524_ = b[991:976];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????:
        _4524_ = b[1007:992];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????:
        _4524_ = b[1023:1008];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????:
        _4524_ = b[1039:1024];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????:
        _4524_ = b[1055:1040];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????:
        _4524_ = b[1071:1056];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????:
        _4524_ = b[1087:1072];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????:
        _4524_ = b[1103:1088];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????:
        _4524_ = b[1119:1104];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????:
        _4524_ = b[1135:1120];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????:
        _4524_ = b[1151:1136];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????:
        _4524_ = b[1167:1152];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????:
        _4524_ = b[1183:1168];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????:
        _4524_ = b[1199:1184];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????:
        _4524_ = b[1215:1200];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????:
        _4524_ = b[1231:1216];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????:
        _4524_ = b[1247:1232];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????:
        _4524_ = b[1263:1248];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????:
        _4524_ = b[1279:1264];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????:
        _4524_ = b[1295:1280];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????:
        _4524_ = b[1311:1296];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????:
        _4524_ = b[1327:1312];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????:
        _4524_ = b[1343:1328];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????:
        _4524_ = b[1359:1344];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????:
        _4524_ = b[1375:1360];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????:
        _4524_ = b[1391:1376];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????:
        _4524_ = b[1407:1392];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????:
        _4524_ = b[1423:1408];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????:
        _4524_ = b[1439:1424];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????:
        _4524_ = b[1455:1440];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????:
        _4524_ = b[1471:1456];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????:
        _4524_ = b[1487:1472];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????:
        _4524_ = b[1503:1488];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????:
        _4524_ = b[1519:1504];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????:
        _4524_ = b[1535:1520];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????:
        _4524_ = b[1551:1536];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????:
        _4524_ = b[1567:1552];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????:
        _4524_ = b[1583:1568];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????:
        _4524_ = b[1599:1584];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4524_ = b[1615:1600];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4524_ = b[1631:1616];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4524_ = b[1647:1632];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4524_ = b[1663:1648];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4524_ = b[1679:1664];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4524_ = b[1695:1680];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4524_ = b[1711:1696];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4524_ = b[1727:1712];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4524_ = b[1743:1728];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4524_ = b[1759:1744];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4524_ = b[1775:1760];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4524_ = b[1791:1776];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4524_ = b[1807:1792];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4524_ = b[1823:1808];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4524_ = b[1839:1824];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4524_ = b[1855:1840];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4524_ = b[1871:1856];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4524_ = b[1887:1872];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4524_ = b[1903:1888];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4524_ = b[1919:1904];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4524_ = b[1935:1920];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4524_ = b[1951:1936];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4524_ = b[1967:1952];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4524_ = b[1983:1968];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4524_ = b[1999:1984];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4524_ = b[2015:2000];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4524_ = b[2031:2016];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4524_ = b[2047:2032];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4524_ = b[2063:2048];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4524_ = b[2079:2064];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4524_ = b[2095:2080];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4524_ = b[2111:2096];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4524_ = b[2127:2112];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4524_ = b[2143:2128];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4524_ = b[2159:2144];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4524_ = b[2175:2160];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4524_ = b[2191:2176];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4524_ = b[2207:2192];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4524_ = b[2223:2208];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4524_ = b[2239:2224];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4524_ = b[2255:2240];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4524_ = b[2271:2256];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4524_ = b[2287:2272];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4524_ = b[2303:2288];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4524_ = b[2319:2304];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4524_ = b[2335:2320];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4524_ = b[2351:2336];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4524_ = b[2367:2352];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4524_ = b[2383:2368];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4524_ = b[2399:2384];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4524_ = b[2415:2400];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4524_ = b[2431:2416];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4524_ = b[2447:2432];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4524_ = b[2463:2448];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4524_ = b[2479:2464];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4524_ = b[2495:2480];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4524_ = b[2511:2496];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4524_ = b[2527:2512];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4524_ = b[2543:2528];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4524_ = b[2559:2544];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4524_ = b[2575:2560];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4524_ = b[2591:2576];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4524_ = b[2607:2592];
      256'b????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4524_ = b[2623:2608];
      256'b???????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4524_ = b[2639:2624];
      256'b??????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4524_ = b[2655:2640];
      256'b?????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4524_ = b[2671:2656];
      256'b????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4524_ = b[2687:2672];
      256'b???????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4524_ = b[2703:2688];
      256'b??????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4524_ = b[2719:2704];
      256'b?????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4524_ = b[2735:2720];
      256'b????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4524_ = b[2751:2736];
      256'b???????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4524_ = b[2767:2752];
      256'b??????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4524_ = b[2783:2768];
      256'b?????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4524_ = b[2799:2784];
      256'b????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4524_ = b[2815:2800];
      256'b???????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4524_ = b[2831:2816];
      256'b??????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4524_ = b[2847:2832];
      256'b?????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4524_ = b[2863:2848];
      256'b????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4524_ = b[2879:2864];
      256'b???????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4524_ = b[2895:2880];
      256'b??????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4524_ = b[2911:2896];
      256'b?????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4524_ = b[2927:2912];
      256'b????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4524_ = b[2943:2928];
      256'b???????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4524_ = b[2959:2944];
      256'b??????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4524_ = b[2975:2960];
      256'b?????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4524_ = b[2991:2976];
      256'b????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4524_ = b[3007:2992];
      256'b???????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4524_ = b[3023:3008];
      256'b??????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4524_ = b[3039:3024];
      256'b?????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4524_ = b[3055:3040];
      256'b????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4524_ = b[3071:3056];
      256'b???????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4524_ = b[3087:3072];
      256'b??????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4524_ = b[3103:3088];
      256'b?????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4524_ = b[3119:3104];
      256'b????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4524_ = b[3135:3120];
      256'b???????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4524_ = b[3151:3136];
      256'b??????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4524_ = b[3167:3152];
      256'b?????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4524_ = b[3183:3168];
      256'b????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4524_ = b[3199:3184];
      256'b???????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4524_ = b[3215:3200];
      256'b??????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4524_ = b[3231:3216];
      256'b?????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4524_ = b[3247:3232];
      256'b????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4524_ = b[3263:3248];
      256'b???????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4524_ = b[3279:3264];
      256'b??????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4524_ = b[3295:3280];
      256'b?????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4524_ = b[3311:3296];
      256'b????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4524_ = b[3327:3312];
      256'b???????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4524_ = b[3343:3328];
      256'b??????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4524_ = b[3359:3344];
      256'b?????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4524_ = b[3375:3360];
      256'b????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4524_ = b[3391:3376];
      256'b???????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4524_ = b[3407:3392];
      256'b??????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4524_ = b[3423:3408];
      256'b?????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4524_ = b[3439:3424];
      256'b????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4524_ = b[3455:3440];
      256'b???????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4524_ = b[3471:3456];
      256'b??????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4524_ = b[3487:3472];
      256'b?????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4524_ = b[3503:3488];
      256'b????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4524_ = b[3519:3504];
      256'b???????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4524_ = b[3535:3520];
      256'b??????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4524_ = b[3551:3536];
      256'b?????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4524_ = b[3567:3552];
      256'b????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4524_ = b[3583:3568];
      256'b???????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4524_ = b[3599:3584];
      256'b??????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4524_ = b[3615:3600];
      256'b?????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4524_ = b[3631:3616];
      256'b????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4524_ = b[3647:3632];
      256'b???????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4524_ = b[3663:3648];
      256'b??????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4524_ = b[3679:3664];
      256'b?????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4524_ = b[3695:3680];
      256'b????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4524_ = b[3711:3696];
      256'b???????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4524_ = b[3727:3712];
      256'b??????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4524_ = b[3743:3728];
      256'b?????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4524_ = b[3759:3744];
      256'b????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4524_ = b[3775:3760];
      256'b???????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4524_ = b[3791:3776];
      256'b??????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4524_ = b[3807:3792];
      256'b?????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4524_ = b[3823:3808];
      256'b????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4524_ = b[3839:3824];
      256'b???????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4524_ = b[3855:3840];
      256'b??????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4524_ = b[3871:3856];
      256'b?????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4524_ = b[3887:3872];
      256'b????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4524_ = b[3903:3888];
      256'b???????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4524_ = b[3919:3904];
      256'b??????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4524_ = b[3935:3920];
      256'b?????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4524_ = b[3951:3936];
      256'b????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4524_ = b[3967:3952];
      256'b???????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4524_ = b[3983:3968];
      256'b??????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4524_ = b[3999:3984];
      256'b?????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4524_ = b[4015:4000];
      256'b????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4524_ = b[4031:4016];
      256'b???1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4524_ = b[4047:4032];
      256'b??1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4524_ = b[4063:4048];
      256'b?1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4524_ = b[4079:4064];
      256'b1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4524_ = b[4095:4080];
      default:
        _4524_ = a;
    endcase
  endfunction
  assign _0681_ = _4524_(density_reg0, { density_reg1, density_reg2, density_reg3, density_reg4, density_reg5, density_reg6, density_reg7, density_reg8, density_reg9, density_reg10, density_reg11, density_reg12, density_reg13, density_reg14, density_reg15, density_reg16, density_reg17, density_reg18, density_reg19, density_reg20, density_reg21, density_reg22, density_reg23, density_reg24, density_reg25, density_reg26, density_reg27, density_reg28, density_reg29, density_reg30, density_reg31, density_reg32, density_reg33, density_reg34, density_reg35, density_reg36, density_reg37, density_reg38, density_reg39, density_reg40, density_reg41, density_reg42, density_reg43, density_reg44, density_reg45, density_reg46, density_reg47, density_reg48, density_reg49, density_reg50, density_reg51, density_reg52, density_reg53, density_reg54, density_reg55, density_reg56, density_reg57, density_reg58, density_reg59, density_reg60, density_reg61, density_reg62, density_reg63, density_reg64, density_reg65, density_reg66, density_reg67, density_reg68, density_reg69, density_reg70, density_reg71, density_reg72, density_reg73, density_reg74, density_reg75, density_reg76, density_reg77, density_reg78, density_reg79, density_reg80, density_reg81, density_reg82, density_reg83, density_reg84, density_reg85, density_reg86, density_reg87, density_reg88, density_reg89, density_reg90, density_reg91, density_reg92, density_reg93, density_reg94, density_reg95, density_reg96, density_reg97, density_reg98, density_reg99, density_reg100, density_reg101, density_reg102, density_reg103, density_reg104, density_reg105, density_reg106, density_reg107, density_reg108, density_reg109, density_reg110, density_reg111, density_reg112, density_reg113, density_reg114, density_reg115, density_reg116, density_reg117, density_reg118, density_reg119, density_reg120, density_reg121, density_reg122, density_reg123, density_reg124, density_reg125, density_reg126, density_reg127, density_reg128, density_reg129, density_reg130, density_reg131, density_reg132, density_reg133, density_reg134, density_reg135, density_reg136, density_reg137, density_reg138, density_reg139, density_reg140, density_reg141, density_reg142, density_reg143, density_reg144, density_reg145, density_reg146, density_reg147, density_reg148, density_reg149, density_reg150, density_reg151, density_reg152, density_reg153, density_reg154, density_reg155, density_reg156, density_reg157, density_reg158, density_reg159, density_reg160, density_reg161, density_reg162, density_reg163, density_reg164, density_reg165, density_reg166, density_reg167, density_reg168, density_reg169, density_reg170, density_reg171, density_reg172, density_reg173, density_reg174, density_reg175, density_reg176, density_reg177, density_reg178, density_reg179, density_reg180, density_reg181, density_reg182, density_reg183, density_reg184, density_reg185, density_reg186, density_reg187, density_reg188, density_reg189, density_reg190, density_reg191, density_reg192, density_reg193, density_reg194, density_reg195, density_reg196, density_reg197, density_reg198, density_reg199, density_reg200, density_reg201, density_reg202, density_reg203, density_reg204, density_reg205, density_reg206, density_reg207, density_reg208, density_reg209, density_reg210, density_reg211, density_reg212, density_reg213, density_reg214, density_reg215, density_reg216, density_reg217, density_reg218, density_reg219, density_reg220, density_reg221, density_reg222, density_reg223, density_reg224, density_reg225, density_reg226, density_reg227, density_reg228, density_reg229, density_reg230, density_reg231, density_reg232, density_reg233, density_reg234, density_reg235, density_reg236, density_reg237, density_reg238, density_reg239, density_reg240, density_reg241, density_reg242, density_reg243, density_reg244, density_reg245, density_reg246, density_reg247, density_reg248, density_reg249, density_reg250, density_reg251, density_reg252, density_reg253, density_reg254, density_reg255, density_reg256 }, { _0938_, _0937_, _0936_, _0935_, _0934_, _0933_, _0932_, _0931_, _0930_, _0929_, _0928_, _0927_, _0926_, _0925_, _0924_, _0923_, _0922_, _0921_, _0920_, _0919_, _0918_, _0917_, _0916_, _0915_, _0914_, _0913_, _0912_, _0911_, _0910_, _0909_, _0908_, _0907_, _0906_, _0905_, _0904_, _0903_, _0902_, _0901_, _0900_, _0899_, _0898_, _0897_, _0896_, _0895_, _0894_, _0893_, _0892_, _0891_, _0890_, _0889_, _0888_, _0887_, _0886_, _0885_, _0884_, _0883_, _0882_, _0881_, _0880_, _0879_, _0878_, _0877_, _0876_, _0875_, _0874_, _0873_, _0872_, _0871_, _0870_, _0869_, _0868_, _0867_, _0866_, _0865_, _0864_, _0863_, _0862_, _0861_, _0860_, _0859_, _0858_, _0857_, _0856_, _0855_, _0854_, _0853_, _0852_, _0851_, _0850_, _0849_, _0848_, _0847_, _0846_, _0845_, _0844_, _0843_, _0842_, _0841_, _0840_, _0839_, _0838_, _0837_, _0836_, _0835_, _0834_, _0833_, _0832_, _0831_, _0830_, _0829_, _0828_, _0827_, _0826_, _0825_, _0824_, _0823_, _0822_, _0821_, _0820_, _0819_, _0818_, _0817_, _0816_, _0815_, _0814_, _0813_, _0812_, _0811_, _0810_, _0809_, _0808_, _0807_, _0806_, _0805_, _0804_, _0803_, _0802_, _0801_, _0800_, _0799_, _0798_, _0797_, _0796_, _0795_, _0794_, _0793_, _0792_, _0791_, _0790_, _0789_, _0788_, _0787_, _0786_, _0785_, _0784_, _0783_, _0782_, _0781_, _0780_, _0779_, _0778_, _0777_, _0776_, _0775_, _0774_, _0773_, _0772_, _0771_, _0770_, _0769_, _0768_, _0767_, _0766_, _0765_, _0764_, _0763_, _0762_, _0761_, _0760_, _0759_, _0758_, _0757_, _0756_, _0755_, _0754_, _0753_, _0752_, _0751_, _0750_, _0749_, _0748_, _0747_, _0746_, _0745_, _0744_, _0743_, _0742_, _0741_, _0740_, _0739_, _0738_, _0737_, _0736_, _0735_, _0734_, _0733_, _0732_, _0731_, _0730_, _0729_, _0728_, _0727_, _0726_, _0725_, _0724_, _0723_, _0722_, _0721_, _0720_, _0719_, _0718_, _0717_, _0716_, _0715_, _0714_, _0713_, _0712_, _0711_, _0710_, _0709_, _0708_, _0707_, _0706_, _0705_, _0704_, _0703_, _0702_, _0701_, _0700_, _0699_, _0698_, _0697_, _0696_, _0695_, _0694_, _0693_, _0692_, _0691_, _0690_, _0689_, _0688_, _0687_, _0686_, _0685_, _0684_, _0412_ });
  assign _0682_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:15605|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 9'b100000000;
  assign _0683_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:15601|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 8'b11111111;
  assign _0684_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:15597|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 8'b11111110;
  assign _0685_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:15593|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 8'b11111101;
  assign _0686_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:15589|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 8'b11111100;
  assign _0687_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:15585|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 8'b11111011;
  assign _0688_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:15581|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 8'b11111010;
  assign _0689_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:15577|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 8'b11111001;
  assign _0690_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:15573|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 8'b11111000;
  assign _0691_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:15569|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 8'b11110111;
  assign _0692_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:15565|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 8'b11110110;
  assign _0693_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:15561|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 8'b11110101;
  assign _0694_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:15557|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 8'b11110100;
  assign _0695_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:15553|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 8'b11110011;
  assign _0696_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:15549|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 8'b11110010;
  assign _0697_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:15545|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 8'b11110001;
  assign _0698_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:15541|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 8'b11110000;
  assign _0699_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:15537|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 8'b11101111;
  assign _0700_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:15533|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 8'b11101110;
  assign _0701_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:15529|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 8'b11101101;
  assign _0702_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:15525|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 8'b11101100;
  assign _0703_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:15521|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 8'b11101011;
  assign _0704_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:15517|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 8'b11101010;
  assign _0705_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:15513|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 8'b11101001;
  assign _0706_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:15509|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 8'b11101000;
  assign _0707_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:15505|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 8'b11100111;
  assign _0708_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:15501|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 8'b11100110;
  assign _0709_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:15497|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 8'b11100101;
  assign _0710_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:15493|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 8'b11100100;
  assign _0711_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:15489|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 8'b11100011;
  assign _0712_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:15485|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 8'b11100010;
  assign _0713_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:15481|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 8'b11100001;
  assign _0714_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:15477|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 8'b11100000;
  assign _0715_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:15473|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 8'b11011111;
  assign _0716_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:15469|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 8'b11011110;
  assign _0717_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:15465|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 8'b11011101;
  assign _0718_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:15461|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 8'b11011100;
  assign _0719_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:15457|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 8'b11011011;
  assign _0720_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:15453|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 8'b11011010;
  assign _0721_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:15449|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 8'b11011001;
  assign _0722_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:15445|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 8'b11011000;
  assign _0723_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:15441|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 8'b11010111;
  assign _0724_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:15437|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 8'b11010110;
  assign _0725_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:15433|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 8'b11010101;
  assign _0726_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:15429|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 8'b11010100;
  assign _0727_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:15425|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 8'b11010011;
  assign _0728_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:15421|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 8'b11010010;
  assign _0729_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:15417|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 8'b11010001;
  assign _0730_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:15413|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 8'b11010000;
  assign _0731_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:15409|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 8'b11001111;
  assign _0732_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:15405|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 8'b11001110;
  assign _0733_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:15401|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 8'b11001101;
  assign _0734_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:15397|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 8'b11001100;
  assign _0735_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:15393|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 8'b11001011;
  assign _0736_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:15389|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 8'b11001010;
  assign _0737_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:15385|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 8'b11001001;
  assign _0738_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:15381|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 8'b11001000;
  assign _0739_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:15377|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 8'b11000111;
  assign _0740_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:15373|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 8'b11000110;
  assign _0741_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:15369|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 8'b11000101;
  assign _0742_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:15365|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 8'b11000100;
  assign _0743_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:15361|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 8'b11000011;
  assign _0744_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:15357|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 8'b11000010;
  assign _0745_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:15353|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 8'b11000001;
  assign _0746_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:15349|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 8'b11000000;
  assign _0747_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:15345|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 8'b10111111;
  assign _0748_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:15341|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 8'b10111110;
  assign _0749_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:15337|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 8'b10111101;
  assign _0750_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:15333|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 8'b10111100;
  assign _0751_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:15329|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 8'b10111011;
  assign _0752_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:15325|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 8'b10111010;
  assign _0753_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:15321|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 8'b10111001;
  assign _0754_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:15317|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 8'b10111000;
  assign _0755_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:15313|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 8'b10110111;
  assign _0756_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:15309|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 8'b10110110;
  assign _0757_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:15305|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 8'b10110101;
  assign _0758_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:15301|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 8'b10110100;
  assign _0759_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:15297|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 8'b10110011;
  assign _0760_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:15293|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 8'b10110010;
  assign _0761_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:15289|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 8'b10110001;
  assign _0762_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:15285|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 8'b10110000;
  assign _0763_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:15281|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 8'b10101111;
  assign _0764_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:15277|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 8'b10101110;
  assign _0765_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:15273|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 8'b10101101;
  assign _0766_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:15269|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 8'b10101100;
  assign _0767_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:15265|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 8'b10101011;
  assign _0768_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:15261|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 8'b10101010;
  assign _0769_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:15257|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 8'b10101001;
  assign _0770_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:15253|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 8'b10101000;
  assign _0771_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:15249|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 8'b10100111;
  assign _0772_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:15245|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 8'b10100110;
  assign _0773_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:15241|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 8'b10100101;
  assign _0774_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:15237|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 8'b10100100;
  assign _0775_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:15233|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 8'b10100011;
  assign _0776_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:15229|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 8'b10100010;
  assign _0777_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:15225|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 8'b10100001;
  assign _0778_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:15221|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 8'b10100000;
  assign _0779_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:15217|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 8'b10011111;
  assign _0780_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:15213|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 8'b10011110;
  assign _0781_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:15209|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 8'b10011101;
  assign _0782_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:15205|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 8'b10011100;
  assign _0783_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:15201|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 8'b10011011;
  assign _0784_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:15197|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 8'b10011010;
  assign _0785_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:15193|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 8'b10011001;
  assign _0786_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:15189|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 8'b10011000;
  assign _0787_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:15185|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 8'b10010111;
  assign _0788_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:15181|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 8'b10010110;
  assign _0789_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:15177|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 8'b10010101;
  assign _0790_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:15173|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 8'b10010100;
  assign _0791_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:15169|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 8'b10010011;
  assign _0792_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:15165|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 8'b10010010;
  assign _0793_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:15161|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 8'b10010001;
  assign _0794_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:15157|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 8'b10010000;
  assign _0795_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:15153|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 8'b10001111;
  assign _0796_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:15149|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 8'b10001110;
  assign _0797_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:15145|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 8'b10001101;
  assign _0798_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:15141|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 8'b10001100;
  assign _0799_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:15137|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 8'b10001011;
  assign _0800_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:15133|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 8'b10001010;
  assign _0801_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:15129|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 8'b10001001;
  assign _0802_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:15125|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 8'b10001000;
  assign _0803_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:15121|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 8'b10000111;
  assign _0804_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:15117|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 8'b10000110;
  assign _0805_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:15113|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 8'b10000101;
  assign _0806_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:15109|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 8'b10000100;
  assign _0807_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:15105|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 8'b10000011;
  assign _0808_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:15101|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 8'b10000010;
  assign _0809_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:15097|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 8'b10000001;
  assign _0810_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:15093|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 8'b10000000;
  assign _0811_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:15089|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 7'b1111111;
  assign _0812_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:15085|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 7'b1111110;
  assign _0813_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:15081|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 7'b1111101;
  assign _0814_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:15077|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 7'b1111100;
  assign _0815_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:15073|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 7'b1111011;
  assign _0816_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:15069|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 7'b1111010;
  assign _0817_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:15065|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 7'b1111001;
  assign _0818_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:15061|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 7'b1111000;
  assign _0819_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:15057|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 7'b1110111;
  assign _0820_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:15053|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 7'b1110110;
  assign _0821_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:15049|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 7'b1110101;
  assign _0822_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:15045|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 7'b1110100;
  assign _0823_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:15041|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 7'b1110011;
  assign _0824_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:15037|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 7'b1110010;
  assign _0825_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:15033|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 7'b1110001;
  assign _0826_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:15029|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 7'b1110000;
  assign _0827_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:15025|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 7'b1101111;
  assign _0828_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:15021|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 7'b1101110;
  assign _0829_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:15017|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 7'b1101101;
  assign _0830_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:15013|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 7'b1101100;
  assign _0831_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:15009|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 7'b1101011;
  assign _0832_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:15005|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 7'b1101010;
  assign _0833_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:15001|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 7'b1101001;
  assign _0834_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14997|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 7'b1101000;
  assign _0835_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14993|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 7'b1100111;
  assign _0836_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14989|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 7'b1100110;
  assign _0837_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14985|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 7'b1100101;
  assign _0838_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14981|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 7'b1100100;
  assign _0839_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14977|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 7'b1100011;
  assign _0840_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14973|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 7'b1100010;
  assign _0841_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14969|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 7'b1100001;
  assign _0842_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14965|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 7'b1100000;
  assign _0843_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14961|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 7'b1011111;
  assign _0844_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14957|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 7'b1011110;
  assign _0845_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14953|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 7'b1011101;
  assign _0846_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14949|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 7'b1011100;
  assign _0847_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14945|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 7'b1011011;
  assign _0848_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14941|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 7'b1011010;
  assign _0849_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14937|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 7'b1011001;
  assign _0850_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14933|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 7'b1011000;
  assign _0851_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14929|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 7'b1010111;
  assign _0852_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14925|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 7'b1010110;
  assign _0853_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14921|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 7'b1010101;
  assign _0854_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14917|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 7'b1010100;
  assign _0855_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14913|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 7'b1010011;
  assign _0856_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14909|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 7'b1010010;
  assign _0857_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14905|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 7'b1010001;
  assign _0858_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14901|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 7'b1010000;
  assign _0859_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14897|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 7'b1001111;
  assign _0860_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14893|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 7'b1001110;
  assign _0861_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14889|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 7'b1001101;
  assign _0862_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14885|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 7'b1001100;
  assign _0863_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14881|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 7'b1001011;
  assign _0864_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14877|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 7'b1001010;
  assign _0865_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14873|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 7'b1001001;
  assign _0866_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14869|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 7'b1001000;
  assign _0867_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14865|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 7'b1000111;
  assign _0868_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14861|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 7'b1000110;
  assign _0869_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14857|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 7'b1000101;
  assign _0870_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14853|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 7'b1000100;
  assign _0871_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14849|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 7'b1000011;
  assign _0872_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14845|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 7'b1000010;
  assign _0873_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14841|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 7'b1000001;
  assign _0874_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14837|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 7'b1000000;
  assign _0875_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14833|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 6'b111111;
  assign _0876_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14829|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 6'b111110;
  assign _0877_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14825|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 6'b111101;
  assign _0878_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14821|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 6'b111100;
  assign _0879_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14817|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 6'b111011;
  assign _0880_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14813|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 6'b111010;
  assign _0881_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14809|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 6'b111001;
  assign _0882_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14805|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 6'b111000;
  assign _0883_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14801|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 6'b110111;
  assign _0884_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14797|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 6'b110110;
  assign _0885_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14793|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 6'b110101;
  assign _0886_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14789|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 6'b110100;
  assign _0887_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14785|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 6'b110011;
  assign _0888_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14781|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 6'b110010;
  assign _0889_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14777|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 6'b110001;
  assign _0890_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14773|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 6'b110000;
  assign _0891_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14769|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 6'b101111;
  assign _0892_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14765|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 6'b101110;
  assign _0893_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14761|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 6'b101101;
  assign _0894_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14757|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 6'b101100;
  assign _0895_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14753|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 6'b101011;
  assign _0896_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14749|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 6'b101010;
  assign _0897_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14745|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 6'b101001;
  assign _0898_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14741|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 6'b101000;
  assign _0899_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14737|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 6'b100111;
  assign _0900_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14733|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 6'b100110;
  assign _0901_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14729|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 6'b100101;
  assign _0902_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14725|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 6'b100100;
  assign _0903_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14721|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 6'b100011;
  assign _0904_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14717|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 6'b100010;
  assign _0905_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14713|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 6'b100001;
  assign _0906_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14709|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 6'b100000;
  assign _0907_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14705|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 5'b11111;
  assign _0908_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14701|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 5'b11110;
  assign _0909_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14697|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 5'b11101;
  assign _0910_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14693|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 5'b11100;
  assign _0911_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14689|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 5'b11011;
  assign _0912_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14685|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 5'b11010;
  assign _0913_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14681|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 5'b11001;
  assign _0914_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14677|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 5'b11000;
  assign _0915_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14673|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 5'b10111;
  assign _0916_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14669|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 5'b10110;
  assign _0917_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14665|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 5'b10101;
  assign _0918_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14661|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 5'b10100;
  assign _0919_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14657|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 5'b10011;
  assign _0920_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14653|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 5'b10010;
  assign _0921_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14649|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 5'b10001;
  assign _0922_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14645|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 5'b10000;
  assign _0923_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14641|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 4'b1111;
  assign _0924_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14637|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 4'b1110;
  assign _0925_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14633|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 4'b1101;
  assign _0926_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14629|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 4'b1100;
  assign _0927_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14625|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 4'b1011;
  assign _0928_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14621|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 4'b1010;
  assign _0929_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14617|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 4'b1001;
  assign _0930_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14613|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 4'b1000;
  assign _0931_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14609|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 3'b111;
  assign _0932_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14605|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 3'b110;
  assign _0933_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14601|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 3'b101;
  assign _0934_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14597|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 3'b100;
  assign _0935_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14593|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 2'b11;
  assign _0936_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14589|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 2'b10;
  assign _0937_ = dp2lut_Y_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14585|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) 1'b1;
  assign _0938_ = ! (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14581|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *) dp2lut_Y_entry_7;
  assign _0939_ = dp2lut_Yinfo_7[17] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14576" *) density_reg256 : _0681_;
  assign _0940_ = dp2lut_Yinfo_7[16] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14573" *) density_reg0 : _0939_;
  assign _0300_ = _0391_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14572" *) _0940_ : lut_Y_data_71;
  function [15:0] _4785_;
    input [15:0] a;
    input [4095:0] b;
    input [255:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:15605|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14580" *)
    (* parallel_case *)
    casez (s)
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1:
        _4785_ = b[15:0];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?:
        _4785_ = b[31:16];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??:
        _4785_ = b[47:32];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???:
        _4785_ = b[63:48];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????:
        _4785_ = b[79:64];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????:
        _4785_ = b[95:80];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????:
        _4785_ = b[111:96];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????:
        _4785_ = b[127:112];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????:
        _4785_ = b[143:128];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????:
        _4785_ = b[159:144];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????:
        _4785_ = b[175:160];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????:
        _4785_ = b[191:176];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????:
        _4785_ = b[207:192];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????:
        _4785_ = b[223:208];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????:
        _4785_ = b[239:224];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????:
        _4785_ = b[255:240];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????:
        _4785_ = b[271:256];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????:
        _4785_ = b[287:272];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????:
        _4785_ = b[303:288];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????:
        _4785_ = b[319:304];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????:
        _4785_ = b[335:320];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????:
        _4785_ = b[351:336];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????:
        _4785_ = b[367:352];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????:
        _4785_ = b[383:368];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????:
        _4785_ = b[399:384];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????:
        _4785_ = b[415:400];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????:
        _4785_ = b[431:416];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????:
        _4785_ = b[447:432];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????:
        _4785_ = b[463:448];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????:
        _4785_ = b[479:464];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????:
        _4785_ = b[495:480];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????:
        _4785_ = b[511:496];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????:
        _4785_ = b[527:512];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????:
        _4785_ = b[543:528];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????:
        _4785_ = b[559:544];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????:
        _4785_ = b[575:560];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????:
        _4785_ = b[591:576];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????:
        _4785_ = b[607:592];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????:
        _4785_ = b[623:608];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????:
        _4785_ = b[639:624];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????:
        _4785_ = b[655:640];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????:
        _4785_ = b[671:656];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????:
        _4785_ = b[687:672];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????:
        _4785_ = b[703:688];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????:
        _4785_ = b[719:704];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????:
        _4785_ = b[735:720];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????:
        _4785_ = b[751:736];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????:
        _4785_ = b[767:752];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????:
        _4785_ = b[783:768];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????:
        _4785_ = b[799:784];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????:
        _4785_ = b[815:800];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????:
        _4785_ = b[831:816];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????:
        _4785_ = b[847:832];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????:
        _4785_ = b[863:848];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????:
        _4785_ = b[879:864];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????:
        _4785_ = b[895:880];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????:
        _4785_ = b[911:896];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????:
        _4785_ = b[927:912];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????:
        _4785_ = b[943:928];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????:
        _4785_ = b[959:944];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????:
        _4785_ = b[975:960];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????:
        _4785_ = b[991:976];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????:
        _4785_ = b[1007:992];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????:
        _4785_ = b[1023:1008];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????:
        _4785_ = b[1039:1024];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????:
        _4785_ = b[1055:1040];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????:
        _4785_ = b[1071:1056];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????:
        _4785_ = b[1087:1072];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????:
        _4785_ = b[1103:1088];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????:
        _4785_ = b[1119:1104];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????:
        _4785_ = b[1135:1120];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????:
        _4785_ = b[1151:1136];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????:
        _4785_ = b[1167:1152];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????:
        _4785_ = b[1183:1168];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????:
        _4785_ = b[1199:1184];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????:
        _4785_ = b[1215:1200];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????:
        _4785_ = b[1231:1216];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????:
        _4785_ = b[1247:1232];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????:
        _4785_ = b[1263:1248];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????:
        _4785_ = b[1279:1264];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????:
        _4785_ = b[1295:1280];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????:
        _4785_ = b[1311:1296];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????:
        _4785_ = b[1327:1312];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????:
        _4785_ = b[1343:1328];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????:
        _4785_ = b[1359:1344];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????:
        _4785_ = b[1375:1360];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????:
        _4785_ = b[1391:1376];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????:
        _4785_ = b[1407:1392];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????:
        _4785_ = b[1423:1408];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????:
        _4785_ = b[1439:1424];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????:
        _4785_ = b[1455:1440];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????:
        _4785_ = b[1471:1456];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????:
        _4785_ = b[1487:1472];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????:
        _4785_ = b[1503:1488];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????:
        _4785_ = b[1519:1504];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????:
        _4785_ = b[1535:1520];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????:
        _4785_ = b[1551:1536];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????:
        _4785_ = b[1567:1552];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????:
        _4785_ = b[1583:1568];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????:
        _4785_ = b[1599:1584];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4785_ = b[1615:1600];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4785_ = b[1631:1616];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4785_ = b[1647:1632];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4785_ = b[1663:1648];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4785_ = b[1679:1664];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4785_ = b[1695:1680];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4785_ = b[1711:1696];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4785_ = b[1727:1712];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4785_ = b[1743:1728];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4785_ = b[1759:1744];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4785_ = b[1775:1760];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4785_ = b[1791:1776];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4785_ = b[1807:1792];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4785_ = b[1823:1808];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4785_ = b[1839:1824];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4785_ = b[1855:1840];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4785_ = b[1871:1856];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4785_ = b[1887:1872];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4785_ = b[1903:1888];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4785_ = b[1919:1904];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4785_ = b[1935:1920];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4785_ = b[1951:1936];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4785_ = b[1967:1952];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4785_ = b[1983:1968];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4785_ = b[1999:1984];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4785_ = b[2015:2000];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4785_ = b[2031:2016];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4785_ = b[2047:2032];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4785_ = b[2063:2048];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4785_ = b[2079:2064];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4785_ = b[2095:2080];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4785_ = b[2111:2096];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4785_ = b[2127:2112];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4785_ = b[2143:2128];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4785_ = b[2159:2144];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4785_ = b[2175:2160];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4785_ = b[2191:2176];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4785_ = b[2207:2192];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4785_ = b[2223:2208];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4785_ = b[2239:2224];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4785_ = b[2255:2240];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4785_ = b[2271:2256];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4785_ = b[2287:2272];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4785_ = b[2303:2288];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4785_ = b[2319:2304];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4785_ = b[2335:2320];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4785_ = b[2351:2336];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4785_ = b[2367:2352];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4785_ = b[2383:2368];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4785_ = b[2399:2384];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4785_ = b[2415:2400];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4785_ = b[2431:2416];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4785_ = b[2447:2432];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4785_ = b[2463:2448];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4785_ = b[2479:2464];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4785_ = b[2495:2480];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4785_ = b[2511:2496];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4785_ = b[2527:2512];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4785_ = b[2543:2528];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4785_ = b[2559:2544];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4785_ = b[2575:2560];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4785_ = b[2591:2576];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4785_ = b[2607:2592];
      256'b????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4785_ = b[2623:2608];
      256'b???????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4785_ = b[2639:2624];
      256'b??????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4785_ = b[2655:2640];
      256'b?????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4785_ = b[2671:2656];
      256'b????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4785_ = b[2687:2672];
      256'b???????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4785_ = b[2703:2688];
      256'b??????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4785_ = b[2719:2704];
      256'b?????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4785_ = b[2735:2720];
      256'b????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4785_ = b[2751:2736];
      256'b???????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4785_ = b[2767:2752];
      256'b??????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4785_ = b[2783:2768];
      256'b?????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4785_ = b[2799:2784];
      256'b????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4785_ = b[2815:2800];
      256'b???????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4785_ = b[2831:2816];
      256'b??????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4785_ = b[2847:2832];
      256'b?????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4785_ = b[2863:2848];
      256'b????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4785_ = b[2879:2864];
      256'b???????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4785_ = b[2895:2880];
      256'b??????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4785_ = b[2911:2896];
      256'b?????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4785_ = b[2927:2912];
      256'b????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4785_ = b[2943:2928];
      256'b???????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4785_ = b[2959:2944];
      256'b??????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4785_ = b[2975:2960];
      256'b?????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4785_ = b[2991:2976];
      256'b????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4785_ = b[3007:2992];
      256'b???????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4785_ = b[3023:3008];
      256'b??????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4785_ = b[3039:3024];
      256'b?????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4785_ = b[3055:3040];
      256'b????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4785_ = b[3071:3056];
      256'b???????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4785_ = b[3087:3072];
      256'b??????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4785_ = b[3103:3088];
      256'b?????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4785_ = b[3119:3104];
      256'b????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4785_ = b[3135:3120];
      256'b???????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4785_ = b[3151:3136];
      256'b??????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4785_ = b[3167:3152];
      256'b?????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4785_ = b[3183:3168];
      256'b????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4785_ = b[3199:3184];
      256'b???????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4785_ = b[3215:3200];
      256'b??????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4785_ = b[3231:3216];
      256'b?????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4785_ = b[3247:3232];
      256'b????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4785_ = b[3263:3248];
      256'b???????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4785_ = b[3279:3264];
      256'b??????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4785_ = b[3295:3280];
      256'b?????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4785_ = b[3311:3296];
      256'b????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4785_ = b[3327:3312];
      256'b???????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4785_ = b[3343:3328];
      256'b??????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4785_ = b[3359:3344];
      256'b?????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4785_ = b[3375:3360];
      256'b????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4785_ = b[3391:3376];
      256'b???????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4785_ = b[3407:3392];
      256'b??????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4785_ = b[3423:3408];
      256'b?????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4785_ = b[3439:3424];
      256'b????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4785_ = b[3455:3440];
      256'b???????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4785_ = b[3471:3456];
      256'b??????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4785_ = b[3487:3472];
      256'b?????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4785_ = b[3503:3488];
      256'b????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4785_ = b[3519:3504];
      256'b???????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4785_ = b[3535:3520];
      256'b??????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4785_ = b[3551:3536];
      256'b?????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4785_ = b[3567:3552];
      256'b????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4785_ = b[3583:3568];
      256'b???????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4785_ = b[3599:3584];
      256'b??????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4785_ = b[3615:3600];
      256'b?????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4785_ = b[3631:3616];
      256'b????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4785_ = b[3647:3632];
      256'b???????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4785_ = b[3663:3648];
      256'b??????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4785_ = b[3679:3664];
      256'b?????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4785_ = b[3695:3680];
      256'b????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4785_ = b[3711:3696];
      256'b???????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4785_ = b[3727:3712];
      256'b??????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4785_ = b[3743:3728];
      256'b?????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4785_ = b[3759:3744];
      256'b????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4785_ = b[3775:3760];
      256'b???????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4785_ = b[3791:3776];
      256'b??????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4785_ = b[3807:3792];
      256'b?????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4785_ = b[3823:3808];
      256'b????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4785_ = b[3839:3824];
      256'b???????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4785_ = b[3855:3840];
      256'b??????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4785_ = b[3871:3856];
      256'b?????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4785_ = b[3887:3872];
      256'b????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4785_ = b[3903:3888];
      256'b???????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4785_ = b[3919:3904];
      256'b??????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4785_ = b[3935:3920];
      256'b?????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4785_ = b[3951:3936];
      256'b????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4785_ = b[3967:3952];
      256'b???????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4785_ = b[3983:3968];
      256'b??????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4785_ = b[3999:3984];
      256'b?????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4785_ = b[4015:4000];
      256'b????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4785_ = b[4031:4016];
      256'b???1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4785_ = b[4047:4032];
      256'b??1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4785_ = b[4063:4048];
      256'b?1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4785_ = b[4079:4064];
      256'b1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4785_ = b[4095:4080];
      default:
        _4785_ = a;
    endcase
  endfunction
  assign _0941_ = _4785_(density_reg0, { density_reg1, density_reg2, density_reg3, density_reg4, density_reg5, density_reg6, density_reg7, density_reg8, density_reg9, density_reg10, density_reg11, density_reg12, density_reg13, density_reg14, density_reg15, density_reg16, density_reg17, density_reg18, density_reg19, density_reg20, density_reg21, density_reg22, density_reg23, density_reg24, density_reg25, density_reg26, density_reg27, density_reg28, density_reg29, density_reg30, density_reg31, density_reg32, density_reg33, density_reg34, density_reg35, density_reg36, density_reg37, density_reg38, density_reg39, density_reg40, density_reg41, density_reg42, density_reg43, density_reg44, density_reg45, density_reg46, density_reg47, density_reg48, density_reg49, density_reg50, density_reg51, density_reg52, density_reg53, density_reg54, density_reg55, density_reg56, density_reg57, density_reg58, density_reg59, density_reg60, density_reg61, density_reg62, density_reg63, density_reg64, density_reg65, density_reg66, density_reg67, density_reg68, density_reg69, density_reg70, density_reg71, density_reg72, density_reg73, density_reg74, density_reg75, density_reg76, density_reg77, density_reg78, density_reg79, density_reg80, density_reg81, density_reg82, density_reg83, density_reg84, density_reg85, density_reg86, density_reg87, density_reg88, density_reg89, density_reg90, density_reg91, density_reg92, density_reg93, density_reg94, density_reg95, density_reg96, density_reg97, density_reg98, density_reg99, density_reg100, density_reg101, density_reg102, density_reg103, density_reg104, density_reg105, density_reg106, density_reg107, density_reg108, density_reg109, density_reg110, density_reg111, density_reg112, density_reg113, density_reg114, density_reg115, density_reg116, density_reg117, density_reg118, density_reg119, density_reg120, density_reg121, density_reg122, density_reg123, density_reg124, density_reg125, density_reg126, density_reg127, density_reg128, density_reg129, density_reg130, density_reg131, density_reg132, density_reg133, density_reg134, density_reg135, density_reg136, density_reg137, density_reg138, density_reg139, density_reg140, density_reg141, density_reg142, density_reg143, density_reg144, density_reg145, density_reg146, density_reg147, density_reg148, density_reg149, density_reg150, density_reg151, density_reg152, density_reg153, density_reg154, density_reg155, density_reg156, density_reg157, density_reg158, density_reg159, density_reg160, density_reg161, density_reg162, density_reg163, density_reg164, density_reg165, density_reg166, density_reg167, density_reg168, density_reg169, density_reg170, density_reg171, density_reg172, density_reg173, density_reg174, density_reg175, density_reg176, density_reg177, density_reg178, density_reg179, density_reg180, density_reg181, density_reg182, density_reg183, density_reg184, density_reg185, density_reg186, density_reg187, density_reg188, density_reg189, density_reg190, density_reg191, density_reg192, density_reg193, density_reg194, density_reg195, density_reg196, density_reg197, density_reg198, density_reg199, density_reg200, density_reg201, density_reg202, density_reg203, density_reg204, density_reg205, density_reg206, density_reg207, density_reg208, density_reg209, density_reg210, density_reg211, density_reg212, density_reg213, density_reg214, density_reg215, density_reg216, density_reg217, density_reg218, density_reg219, density_reg220, density_reg221, density_reg222, density_reg223, density_reg224, density_reg225, density_reg226, density_reg227, density_reg228, density_reg229, density_reg230, density_reg231, density_reg232, density_reg233, density_reg234, density_reg235, density_reg236, density_reg237, density_reg238, density_reg239, density_reg240, density_reg241, density_reg242, density_reg243, density_reg244, density_reg245, density_reg246, density_reg247, density_reg248, density_reg249, density_reg250, density_reg251, density_reg252, density_reg253, density_reg254, density_reg255, density_reg256 }, { _0937_, _0936_, _0935_, _0934_, _0933_, _0932_, _0931_, _0930_, _0929_, _0928_, _0927_, _0926_, _0925_, _0924_, _0923_, _0922_, _0921_, _0920_, _0919_, _0918_, _0917_, _0916_, _0915_, _0914_, _0913_, _0912_, _0911_, _0910_, _0909_, _0908_, _0907_, _0906_, _0905_, _0904_, _0903_, _0902_, _0901_, _0900_, _0899_, _0898_, _0897_, _0896_, _0895_, _0894_, _0893_, _0892_, _0891_, _0890_, _0889_, _0888_, _0887_, _0886_, _0885_, _0884_, _0883_, _0882_, _0881_, _0880_, _0879_, _0878_, _0877_, _0876_, _0875_, _0874_, _0873_, _0872_, _0871_, _0870_, _0869_, _0868_, _0867_, _0866_, _0865_, _0864_, _0863_, _0862_, _0861_, _0860_, _0859_, _0858_, _0857_, _0856_, _0855_, _0854_, _0853_, _0852_, _0851_, _0850_, _0849_, _0848_, _0847_, _0846_, _0845_, _0844_, _0843_, _0842_, _0841_, _0840_, _0839_, _0838_, _0837_, _0836_, _0835_, _0834_, _0833_, _0832_, _0831_, _0830_, _0829_, _0828_, _0827_, _0826_, _0825_, _0824_, _0823_, _0822_, _0821_, _0820_, _0819_, _0818_, _0817_, _0816_, _0815_, _0814_, _0813_, _0812_, _0811_, _0810_, _0809_, _0808_, _0807_, _0806_, _0805_, _0804_, _0803_, _0802_, _0801_, _0800_, _0799_, _0798_, _0797_, _0796_, _0795_, _0794_, _0793_, _0792_, _0791_, _0790_, _0789_, _0788_, _0787_, _0786_, _0785_, _0784_, _0783_, _0782_, _0781_, _0780_, _0779_, _0778_, _0777_, _0776_, _0775_, _0774_, _0773_, _0772_, _0771_, _0770_, _0769_, _0768_, _0767_, _0766_, _0765_, _0764_, _0763_, _0762_, _0761_, _0760_, _0759_, _0758_, _0757_, _0756_, _0755_, _0754_, _0753_, _0752_, _0751_, _0750_, _0749_, _0748_, _0747_, _0746_, _0745_, _0744_, _0743_, _0742_, _0741_, _0740_, _0739_, _0738_, _0737_, _0736_, _0735_, _0734_, _0733_, _0732_, _0731_, _0730_, _0729_, _0728_, _0727_, _0726_, _0725_, _0724_, _0723_, _0722_, _0721_, _0720_, _0719_, _0718_, _0717_, _0716_, _0715_, _0714_, _0713_, _0712_, _0711_, _0710_, _0709_, _0708_, _0707_, _0706_, _0705_, _0704_, _0703_, _0702_, _0701_, _0700_, _0699_, _0698_, _0697_, _0696_, _0695_, _0694_, _0693_, _0692_, _0691_, _0690_, _0689_, _0688_, _0687_, _0686_, _0685_, _0684_, _0683_, _0682_ });
  assign _0942_ = dp2lut_Yinfo_7[17] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14576" *) density_reg256 : _0941_;
  assign _0943_ = dp2lut_Yinfo_7[16] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14573" *) density_reg0 : _0942_;
  assign _0299_ = _0391_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14572" *) _0943_ : lut_Y_data_70;
  function [15:0] _4789_;
    input [15:0] a;
    input [4095:0] b;
    input [255:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14554|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *)
    (* parallel_case *)
    casez (s)
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1:
        _4789_ = b[15:0];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?:
        _4789_ = b[31:16];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??:
        _4789_ = b[47:32];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???:
        _4789_ = b[63:48];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????:
        _4789_ = b[79:64];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????:
        _4789_ = b[95:80];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????:
        _4789_ = b[111:96];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????:
        _4789_ = b[127:112];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????:
        _4789_ = b[143:128];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????:
        _4789_ = b[159:144];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????:
        _4789_ = b[175:160];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????:
        _4789_ = b[191:176];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????:
        _4789_ = b[207:192];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????:
        _4789_ = b[223:208];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????:
        _4789_ = b[239:224];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????:
        _4789_ = b[255:240];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????:
        _4789_ = b[271:256];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????:
        _4789_ = b[287:272];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????:
        _4789_ = b[303:288];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????:
        _4789_ = b[319:304];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????:
        _4789_ = b[335:320];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????:
        _4789_ = b[351:336];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????:
        _4789_ = b[367:352];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????:
        _4789_ = b[383:368];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????:
        _4789_ = b[399:384];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????:
        _4789_ = b[415:400];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????:
        _4789_ = b[431:416];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????:
        _4789_ = b[447:432];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????:
        _4789_ = b[463:448];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????:
        _4789_ = b[479:464];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????:
        _4789_ = b[495:480];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????:
        _4789_ = b[511:496];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????:
        _4789_ = b[527:512];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????:
        _4789_ = b[543:528];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????:
        _4789_ = b[559:544];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????:
        _4789_ = b[575:560];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????:
        _4789_ = b[591:576];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????:
        _4789_ = b[607:592];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????:
        _4789_ = b[623:608];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????:
        _4789_ = b[639:624];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????:
        _4789_ = b[655:640];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????:
        _4789_ = b[671:656];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????:
        _4789_ = b[687:672];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????:
        _4789_ = b[703:688];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????:
        _4789_ = b[719:704];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????:
        _4789_ = b[735:720];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????:
        _4789_ = b[751:736];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????:
        _4789_ = b[767:752];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????:
        _4789_ = b[783:768];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????:
        _4789_ = b[799:784];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????:
        _4789_ = b[815:800];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????:
        _4789_ = b[831:816];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????:
        _4789_ = b[847:832];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????:
        _4789_ = b[863:848];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????:
        _4789_ = b[879:864];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????:
        _4789_ = b[895:880];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????:
        _4789_ = b[911:896];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????:
        _4789_ = b[927:912];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????:
        _4789_ = b[943:928];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????:
        _4789_ = b[959:944];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????:
        _4789_ = b[975:960];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????:
        _4789_ = b[991:976];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????:
        _4789_ = b[1007:992];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????:
        _4789_ = b[1023:1008];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????:
        _4789_ = b[1039:1024];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????:
        _4789_ = b[1055:1040];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????:
        _4789_ = b[1071:1056];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????:
        _4789_ = b[1087:1072];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????:
        _4789_ = b[1103:1088];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????:
        _4789_ = b[1119:1104];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????:
        _4789_ = b[1135:1120];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????:
        _4789_ = b[1151:1136];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????:
        _4789_ = b[1167:1152];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????:
        _4789_ = b[1183:1168];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????:
        _4789_ = b[1199:1184];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????:
        _4789_ = b[1215:1200];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????:
        _4789_ = b[1231:1216];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????:
        _4789_ = b[1247:1232];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????:
        _4789_ = b[1263:1248];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????:
        _4789_ = b[1279:1264];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????:
        _4789_ = b[1295:1280];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????:
        _4789_ = b[1311:1296];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????:
        _4789_ = b[1327:1312];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????:
        _4789_ = b[1343:1328];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????:
        _4789_ = b[1359:1344];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????:
        _4789_ = b[1375:1360];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????:
        _4789_ = b[1391:1376];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????:
        _4789_ = b[1407:1392];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????:
        _4789_ = b[1423:1408];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????:
        _4789_ = b[1439:1424];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????:
        _4789_ = b[1455:1440];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????:
        _4789_ = b[1471:1456];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????:
        _4789_ = b[1487:1472];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????:
        _4789_ = b[1503:1488];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????:
        _4789_ = b[1519:1504];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????:
        _4789_ = b[1535:1520];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????:
        _4789_ = b[1551:1536];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????:
        _4789_ = b[1567:1552];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????:
        _4789_ = b[1583:1568];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????:
        _4789_ = b[1599:1584];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4789_ = b[1615:1600];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4789_ = b[1631:1616];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4789_ = b[1647:1632];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4789_ = b[1663:1648];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4789_ = b[1679:1664];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4789_ = b[1695:1680];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4789_ = b[1711:1696];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4789_ = b[1727:1712];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4789_ = b[1743:1728];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4789_ = b[1759:1744];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4789_ = b[1775:1760];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4789_ = b[1791:1776];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4789_ = b[1807:1792];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4789_ = b[1823:1808];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4789_ = b[1839:1824];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4789_ = b[1855:1840];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4789_ = b[1871:1856];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4789_ = b[1887:1872];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4789_ = b[1903:1888];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4789_ = b[1919:1904];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4789_ = b[1935:1920];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4789_ = b[1951:1936];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4789_ = b[1967:1952];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4789_ = b[1983:1968];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4789_ = b[1999:1984];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4789_ = b[2015:2000];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4789_ = b[2031:2016];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4789_ = b[2047:2032];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4789_ = b[2063:2048];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4789_ = b[2079:2064];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4789_ = b[2095:2080];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4789_ = b[2111:2096];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4789_ = b[2127:2112];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4789_ = b[2143:2128];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4789_ = b[2159:2144];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4789_ = b[2175:2160];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4789_ = b[2191:2176];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4789_ = b[2207:2192];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4789_ = b[2223:2208];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4789_ = b[2239:2224];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4789_ = b[2255:2240];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4789_ = b[2271:2256];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4789_ = b[2287:2272];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4789_ = b[2303:2288];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4789_ = b[2319:2304];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4789_ = b[2335:2320];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4789_ = b[2351:2336];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4789_ = b[2367:2352];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4789_ = b[2383:2368];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4789_ = b[2399:2384];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4789_ = b[2415:2400];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4789_ = b[2431:2416];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4789_ = b[2447:2432];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4789_ = b[2463:2448];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4789_ = b[2479:2464];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4789_ = b[2495:2480];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4789_ = b[2511:2496];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4789_ = b[2527:2512];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4789_ = b[2543:2528];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4789_ = b[2559:2544];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4789_ = b[2575:2560];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4789_ = b[2591:2576];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4789_ = b[2607:2592];
      256'b????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4789_ = b[2623:2608];
      256'b???????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4789_ = b[2639:2624];
      256'b??????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4789_ = b[2655:2640];
      256'b?????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4789_ = b[2671:2656];
      256'b????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4789_ = b[2687:2672];
      256'b???????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4789_ = b[2703:2688];
      256'b??????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4789_ = b[2719:2704];
      256'b?????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4789_ = b[2735:2720];
      256'b????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4789_ = b[2751:2736];
      256'b???????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4789_ = b[2767:2752];
      256'b??????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4789_ = b[2783:2768];
      256'b?????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4789_ = b[2799:2784];
      256'b????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4789_ = b[2815:2800];
      256'b???????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4789_ = b[2831:2816];
      256'b??????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4789_ = b[2847:2832];
      256'b?????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4789_ = b[2863:2848];
      256'b????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4789_ = b[2879:2864];
      256'b???????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4789_ = b[2895:2880];
      256'b??????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4789_ = b[2911:2896];
      256'b?????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4789_ = b[2927:2912];
      256'b????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4789_ = b[2943:2928];
      256'b???????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4789_ = b[2959:2944];
      256'b??????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4789_ = b[2975:2960];
      256'b?????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4789_ = b[2991:2976];
      256'b????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4789_ = b[3007:2992];
      256'b???????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4789_ = b[3023:3008];
      256'b??????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4789_ = b[3039:3024];
      256'b?????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4789_ = b[3055:3040];
      256'b????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4789_ = b[3071:3056];
      256'b???????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4789_ = b[3087:3072];
      256'b??????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4789_ = b[3103:3088];
      256'b?????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4789_ = b[3119:3104];
      256'b????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4789_ = b[3135:3120];
      256'b???????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4789_ = b[3151:3136];
      256'b??????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4789_ = b[3167:3152];
      256'b?????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4789_ = b[3183:3168];
      256'b????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4789_ = b[3199:3184];
      256'b???????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4789_ = b[3215:3200];
      256'b??????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4789_ = b[3231:3216];
      256'b?????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4789_ = b[3247:3232];
      256'b????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4789_ = b[3263:3248];
      256'b???????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4789_ = b[3279:3264];
      256'b??????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4789_ = b[3295:3280];
      256'b?????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4789_ = b[3311:3296];
      256'b????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4789_ = b[3327:3312];
      256'b???????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4789_ = b[3343:3328];
      256'b??????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4789_ = b[3359:3344];
      256'b?????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4789_ = b[3375:3360];
      256'b????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4789_ = b[3391:3376];
      256'b???????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4789_ = b[3407:3392];
      256'b??????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4789_ = b[3423:3408];
      256'b?????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4789_ = b[3439:3424];
      256'b????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4789_ = b[3455:3440];
      256'b???????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4789_ = b[3471:3456];
      256'b??????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4789_ = b[3487:3472];
      256'b?????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4789_ = b[3503:3488];
      256'b????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4789_ = b[3519:3504];
      256'b???????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4789_ = b[3535:3520];
      256'b??????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4789_ = b[3551:3536];
      256'b?????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4789_ = b[3567:3552];
      256'b????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4789_ = b[3583:3568];
      256'b???????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4789_ = b[3599:3584];
      256'b??????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4789_ = b[3615:3600];
      256'b?????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4789_ = b[3631:3616];
      256'b????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4789_ = b[3647:3632];
      256'b???????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4789_ = b[3663:3648];
      256'b??????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4789_ = b[3679:3664];
      256'b?????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4789_ = b[3695:3680];
      256'b????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4789_ = b[3711:3696];
      256'b???????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4789_ = b[3727:3712];
      256'b??????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4789_ = b[3743:3728];
      256'b?????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4789_ = b[3759:3744];
      256'b????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4789_ = b[3775:3760];
      256'b???????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4789_ = b[3791:3776];
      256'b??????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4789_ = b[3807:3792];
      256'b?????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4789_ = b[3823:3808];
      256'b????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4789_ = b[3839:3824];
      256'b???????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4789_ = b[3855:3840];
      256'b??????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4789_ = b[3871:3856];
      256'b?????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4789_ = b[3887:3872];
      256'b????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4789_ = b[3903:3888];
      256'b???????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4789_ = b[3919:3904];
      256'b??????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4789_ = b[3935:3920];
      256'b?????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4789_ = b[3951:3936];
      256'b????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4789_ = b[3967:3952];
      256'b???????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4789_ = b[3983:3968];
      256'b??????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4789_ = b[3999:3984];
      256'b?????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4789_ = b[4015:4000];
      256'b????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4789_ = b[4031:4016];
      256'b???1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4789_ = b[4047:4032];
      256'b??1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4789_ = b[4063:4048];
      256'b?1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4789_ = b[4079:4064];
      256'b1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _4789_ = b[4095:4080];
      default:
        _4789_ = a;
    endcase
  endfunction
  assign _0944_ = _4789_(density_reg0, { density_reg1, density_reg2, density_reg3, density_reg4, density_reg5, density_reg6, density_reg7, density_reg8, density_reg9, density_reg10, density_reg11, density_reg12, density_reg13, density_reg14, density_reg15, density_reg16, density_reg17, density_reg18, density_reg19, density_reg20, density_reg21, density_reg22, density_reg23, density_reg24, density_reg25, density_reg26, density_reg27, density_reg28, density_reg29, density_reg30, density_reg31, density_reg32, density_reg33, density_reg34, density_reg35, density_reg36, density_reg37, density_reg38, density_reg39, density_reg40, density_reg41, density_reg42, density_reg43, density_reg44, density_reg45, density_reg46, density_reg47, density_reg48, density_reg49, density_reg50, density_reg51, density_reg52, density_reg53, density_reg54, density_reg55, density_reg56, density_reg57, density_reg58, density_reg59, density_reg60, density_reg61, density_reg62, density_reg63, density_reg64, density_reg65, density_reg66, density_reg67, density_reg68, density_reg69, density_reg70, density_reg71, density_reg72, density_reg73, density_reg74, density_reg75, density_reg76, density_reg77, density_reg78, density_reg79, density_reg80, density_reg81, density_reg82, density_reg83, density_reg84, density_reg85, density_reg86, density_reg87, density_reg88, density_reg89, density_reg90, density_reg91, density_reg92, density_reg93, density_reg94, density_reg95, density_reg96, density_reg97, density_reg98, density_reg99, density_reg100, density_reg101, density_reg102, density_reg103, density_reg104, density_reg105, density_reg106, density_reg107, density_reg108, density_reg109, density_reg110, density_reg111, density_reg112, density_reg113, density_reg114, density_reg115, density_reg116, density_reg117, density_reg118, density_reg119, density_reg120, density_reg121, density_reg122, density_reg123, density_reg124, density_reg125, density_reg126, density_reg127, density_reg128, density_reg129, density_reg130, density_reg131, density_reg132, density_reg133, density_reg134, density_reg135, density_reg136, density_reg137, density_reg138, density_reg139, density_reg140, density_reg141, density_reg142, density_reg143, density_reg144, density_reg145, density_reg146, density_reg147, density_reg148, density_reg149, density_reg150, density_reg151, density_reg152, density_reg153, density_reg154, density_reg155, density_reg156, density_reg157, density_reg158, density_reg159, density_reg160, density_reg161, density_reg162, density_reg163, density_reg164, density_reg165, density_reg166, density_reg167, density_reg168, density_reg169, density_reg170, density_reg171, density_reg172, density_reg173, density_reg174, density_reg175, density_reg176, density_reg177, density_reg178, density_reg179, density_reg180, density_reg181, density_reg182, density_reg183, density_reg184, density_reg185, density_reg186, density_reg187, density_reg188, density_reg189, density_reg190, density_reg191, density_reg192, density_reg193, density_reg194, density_reg195, density_reg196, density_reg197, density_reg198, density_reg199, density_reg200, density_reg201, density_reg202, density_reg203, density_reg204, density_reg205, density_reg206, density_reg207, density_reg208, density_reg209, density_reg210, density_reg211, density_reg212, density_reg213, density_reg214, density_reg215, density_reg216, density_reg217, density_reg218, density_reg219, density_reg220, density_reg221, density_reg222, density_reg223, density_reg224, density_reg225, density_reg226, density_reg227, density_reg228, density_reg229, density_reg230, density_reg231, density_reg232, density_reg233, density_reg234, density_reg235, density_reg236, density_reg237, density_reg238, density_reg239, density_reg240, density_reg241, density_reg242, density_reg243, density_reg244, density_reg245, density_reg246, density_reg247, density_reg248, density_reg249, density_reg250, density_reg251, density_reg252, density_reg253, density_reg254, density_reg255, density_reg256 }, { _1201_, _1200_, _1199_, _1198_, _1197_, _1196_, _1195_, _1194_, _1193_, _1192_, _1191_, _1190_, _1189_, _1188_, _1187_, _1186_, _1185_, _1184_, _1183_, _1182_, _1181_, _1180_, _1179_, _1178_, _1177_, _1176_, _1175_, _1174_, _1173_, _1172_, _1171_, _1170_, _1169_, _1168_, _1167_, _1166_, _1165_, _1164_, _1163_, _1162_, _1161_, _1160_, _1159_, _1158_, _1157_, _1156_, _1155_, _1154_, _1153_, _1152_, _1151_, _1150_, _1149_, _1148_, _1147_, _1146_, _1145_, _1144_, _1143_, _1142_, _1141_, _1140_, _1139_, _1138_, _1137_, _1136_, _1135_, _1134_, _1133_, _1132_, _1131_, _1130_, _1129_, _1128_, _1127_, _1126_, _1125_, _1124_, _1123_, _1122_, _1121_, _1120_, _1119_, _1118_, _1117_, _1116_, _1115_, _1114_, _1113_, _1112_, _1111_, _1110_, _1109_, _1108_, _1107_, _1106_, _1105_, _1104_, _1103_, _1102_, _1101_, _1100_, _1099_, _1098_, _1097_, _1096_, _1095_, _1094_, _1093_, _1092_, _1091_, _1090_, _1089_, _1088_, _1087_, _1086_, _1085_, _1084_, _1083_, _1082_, _1081_, _1080_, _1079_, _1078_, _1077_, _1076_, _1075_, _1074_, _1073_, _1072_, _1071_, _1070_, _1069_, _1068_, _1067_, _1066_, _1065_, _1064_, _1063_, _1062_, _1061_, _1060_, _1059_, _1058_, _1057_, _1056_, _1055_, _1054_, _1053_, _1052_, _1051_, _1050_, _1049_, _1048_, _1047_, _1046_, _1045_, _1044_, _1043_, _1042_, _1041_, _1040_, _1039_, _1038_, _1037_, _1036_, _1035_, _1034_, _1033_, _1032_, _1031_, _1030_, _1029_, _1028_, _1027_, _1026_, _1025_, _1024_, _1023_, _1022_, _1021_, _1020_, _1019_, _1018_, _1017_, _1016_, _1015_, _1014_, _1013_, _1012_, _1011_, _1010_, _1009_, _1008_, _1007_, _1006_, _1005_, _1004_, _1003_, _1002_, _1001_, _1000_, _0999_, _0998_, _0997_, _0996_, _0995_, _0994_, _0993_, _0992_, _0991_, _0990_, _0989_, _0988_, _0987_, _0986_, _0985_, _0984_, _0983_, _0982_, _0981_, _0980_, _0979_, _0978_, _0977_, _0976_, _0975_, _0974_, _0973_, _0972_, _0971_, _0970_, _0969_, _0968_, _0967_, _0966_, _0965_, _0964_, _0963_, _0962_, _0961_, _0960_, _0959_, _0958_, _0957_, _0956_, _0955_, _0954_, _0953_, _0952_, _0951_, _0950_, _0949_, _0948_, _0947_, _0403_ });
  assign _0945_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14554|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 9'b100000000;
  assign _0946_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14550|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 8'b11111111;
  assign _0947_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14546|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 8'b11111110;
  assign _0948_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14542|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 8'b11111101;
  assign _0949_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14538|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 8'b11111100;
  assign _0950_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14534|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 8'b11111011;
  assign _0951_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14530|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 8'b11111010;
  assign _0952_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14526|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 8'b11111001;
  assign _0953_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14522|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 8'b11111000;
  assign _0954_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14518|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 8'b11110111;
  assign _0955_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14514|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 8'b11110110;
  assign _0956_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14510|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 8'b11110101;
  assign _0957_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14506|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 8'b11110100;
  assign _0958_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14502|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 8'b11110011;
  assign _0959_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14498|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 8'b11110010;
  assign _0960_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14494|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 8'b11110001;
  assign _0961_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14490|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 8'b11110000;
  assign _0962_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14486|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 8'b11101111;
  assign _0963_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14482|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 8'b11101110;
  assign _0964_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14478|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 8'b11101101;
  assign _0965_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14474|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 8'b11101100;
  assign _0966_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14470|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 8'b11101011;
  assign _0967_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14466|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 8'b11101010;
  assign _0968_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14462|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 8'b11101001;
  assign _0969_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14458|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 8'b11101000;
  assign _0970_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14454|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 8'b11100111;
  assign _0971_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14450|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 8'b11100110;
  assign _0972_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14446|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 8'b11100101;
  assign _0973_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14442|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 8'b11100100;
  assign _0974_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14438|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 8'b11100011;
  assign _0975_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14434|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 8'b11100010;
  assign _0976_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14430|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 8'b11100001;
  assign _0977_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14426|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 8'b11100000;
  assign _0978_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14422|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 8'b11011111;
  assign _0979_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14418|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 8'b11011110;
  assign _0980_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14414|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 8'b11011101;
  assign _0981_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14410|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 8'b11011100;
  assign _0982_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14406|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 8'b11011011;
  assign _0983_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14402|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 8'b11011010;
  assign _0984_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14398|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 8'b11011001;
  assign _0985_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14394|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 8'b11011000;
  assign _0986_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14390|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 8'b11010111;
  assign _0987_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14386|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 8'b11010110;
  assign _0988_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14382|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 8'b11010101;
  assign _0989_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14378|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 8'b11010100;
  assign _0990_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14374|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 8'b11010011;
  assign _0991_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14370|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 8'b11010010;
  assign _0992_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14366|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 8'b11010001;
  assign _0993_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14362|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 8'b11010000;
  assign _0994_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14358|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 8'b11001111;
  assign _0995_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14354|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 8'b11001110;
  assign _0996_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14350|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 8'b11001101;
  assign _0997_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14346|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 8'b11001100;
  assign _0998_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14342|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 8'b11001011;
  assign _0999_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14338|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 8'b11001010;
  assign _1000_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14334|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 8'b11001001;
  assign _1001_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14330|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 8'b11001000;
  assign _1002_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14326|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 8'b11000111;
  assign _1003_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14322|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 8'b11000110;
  assign _1004_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14318|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 8'b11000101;
  assign _1005_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14314|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 8'b11000100;
  assign _1006_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14310|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 8'b11000011;
  assign _1007_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14306|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 8'b11000010;
  assign _1008_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14302|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 8'b11000001;
  assign _1009_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14298|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 8'b11000000;
  assign _1010_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14294|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 8'b10111111;
  assign _1011_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14290|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 8'b10111110;
  assign _1012_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14286|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 8'b10111101;
  assign _1013_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14282|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 8'b10111100;
  assign _1014_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14278|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 8'b10111011;
  assign _1015_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14274|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 8'b10111010;
  assign _1016_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14270|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 8'b10111001;
  assign _1017_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14266|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 8'b10111000;
  assign _1018_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14262|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 8'b10110111;
  assign _1019_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14258|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 8'b10110110;
  assign _1020_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14254|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 8'b10110101;
  assign _1021_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14250|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 8'b10110100;
  assign _1022_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14246|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 8'b10110011;
  assign _1023_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14242|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 8'b10110010;
  assign _1024_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14238|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 8'b10110001;
  assign _1025_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14234|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 8'b10110000;
  assign _1026_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14230|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 8'b10101111;
  assign _1027_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14226|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 8'b10101110;
  assign _1028_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14222|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 8'b10101101;
  assign _1029_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14218|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 8'b10101100;
  assign _1030_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14214|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 8'b10101011;
  assign _1031_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14210|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 8'b10101010;
  assign _1032_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14206|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 8'b10101001;
  assign _1033_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14202|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 8'b10101000;
  assign _1034_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14198|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 8'b10100111;
  assign _1035_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14194|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 8'b10100110;
  assign _1036_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14190|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 8'b10100101;
  assign _1037_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14186|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 8'b10100100;
  assign _1038_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14182|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 8'b10100011;
  assign _1039_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14178|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 8'b10100010;
  assign _1040_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14174|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 8'b10100001;
  assign _1041_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14170|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 8'b10100000;
  assign _1042_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14166|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 8'b10011111;
  assign _1043_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14162|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 8'b10011110;
  assign _1044_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14158|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 8'b10011101;
  assign _1045_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14154|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 8'b10011100;
  assign _1046_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14150|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 8'b10011011;
  assign _1047_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14146|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 8'b10011010;
  assign _1048_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14142|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 8'b10011001;
  assign _1049_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14138|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 8'b10011000;
  assign _1050_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14134|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 8'b10010111;
  assign _1051_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14130|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 8'b10010110;
  assign _1052_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14126|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 8'b10010101;
  assign _1053_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14122|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 8'b10010100;
  assign _1054_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14118|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 8'b10010011;
  assign _1055_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14114|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 8'b10010010;
  assign _1056_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14110|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 8'b10010001;
  assign _1057_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14106|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 8'b10010000;
  assign _1058_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14102|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 8'b10001111;
  assign _1059_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14098|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 8'b10001110;
  assign _1060_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14094|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 8'b10001101;
  assign _1061_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14090|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 8'b10001100;
  assign _1062_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14086|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 8'b10001011;
  assign _1063_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14082|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 8'b10001010;
  assign _1064_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14078|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 8'b10001001;
  assign _1065_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14074|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 8'b10001000;
  assign _1066_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14070|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 8'b10000111;
  assign _1067_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14066|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 8'b10000110;
  assign _1068_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14062|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 8'b10000101;
  assign _1069_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14058|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 8'b10000100;
  assign _1070_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14054|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 8'b10000011;
  assign _1071_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14050|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 8'b10000010;
  assign _1072_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14046|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 8'b10000001;
  assign _1073_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14042|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 8'b10000000;
  assign _1074_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14038|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 7'b1111111;
  assign _1075_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14034|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 7'b1111110;
  assign _1076_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14030|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 7'b1111101;
  assign _1077_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14026|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 7'b1111100;
  assign _1078_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14022|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 7'b1111011;
  assign _1079_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14018|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 7'b1111010;
  assign _1080_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14014|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 7'b1111001;
  assign _1081_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14010|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 7'b1111000;
  assign _1082_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14006|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 7'b1110111;
  assign _1083_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14002|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 7'b1110110;
  assign _1084_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13998|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 7'b1110101;
  assign _1085_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13994|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 7'b1110100;
  assign _1086_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13990|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 7'b1110011;
  assign _1087_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13986|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 7'b1110010;
  assign _1088_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13982|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 7'b1110001;
  assign _1089_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13978|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 7'b1110000;
  assign _1090_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13974|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 7'b1101111;
  assign _1091_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13970|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 7'b1101110;
  assign _1092_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13966|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 7'b1101101;
  assign _1093_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13962|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 7'b1101100;
  assign _1094_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13958|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 7'b1101011;
  assign _1095_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13954|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 7'b1101010;
  assign _1096_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13950|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 7'b1101001;
  assign _1097_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13946|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 7'b1101000;
  assign _1098_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13942|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 7'b1100111;
  assign _1099_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13938|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 7'b1100110;
  assign _1100_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13934|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 7'b1100101;
  assign _1101_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13930|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 7'b1100100;
  assign _1102_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13926|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 7'b1100011;
  assign _1103_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13922|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 7'b1100010;
  assign _1104_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13918|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 7'b1100001;
  assign _1105_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13914|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 7'b1100000;
  assign _1106_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13910|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 7'b1011111;
  assign _1107_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13906|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 7'b1011110;
  assign _1108_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13902|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 7'b1011101;
  assign _1109_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13898|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 7'b1011100;
  assign _1110_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13894|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 7'b1011011;
  assign _1111_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13890|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 7'b1011010;
  assign _1112_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13886|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 7'b1011001;
  assign _1113_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13882|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 7'b1011000;
  assign _1114_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13878|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 7'b1010111;
  assign _1115_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13874|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 7'b1010110;
  assign _1116_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13870|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 7'b1010101;
  assign _1117_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13866|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 7'b1010100;
  assign _1118_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13862|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 7'b1010011;
  assign _1119_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13858|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 7'b1010010;
  assign _1120_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13854|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 7'b1010001;
  assign _1121_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13850|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 7'b1010000;
  assign _1122_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13846|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 7'b1001111;
  assign _1123_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13842|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 7'b1001110;
  assign _1124_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13838|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 7'b1001101;
  assign _1125_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13834|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 7'b1001100;
  assign _1126_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13830|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 7'b1001011;
  assign _1127_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13826|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 7'b1001010;
  assign _1128_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13822|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 7'b1001001;
  assign _1129_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13818|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 7'b1001000;
  assign _1130_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13814|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 7'b1000111;
  assign _1131_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13810|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 7'b1000110;
  assign _1132_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13806|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 7'b1000101;
  assign _1133_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13802|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 7'b1000100;
  assign _1134_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13798|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 7'b1000011;
  assign _1135_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13794|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 7'b1000010;
  assign _1136_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13790|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 7'b1000001;
  assign _1137_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13786|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 7'b1000000;
  assign _1138_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13782|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 6'b111111;
  assign _1139_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13778|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 6'b111110;
  assign _1140_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13774|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 6'b111101;
  assign _1141_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13770|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 6'b111100;
  assign _1142_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13766|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 6'b111011;
  assign _1143_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13762|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 6'b111010;
  assign _1144_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13758|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 6'b111001;
  assign _1145_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13754|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 6'b111000;
  assign _1146_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13750|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 6'b110111;
  assign _1147_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13746|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 6'b110110;
  assign _1148_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13742|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 6'b110101;
  assign _1149_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13738|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 6'b110100;
  assign _1150_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13734|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 6'b110011;
  assign _1151_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13730|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 6'b110010;
  assign _1152_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13726|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 6'b110001;
  assign _1153_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13722|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 6'b110000;
  assign _1154_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13718|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 6'b101111;
  assign _1155_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13714|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 6'b101110;
  assign _1156_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13710|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 6'b101101;
  assign _1157_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13706|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 6'b101100;
  assign _1158_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13702|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 6'b101011;
  assign _1159_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13698|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 6'b101010;
  assign _1160_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13694|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 6'b101001;
  assign _1161_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13690|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 6'b101000;
  assign _1162_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13686|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 6'b100111;
  assign _1163_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13682|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 6'b100110;
  assign _1164_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13678|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 6'b100101;
  assign _1165_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13674|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 6'b100100;
  assign _1166_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13670|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 6'b100011;
  assign _1167_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13666|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 6'b100010;
  assign _1168_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13662|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 6'b100001;
  assign _1169_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13658|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 6'b100000;
  assign _1170_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13654|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 5'b11111;
  assign _1171_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13650|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 5'b11110;
  assign _1172_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13646|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 5'b11101;
  assign _1173_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13642|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 5'b11100;
  assign _1174_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13638|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 5'b11011;
  assign _1175_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13634|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 5'b11010;
  assign _1176_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13630|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 5'b11001;
  assign _1177_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13626|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 5'b11000;
  assign _1178_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13622|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 5'b10111;
  assign _1179_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13618|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 5'b10110;
  assign _1180_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13614|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 5'b10101;
  assign _1181_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13610|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 5'b10100;
  assign _1182_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13606|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 5'b10011;
  assign _1183_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13602|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 5'b10010;
  assign _1184_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13598|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 5'b10001;
  assign _1185_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13594|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 5'b10000;
  assign _1186_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13590|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 4'b1111;
  assign _1187_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13586|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 4'b1110;
  assign _1188_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13582|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 4'b1101;
  assign _1189_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13578|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 4'b1100;
  assign _1190_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13574|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 4'b1011;
  assign _1191_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13570|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 4'b1010;
  assign _1192_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13566|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 4'b1001;
  assign _1193_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13562|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 4'b1000;
  assign _1194_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13558|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 3'b111;
  assign _1195_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13554|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 3'b110;
  assign _1196_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13550|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 3'b101;
  assign _1197_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13546|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 3'b100;
  assign _1198_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13542|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 2'b11;
  assign _1199_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13538|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 2'b10;
  assign _1200_ = dp2lut_Y_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13534|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) 1'b1;
  assign _1201_ = ! (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13530|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *) dp2lut_Y_entry_6;
  assign _1202_ = dp2lut_Yinfo_6[17] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13525" *) density_reg256 : _0944_;
  assign _1203_ = dp2lut_Yinfo_6[16] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13522" *) density_reg0 : _1202_;
  assign _0298_ = _0390_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13521" *) _1203_ : lut_Y_data_61;
  function [15:0] _5050_;
    input [15:0] a;
    input [4095:0] b;
    input [255:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:14554|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13529" *)
    (* parallel_case *)
    casez (s)
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1:
        _5050_ = b[15:0];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?:
        _5050_ = b[31:16];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??:
        _5050_ = b[47:32];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???:
        _5050_ = b[63:48];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????:
        _5050_ = b[79:64];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????:
        _5050_ = b[95:80];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????:
        _5050_ = b[111:96];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????:
        _5050_ = b[127:112];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????:
        _5050_ = b[143:128];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????:
        _5050_ = b[159:144];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????:
        _5050_ = b[175:160];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????:
        _5050_ = b[191:176];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????:
        _5050_ = b[207:192];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????:
        _5050_ = b[223:208];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????:
        _5050_ = b[239:224];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????:
        _5050_ = b[255:240];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????:
        _5050_ = b[271:256];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????:
        _5050_ = b[287:272];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????:
        _5050_ = b[303:288];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????:
        _5050_ = b[319:304];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????:
        _5050_ = b[335:320];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????:
        _5050_ = b[351:336];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????:
        _5050_ = b[367:352];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????:
        _5050_ = b[383:368];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????:
        _5050_ = b[399:384];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????:
        _5050_ = b[415:400];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????:
        _5050_ = b[431:416];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????:
        _5050_ = b[447:432];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????:
        _5050_ = b[463:448];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????:
        _5050_ = b[479:464];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????:
        _5050_ = b[495:480];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????:
        _5050_ = b[511:496];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????:
        _5050_ = b[527:512];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????:
        _5050_ = b[543:528];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????:
        _5050_ = b[559:544];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????:
        _5050_ = b[575:560];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????:
        _5050_ = b[591:576];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????:
        _5050_ = b[607:592];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????:
        _5050_ = b[623:608];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????:
        _5050_ = b[639:624];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????:
        _5050_ = b[655:640];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????:
        _5050_ = b[671:656];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????:
        _5050_ = b[687:672];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????:
        _5050_ = b[703:688];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????:
        _5050_ = b[719:704];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????:
        _5050_ = b[735:720];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????:
        _5050_ = b[751:736];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????:
        _5050_ = b[767:752];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????:
        _5050_ = b[783:768];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????:
        _5050_ = b[799:784];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????:
        _5050_ = b[815:800];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????:
        _5050_ = b[831:816];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????:
        _5050_ = b[847:832];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????:
        _5050_ = b[863:848];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????:
        _5050_ = b[879:864];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????:
        _5050_ = b[895:880];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????:
        _5050_ = b[911:896];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????:
        _5050_ = b[927:912];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????:
        _5050_ = b[943:928];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????:
        _5050_ = b[959:944];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????:
        _5050_ = b[975:960];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????:
        _5050_ = b[991:976];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????:
        _5050_ = b[1007:992];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????:
        _5050_ = b[1023:1008];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????:
        _5050_ = b[1039:1024];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????:
        _5050_ = b[1055:1040];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????:
        _5050_ = b[1071:1056];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????:
        _5050_ = b[1087:1072];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????:
        _5050_ = b[1103:1088];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????:
        _5050_ = b[1119:1104];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????:
        _5050_ = b[1135:1120];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????:
        _5050_ = b[1151:1136];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????:
        _5050_ = b[1167:1152];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????:
        _5050_ = b[1183:1168];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????:
        _5050_ = b[1199:1184];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????:
        _5050_ = b[1215:1200];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????:
        _5050_ = b[1231:1216];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????:
        _5050_ = b[1247:1232];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????:
        _5050_ = b[1263:1248];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????:
        _5050_ = b[1279:1264];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????:
        _5050_ = b[1295:1280];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????:
        _5050_ = b[1311:1296];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????:
        _5050_ = b[1327:1312];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????:
        _5050_ = b[1343:1328];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????:
        _5050_ = b[1359:1344];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????:
        _5050_ = b[1375:1360];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????:
        _5050_ = b[1391:1376];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????:
        _5050_ = b[1407:1392];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????:
        _5050_ = b[1423:1408];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????:
        _5050_ = b[1439:1424];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????:
        _5050_ = b[1455:1440];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????:
        _5050_ = b[1471:1456];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????:
        _5050_ = b[1487:1472];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????:
        _5050_ = b[1503:1488];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????:
        _5050_ = b[1519:1504];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????:
        _5050_ = b[1535:1520];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????:
        _5050_ = b[1551:1536];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????:
        _5050_ = b[1567:1552];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????:
        _5050_ = b[1583:1568];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????:
        _5050_ = b[1599:1584];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5050_ = b[1615:1600];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5050_ = b[1631:1616];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5050_ = b[1647:1632];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5050_ = b[1663:1648];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5050_ = b[1679:1664];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5050_ = b[1695:1680];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5050_ = b[1711:1696];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5050_ = b[1727:1712];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5050_ = b[1743:1728];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5050_ = b[1759:1744];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5050_ = b[1775:1760];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5050_ = b[1791:1776];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5050_ = b[1807:1792];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5050_ = b[1823:1808];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5050_ = b[1839:1824];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5050_ = b[1855:1840];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5050_ = b[1871:1856];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5050_ = b[1887:1872];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5050_ = b[1903:1888];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5050_ = b[1919:1904];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5050_ = b[1935:1920];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5050_ = b[1951:1936];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5050_ = b[1967:1952];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5050_ = b[1983:1968];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5050_ = b[1999:1984];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5050_ = b[2015:2000];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5050_ = b[2031:2016];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5050_ = b[2047:2032];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5050_ = b[2063:2048];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5050_ = b[2079:2064];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5050_ = b[2095:2080];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5050_ = b[2111:2096];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5050_ = b[2127:2112];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5050_ = b[2143:2128];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5050_ = b[2159:2144];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5050_ = b[2175:2160];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5050_ = b[2191:2176];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5050_ = b[2207:2192];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5050_ = b[2223:2208];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5050_ = b[2239:2224];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5050_ = b[2255:2240];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5050_ = b[2271:2256];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5050_ = b[2287:2272];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5050_ = b[2303:2288];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5050_ = b[2319:2304];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5050_ = b[2335:2320];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5050_ = b[2351:2336];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5050_ = b[2367:2352];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5050_ = b[2383:2368];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5050_ = b[2399:2384];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5050_ = b[2415:2400];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5050_ = b[2431:2416];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5050_ = b[2447:2432];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5050_ = b[2463:2448];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5050_ = b[2479:2464];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5050_ = b[2495:2480];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5050_ = b[2511:2496];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5050_ = b[2527:2512];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5050_ = b[2543:2528];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5050_ = b[2559:2544];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5050_ = b[2575:2560];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5050_ = b[2591:2576];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5050_ = b[2607:2592];
      256'b????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5050_ = b[2623:2608];
      256'b???????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5050_ = b[2639:2624];
      256'b??????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5050_ = b[2655:2640];
      256'b?????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5050_ = b[2671:2656];
      256'b????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5050_ = b[2687:2672];
      256'b???????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5050_ = b[2703:2688];
      256'b??????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5050_ = b[2719:2704];
      256'b?????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5050_ = b[2735:2720];
      256'b????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5050_ = b[2751:2736];
      256'b???????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5050_ = b[2767:2752];
      256'b??????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5050_ = b[2783:2768];
      256'b?????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5050_ = b[2799:2784];
      256'b????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5050_ = b[2815:2800];
      256'b???????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5050_ = b[2831:2816];
      256'b??????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5050_ = b[2847:2832];
      256'b?????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5050_ = b[2863:2848];
      256'b????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5050_ = b[2879:2864];
      256'b???????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5050_ = b[2895:2880];
      256'b??????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5050_ = b[2911:2896];
      256'b?????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5050_ = b[2927:2912];
      256'b????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5050_ = b[2943:2928];
      256'b???????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5050_ = b[2959:2944];
      256'b??????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5050_ = b[2975:2960];
      256'b?????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5050_ = b[2991:2976];
      256'b????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5050_ = b[3007:2992];
      256'b???????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5050_ = b[3023:3008];
      256'b??????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5050_ = b[3039:3024];
      256'b?????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5050_ = b[3055:3040];
      256'b????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5050_ = b[3071:3056];
      256'b???????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5050_ = b[3087:3072];
      256'b??????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5050_ = b[3103:3088];
      256'b?????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5050_ = b[3119:3104];
      256'b????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5050_ = b[3135:3120];
      256'b???????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5050_ = b[3151:3136];
      256'b??????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5050_ = b[3167:3152];
      256'b?????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5050_ = b[3183:3168];
      256'b????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5050_ = b[3199:3184];
      256'b???????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5050_ = b[3215:3200];
      256'b??????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5050_ = b[3231:3216];
      256'b?????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5050_ = b[3247:3232];
      256'b????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5050_ = b[3263:3248];
      256'b???????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5050_ = b[3279:3264];
      256'b??????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5050_ = b[3295:3280];
      256'b?????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5050_ = b[3311:3296];
      256'b????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5050_ = b[3327:3312];
      256'b???????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5050_ = b[3343:3328];
      256'b??????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5050_ = b[3359:3344];
      256'b?????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5050_ = b[3375:3360];
      256'b????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5050_ = b[3391:3376];
      256'b???????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5050_ = b[3407:3392];
      256'b??????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5050_ = b[3423:3408];
      256'b?????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5050_ = b[3439:3424];
      256'b????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5050_ = b[3455:3440];
      256'b???????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5050_ = b[3471:3456];
      256'b??????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5050_ = b[3487:3472];
      256'b?????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5050_ = b[3503:3488];
      256'b????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5050_ = b[3519:3504];
      256'b???????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5050_ = b[3535:3520];
      256'b??????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5050_ = b[3551:3536];
      256'b?????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5050_ = b[3567:3552];
      256'b????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5050_ = b[3583:3568];
      256'b???????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5050_ = b[3599:3584];
      256'b??????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5050_ = b[3615:3600];
      256'b?????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5050_ = b[3631:3616];
      256'b????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5050_ = b[3647:3632];
      256'b???????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5050_ = b[3663:3648];
      256'b??????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5050_ = b[3679:3664];
      256'b?????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5050_ = b[3695:3680];
      256'b????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5050_ = b[3711:3696];
      256'b???????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5050_ = b[3727:3712];
      256'b??????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5050_ = b[3743:3728];
      256'b?????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5050_ = b[3759:3744];
      256'b????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5050_ = b[3775:3760];
      256'b???????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5050_ = b[3791:3776];
      256'b??????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5050_ = b[3807:3792];
      256'b?????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5050_ = b[3823:3808];
      256'b????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5050_ = b[3839:3824];
      256'b???????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5050_ = b[3855:3840];
      256'b??????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5050_ = b[3871:3856];
      256'b?????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5050_ = b[3887:3872];
      256'b????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5050_ = b[3903:3888];
      256'b???????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5050_ = b[3919:3904];
      256'b??????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5050_ = b[3935:3920];
      256'b?????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5050_ = b[3951:3936];
      256'b????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5050_ = b[3967:3952];
      256'b???????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5050_ = b[3983:3968];
      256'b??????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5050_ = b[3999:3984];
      256'b?????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5050_ = b[4015:4000];
      256'b????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5050_ = b[4031:4016];
      256'b???1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5050_ = b[4047:4032];
      256'b??1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5050_ = b[4063:4048];
      256'b?1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5050_ = b[4079:4064];
      256'b1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5050_ = b[4095:4080];
      default:
        _5050_ = a;
    endcase
  endfunction
  assign _1204_ = _5050_(density_reg0, { density_reg1, density_reg2, density_reg3, density_reg4, density_reg5, density_reg6, density_reg7, density_reg8, density_reg9, density_reg10, density_reg11, density_reg12, density_reg13, density_reg14, density_reg15, density_reg16, density_reg17, density_reg18, density_reg19, density_reg20, density_reg21, density_reg22, density_reg23, density_reg24, density_reg25, density_reg26, density_reg27, density_reg28, density_reg29, density_reg30, density_reg31, density_reg32, density_reg33, density_reg34, density_reg35, density_reg36, density_reg37, density_reg38, density_reg39, density_reg40, density_reg41, density_reg42, density_reg43, density_reg44, density_reg45, density_reg46, density_reg47, density_reg48, density_reg49, density_reg50, density_reg51, density_reg52, density_reg53, density_reg54, density_reg55, density_reg56, density_reg57, density_reg58, density_reg59, density_reg60, density_reg61, density_reg62, density_reg63, density_reg64, density_reg65, density_reg66, density_reg67, density_reg68, density_reg69, density_reg70, density_reg71, density_reg72, density_reg73, density_reg74, density_reg75, density_reg76, density_reg77, density_reg78, density_reg79, density_reg80, density_reg81, density_reg82, density_reg83, density_reg84, density_reg85, density_reg86, density_reg87, density_reg88, density_reg89, density_reg90, density_reg91, density_reg92, density_reg93, density_reg94, density_reg95, density_reg96, density_reg97, density_reg98, density_reg99, density_reg100, density_reg101, density_reg102, density_reg103, density_reg104, density_reg105, density_reg106, density_reg107, density_reg108, density_reg109, density_reg110, density_reg111, density_reg112, density_reg113, density_reg114, density_reg115, density_reg116, density_reg117, density_reg118, density_reg119, density_reg120, density_reg121, density_reg122, density_reg123, density_reg124, density_reg125, density_reg126, density_reg127, density_reg128, density_reg129, density_reg130, density_reg131, density_reg132, density_reg133, density_reg134, density_reg135, density_reg136, density_reg137, density_reg138, density_reg139, density_reg140, density_reg141, density_reg142, density_reg143, density_reg144, density_reg145, density_reg146, density_reg147, density_reg148, density_reg149, density_reg150, density_reg151, density_reg152, density_reg153, density_reg154, density_reg155, density_reg156, density_reg157, density_reg158, density_reg159, density_reg160, density_reg161, density_reg162, density_reg163, density_reg164, density_reg165, density_reg166, density_reg167, density_reg168, density_reg169, density_reg170, density_reg171, density_reg172, density_reg173, density_reg174, density_reg175, density_reg176, density_reg177, density_reg178, density_reg179, density_reg180, density_reg181, density_reg182, density_reg183, density_reg184, density_reg185, density_reg186, density_reg187, density_reg188, density_reg189, density_reg190, density_reg191, density_reg192, density_reg193, density_reg194, density_reg195, density_reg196, density_reg197, density_reg198, density_reg199, density_reg200, density_reg201, density_reg202, density_reg203, density_reg204, density_reg205, density_reg206, density_reg207, density_reg208, density_reg209, density_reg210, density_reg211, density_reg212, density_reg213, density_reg214, density_reg215, density_reg216, density_reg217, density_reg218, density_reg219, density_reg220, density_reg221, density_reg222, density_reg223, density_reg224, density_reg225, density_reg226, density_reg227, density_reg228, density_reg229, density_reg230, density_reg231, density_reg232, density_reg233, density_reg234, density_reg235, density_reg236, density_reg237, density_reg238, density_reg239, density_reg240, density_reg241, density_reg242, density_reg243, density_reg244, density_reg245, density_reg246, density_reg247, density_reg248, density_reg249, density_reg250, density_reg251, density_reg252, density_reg253, density_reg254, density_reg255, density_reg256 }, { _1200_, _1199_, _1198_, _1197_, _1196_, _1195_, _1194_, _1193_, _1192_, _1191_, _1190_, _1189_, _1188_, _1187_, _1186_, _1185_, _1184_, _1183_, _1182_, _1181_, _1180_, _1179_, _1178_, _1177_, _1176_, _1175_, _1174_, _1173_, _1172_, _1171_, _1170_, _1169_, _1168_, _1167_, _1166_, _1165_, _1164_, _1163_, _1162_, _1161_, _1160_, _1159_, _1158_, _1157_, _1156_, _1155_, _1154_, _1153_, _1152_, _1151_, _1150_, _1149_, _1148_, _1147_, _1146_, _1145_, _1144_, _1143_, _1142_, _1141_, _1140_, _1139_, _1138_, _1137_, _1136_, _1135_, _1134_, _1133_, _1132_, _1131_, _1130_, _1129_, _1128_, _1127_, _1126_, _1125_, _1124_, _1123_, _1122_, _1121_, _1120_, _1119_, _1118_, _1117_, _1116_, _1115_, _1114_, _1113_, _1112_, _1111_, _1110_, _1109_, _1108_, _1107_, _1106_, _1105_, _1104_, _1103_, _1102_, _1101_, _1100_, _1099_, _1098_, _1097_, _1096_, _1095_, _1094_, _1093_, _1092_, _1091_, _1090_, _1089_, _1088_, _1087_, _1086_, _1085_, _1084_, _1083_, _1082_, _1081_, _1080_, _1079_, _1078_, _1077_, _1076_, _1075_, _1074_, _1073_, _1072_, _1071_, _1070_, _1069_, _1068_, _1067_, _1066_, _1065_, _1064_, _1063_, _1062_, _1061_, _1060_, _1059_, _1058_, _1057_, _1056_, _1055_, _1054_, _1053_, _1052_, _1051_, _1050_, _1049_, _1048_, _1047_, _1046_, _1045_, _1044_, _1043_, _1042_, _1041_, _1040_, _1039_, _1038_, _1037_, _1036_, _1035_, _1034_, _1033_, _1032_, _1031_, _1030_, _1029_, _1028_, _1027_, _1026_, _1025_, _1024_, _1023_, _1022_, _1021_, _1020_, _1019_, _1018_, _1017_, _1016_, _1015_, _1014_, _1013_, _1012_, _1011_, _1010_, _1009_, _1008_, _1007_, _1006_, _1005_, _1004_, _1003_, _1002_, _1001_, _1000_, _0999_, _0998_, _0997_, _0996_, _0995_, _0994_, _0993_, _0992_, _0991_, _0990_, _0989_, _0988_, _0987_, _0986_, _0985_, _0984_, _0983_, _0982_, _0981_, _0980_, _0979_, _0978_, _0977_, _0976_, _0975_, _0974_, _0973_, _0972_, _0971_, _0970_, _0969_, _0968_, _0967_, _0966_, _0965_, _0964_, _0963_, _0962_, _0961_, _0960_, _0959_, _0958_, _0957_, _0956_, _0955_, _0954_, _0953_, _0952_, _0951_, _0950_, _0949_, _0948_, _0947_, _0946_, _0945_ });
  assign _1205_ = dp2lut_Yinfo_6[17] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13525" *) density_reg256 : _1204_;
  assign _1206_ = dp2lut_Yinfo_6[16] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13522" *) density_reg0 : _1205_;
  assign _0297_ = _0390_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13521" *) _1206_ : lut_Y_data_60;
  function [15:0] _5054_;
    input [15:0] a;
    input [4095:0] b;
    input [255:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13503|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *)
    (* parallel_case *)
    casez (s)
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1:
        _5054_ = b[15:0];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?:
        _5054_ = b[31:16];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??:
        _5054_ = b[47:32];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???:
        _5054_ = b[63:48];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????:
        _5054_ = b[79:64];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????:
        _5054_ = b[95:80];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????:
        _5054_ = b[111:96];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????:
        _5054_ = b[127:112];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????:
        _5054_ = b[143:128];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????:
        _5054_ = b[159:144];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????:
        _5054_ = b[175:160];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????:
        _5054_ = b[191:176];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????:
        _5054_ = b[207:192];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????:
        _5054_ = b[223:208];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????:
        _5054_ = b[239:224];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????:
        _5054_ = b[255:240];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????:
        _5054_ = b[271:256];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????:
        _5054_ = b[287:272];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????:
        _5054_ = b[303:288];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????:
        _5054_ = b[319:304];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????:
        _5054_ = b[335:320];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????:
        _5054_ = b[351:336];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????:
        _5054_ = b[367:352];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????:
        _5054_ = b[383:368];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????:
        _5054_ = b[399:384];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????:
        _5054_ = b[415:400];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????:
        _5054_ = b[431:416];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????:
        _5054_ = b[447:432];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????:
        _5054_ = b[463:448];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????:
        _5054_ = b[479:464];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????:
        _5054_ = b[495:480];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????:
        _5054_ = b[511:496];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????:
        _5054_ = b[527:512];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????:
        _5054_ = b[543:528];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????:
        _5054_ = b[559:544];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????:
        _5054_ = b[575:560];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????:
        _5054_ = b[591:576];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????:
        _5054_ = b[607:592];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????:
        _5054_ = b[623:608];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????:
        _5054_ = b[639:624];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????:
        _5054_ = b[655:640];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????:
        _5054_ = b[671:656];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????:
        _5054_ = b[687:672];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????:
        _5054_ = b[703:688];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????:
        _5054_ = b[719:704];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????:
        _5054_ = b[735:720];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????:
        _5054_ = b[751:736];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????:
        _5054_ = b[767:752];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????:
        _5054_ = b[783:768];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????:
        _5054_ = b[799:784];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????:
        _5054_ = b[815:800];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????:
        _5054_ = b[831:816];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????:
        _5054_ = b[847:832];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????:
        _5054_ = b[863:848];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????:
        _5054_ = b[879:864];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????:
        _5054_ = b[895:880];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????:
        _5054_ = b[911:896];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????:
        _5054_ = b[927:912];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????:
        _5054_ = b[943:928];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????:
        _5054_ = b[959:944];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????:
        _5054_ = b[975:960];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????:
        _5054_ = b[991:976];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????:
        _5054_ = b[1007:992];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????:
        _5054_ = b[1023:1008];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????:
        _5054_ = b[1039:1024];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????:
        _5054_ = b[1055:1040];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????:
        _5054_ = b[1071:1056];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????:
        _5054_ = b[1087:1072];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????:
        _5054_ = b[1103:1088];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????:
        _5054_ = b[1119:1104];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????:
        _5054_ = b[1135:1120];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????:
        _5054_ = b[1151:1136];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????:
        _5054_ = b[1167:1152];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????:
        _5054_ = b[1183:1168];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????:
        _5054_ = b[1199:1184];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????:
        _5054_ = b[1215:1200];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????:
        _5054_ = b[1231:1216];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????:
        _5054_ = b[1247:1232];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????:
        _5054_ = b[1263:1248];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????:
        _5054_ = b[1279:1264];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????:
        _5054_ = b[1295:1280];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????:
        _5054_ = b[1311:1296];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????:
        _5054_ = b[1327:1312];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????:
        _5054_ = b[1343:1328];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????:
        _5054_ = b[1359:1344];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????:
        _5054_ = b[1375:1360];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????:
        _5054_ = b[1391:1376];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????:
        _5054_ = b[1407:1392];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????:
        _5054_ = b[1423:1408];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????:
        _5054_ = b[1439:1424];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????:
        _5054_ = b[1455:1440];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????:
        _5054_ = b[1471:1456];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????:
        _5054_ = b[1487:1472];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????:
        _5054_ = b[1503:1488];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????:
        _5054_ = b[1519:1504];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????:
        _5054_ = b[1535:1520];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????:
        _5054_ = b[1551:1536];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????:
        _5054_ = b[1567:1552];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????:
        _5054_ = b[1583:1568];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????:
        _5054_ = b[1599:1584];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5054_ = b[1615:1600];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5054_ = b[1631:1616];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5054_ = b[1647:1632];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5054_ = b[1663:1648];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5054_ = b[1679:1664];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5054_ = b[1695:1680];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5054_ = b[1711:1696];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5054_ = b[1727:1712];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5054_ = b[1743:1728];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5054_ = b[1759:1744];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5054_ = b[1775:1760];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5054_ = b[1791:1776];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5054_ = b[1807:1792];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5054_ = b[1823:1808];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5054_ = b[1839:1824];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5054_ = b[1855:1840];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5054_ = b[1871:1856];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5054_ = b[1887:1872];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5054_ = b[1903:1888];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5054_ = b[1919:1904];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5054_ = b[1935:1920];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5054_ = b[1951:1936];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5054_ = b[1967:1952];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5054_ = b[1983:1968];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5054_ = b[1999:1984];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5054_ = b[2015:2000];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5054_ = b[2031:2016];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5054_ = b[2047:2032];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5054_ = b[2063:2048];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5054_ = b[2079:2064];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5054_ = b[2095:2080];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5054_ = b[2111:2096];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5054_ = b[2127:2112];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5054_ = b[2143:2128];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5054_ = b[2159:2144];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5054_ = b[2175:2160];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5054_ = b[2191:2176];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5054_ = b[2207:2192];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5054_ = b[2223:2208];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5054_ = b[2239:2224];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5054_ = b[2255:2240];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5054_ = b[2271:2256];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5054_ = b[2287:2272];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5054_ = b[2303:2288];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5054_ = b[2319:2304];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5054_ = b[2335:2320];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5054_ = b[2351:2336];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5054_ = b[2367:2352];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5054_ = b[2383:2368];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5054_ = b[2399:2384];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5054_ = b[2415:2400];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5054_ = b[2431:2416];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5054_ = b[2447:2432];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5054_ = b[2463:2448];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5054_ = b[2479:2464];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5054_ = b[2495:2480];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5054_ = b[2511:2496];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5054_ = b[2527:2512];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5054_ = b[2543:2528];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5054_ = b[2559:2544];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5054_ = b[2575:2560];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5054_ = b[2591:2576];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5054_ = b[2607:2592];
      256'b????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5054_ = b[2623:2608];
      256'b???????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5054_ = b[2639:2624];
      256'b??????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5054_ = b[2655:2640];
      256'b?????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5054_ = b[2671:2656];
      256'b????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5054_ = b[2687:2672];
      256'b???????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5054_ = b[2703:2688];
      256'b??????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5054_ = b[2719:2704];
      256'b?????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5054_ = b[2735:2720];
      256'b????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5054_ = b[2751:2736];
      256'b???????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5054_ = b[2767:2752];
      256'b??????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5054_ = b[2783:2768];
      256'b?????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5054_ = b[2799:2784];
      256'b????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5054_ = b[2815:2800];
      256'b???????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5054_ = b[2831:2816];
      256'b??????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5054_ = b[2847:2832];
      256'b?????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5054_ = b[2863:2848];
      256'b????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5054_ = b[2879:2864];
      256'b???????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5054_ = b[2895:2880];
      256'b??????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5054_ = b[2911:2896];
      256'b?????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5054_ = b[2927:2912];
      256'b????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5054_ = b[2943:2928];
      256'b???????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5054_ = b[2959:2944];
      256'b??????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5054_ = b[2975:2960];
      256'b?????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5054_ = b[2991:2976];
      256'b????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5054_ = b[3007:2992];
      256'b???????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5054_ = b[3023:3008];
      256'b??????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5054_ = b[3039:3024];
      256'b?????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5054_ = b[3055:3040];
      256'b????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5054_ = b[3071:3056];
      256'b???????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5054_ = b[3087:3072];
      256'b??????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5054_ = b[3103:3088];
      256'b?????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5054_ = b[3119:3104];
      256'b????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5054_ = b[3135:3120];
      256'b???????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5054_ = b[3151:3136];
      256'b??????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5054_ = b[3167:3152];
      256'b?????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5054_ = b[3183:3168];
      256'b????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5054_ = b[3199:3184];
      256'b???????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5054_ = b[3215:3200];
      256'b??????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5054_ = b[3231:3216];
      256'b?????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5054_ = b[3247:3232];
      256'b????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5054_ = b[3263:3248];
      256'b???????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5054_ = b[3279:3264];
      256'b??????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5054_ = b[3295:3280];
      256'b?????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5054_ = b[3311:3296];
      256'b????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5054_ = b[3327:3312];
      256'b???????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5054_ = b[3343:3328];
      256'b??????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5054_ = b[3359:3344];
      256'b?????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5054_ = b[3375:3360];
      256'b????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5054_ = b[3391:3376];
      256'b???????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5054_ = b[3407:3392];
      256'b??????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5054_ = b[3423:3408];
      256'b?????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5054_ = b[3439:3424];
      256'b????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5054_ = b[3455:3440];
      256'b???????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5054_ = b[3471:3456];
      256'b??????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5054_ = b[3487:3472];
      256'b?????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5054_ = b[3503:3488];
      256'b????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5054_ = b[3519:3504];
      256'b???????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5054_ = b[3535:3520];
      256'b??????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5054_ = b[3551:3536];
      256'b?????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5054_ = b[3567:3552];
      256'b????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5054_ = b[3583:3568];
      256'b???????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5054_ = b[3599:3584];
      256'b??????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5054_ = b[3615:3600];
      256'b?????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5054_ = b[3631:3616];
      256'b????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5054_ = b[3647:3632];
      256'b???????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5054_ = b[3663:3648];
      256'b??????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5054_ = b[3679:3664];
      256'b?????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5054_ = b[3695:3680];
      256'b????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5054_ = b[3711:3696];
      256'b???????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5054_ = b[3727:3712];
      256'b??????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5054_ = b[3743:3728];
      256'b?????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5054_ = b[3759:3744];
      256'b????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5054_ = b[3775:3760];
      256'b???????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5054_ = b[3791:3776];
      256'b??????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5054_ = b[3807:3792];
      256'b?????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5054_ = b[3823:3808];
      256'b????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5054_ = b[3839:3824];
      256'b???????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5054_ = b[3855:3840];
      256'b??????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5054_ = b[3871:3856];
      256'b?????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5054_ = b[3887:3872];
      256'b????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5054_ = b[3903:3888];
      256'b???????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5054_ = b[3919:3904];
      256'b??????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5054_ = b[3935:3920];
      256'b?????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5054_ = b[3951:3936];
      256'b????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5054_ = b[3967:3952];
      256'b???????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5054_ = b[3983:3968];
      256'b??????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5054_ = b[3999:3984];
      256'b?????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5054_ = b[4015:4000];
      256'b????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5054_ = b[4031:4016];
      256'b???1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5054_ = b[4047:4032];
      256'b??1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5054_ = b[4063:4048];
      256'b?1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5054_ = b[4079:4064];
      256'b1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5054_ = b[4095:4080];
      default:
        _5054_ = a;
    endcase
  endfunction
  assign _1207_ = _5054_(density_reg0, { density_reg1, density_reg2, density_reg3, density_reg4, density_reg5, density_reg6, density_reg7, density_reg8, density_reg9, density_reg10, density_reg11, density_reg12, density_reg13, density_reg14, density_reg15, density_reg16, density_reg17, density_reg18, density_reg19, density_reg20, density_reg21, density_reg22, density_reg23, density_reg24, density_reg25, density_reg26, density_reg27, density_reg28, density_reg29, density_reg30, density_reg31, density_reg32, density_reg33, density_reg34, density_reg35, density_reg36, density_reg37, density_reg38, density_reg39, density_reg40, density_reg41, density_reg42, density_reg43, density_reg44, density_reg45, density_reg46, density_reg47, density_reg48, density_reg49, density_reg50, density_reg51, density_reg52, density_reg53, density_reg54, density_reg55, density_reg56, density_reg57, density_reg58, density_reg59, density_reg60, density_reg61, density_reg62, density_reg63, density_reg64, density_reg65, density_reg66, density_reg67, density_reg68, density_reg69, density_reg70, density_reg71, density_reg72, density_reg73, density_reg74, density_reg75, density_reg76, density_reg77, density_reg78, density_reg79, density_reg80, density_reg81, density_reg82, density_reg83, density_reg84, density_reg85, density_reg86, density_reg87, density_reg88, density_reg89, density_reg90, density_reg91, density_reg92, density_reg93, density_reg94, density_reg95, density_reg96, density_reg97, density_reg98, density_reg99, density_reg100, density_reg101, density_reg102, density_reg103, density_reg104, density_reg105, density_reg106, density_reg107, density_reg108, density_reg109, density_reg110, density_reg111, density_reg112, density_reg113, density_reg114, density_reg115, density_reg116, density_reg117, density_reg118, density_reg119, density_reg120, density_reg121, density_reg122, density_reg123, density_reg124, density_reg125, density_reg126, density_reg127, density_reg128, density_reg129, density_reg130, density_reg131, density_reg132, density_reg133, density_reg134, density_reg135, density_reg136, density_reg137, density_reg138, density_reg139, density_reg140, density_reg141, density_reg142, density_reg143, density_reg144, density_reg145, density_reg146, density_reg147, density_reg148, density_reg149, density_reg150, density_reg151, density_reg152, density_reg153, density_reg154, density_reg155, density_reg156, density_reg157, density_reg158, density_reg159, density_reg160, density_reg161, density_reg162, density_reg163, density_reg164, density_reg165, density_reg166, density_reg167, density_reg168, density_reg169, density_reg170, density_reg171, density_reg172, density_reg173, density_reg174, density_reg175, density_reg176, density_reg177, density_reg178, density_reg179, density_reg180, density_reg181, density_reg182, density_reg183, density_reg184, density_reg185, density_reg186, density_reg187, density_reg188, density_reg189, density_reg190, density_reg191, density_reg192, density_reg193, density_reg194, density_reg195, density_reg196, density_reg197, density_reg198, density_reg199, density_reg200, density_reg201, density_reg202, density_reg203, density_reg204, density_reg205, density_reg206, density_reg207, density_reg208, density_reg209, density_reg210, density_reg211, density_reg212, density_reg213, density_reg214, density_reg215, density_reg216, density_reg217, density_reg218, density_reg219, density_reg220, density_reg221, density_reg222, density_reg223, density_reg224, density_reg225, density_reg226, density_reg227, density_reg228, density_reg229, density_reg230, density_reg231, density_reg232, density_reg233, density_reg234, density_reg235, density_reg236, density_reg237, density_reg238, density_reg239, density_reg240, density_reg241, density_reg242, density_reg243, density_reg244, density_reg245, density_reg246, density_reg247, density_reg248, density_reg249, density_reg250, density_reg251, density_reg252, density_reg253, density_reg254, density_reg255, density_reg256 }, { _1464_, _1463_, _1462_, _1461_, _1460_, _1459_, _1458_, _1457_, _1456_, _1455_, _1454_, _1453_, _1452_, _1451_, _1450_, _1449_, _1448_, _1447_, _1446_, _1445_, _1444_, _1443_, _1442_, _1441_, _1440_, _1439_, _1438_, _1437_, _1436_, _1435_, _1434_, _1433_, _1432_, _1431_, _1430_, _1429_, _1428_, _1427_, _1426_, _1425_, _1424_, _1423_, _1422_, _1421_, _1420_, _1419_, _1418_, _1417_, _1416_, _1415_, _1414_, _1413_, _1412_, _1411_, _1410_, _1409_, _1408_, _1407_, _1406_, _1405_, _1404_, _1403_, _1402_, _1401_, _1400_, _1399_, _1398_, _1397_, _1396_, _1395_, _1394_, _1393_, _1392_, _1391_, _1390_, _1389_, _1388_, _1387_, _1386_, _1385_, _1384_, _1383_, _1382_, _1381_, _1380_, _1379_, _1378_, _1377_, _1376_, _1375_, _1374_, _1373_, _1372_, _1371_, _1370_, _1369_, _1368_, _1367_, _1366_, _1365_, _1364_, _1363_, _1362_, _1361_, _1360_, _1359_, _1358_, _1357_, _1356_, _1355_, _1354_, _1353_, _1352_, _1351_, _1350_, _1349_, _1348_, _1347_, _1346_, _1345_, _1344_, _1343_, _1342_, _1341_, _1340_, _1339_, _1338_, _1337_, _1336_, _1335_, _1334_, _1333_, _1332_, _1331_, _1330_, _1329_, _1328_, _1327_, _1326_, _1325_, _1324_, _1323_, _1322_, _1321_, _1320_, _1319_, _1318_, _1317_, _1316_, _1315_, _1314_, _1313_, _1312_, _1311_, _1310_, _1309_, _1308_, _1307_, _1306_, _1305_, _1304_, _1303_, _1302_, _1301_, _1300_, _1299_, _1298_, _1297_, _1296_, _1295_, _1294_, _1293_, _1292_, _1291_, _1290_, _1289_, _1288_, _1287_, _1286_, _1285_, _1284_, _1283_, _1282_, _1281_, _1280_, _1279_, _1278_, _1277_, _1276_, _1275_, _1274_, _1273_, _1272_, _1271_, _1270_, _1269_, _1268_, _1267_, _1266_, _1265_, _1264_, _1263_, _1262_, _1261_, _1260_, _1259_, _1258_, _1257_, _1256_, _1255_, _1254_, _1253_, _1252_, _1251_, _1250_, _1249_, _1248_, _1247_, _1246_, _1245_, _1244_, _1243_, _1242_, _1241_, _1240_, _1239_, _1238_, _1237_, _1236_, _1235_, _1234_, _1233_, _1232_, _1231_, _1230_, _1229_, _1228_, _1227_, _1226_, _1225_, _1224_, _1223_, _1222_, _1221_, _1220_, _1219_, _1218_, _1217_, _1216_, _1215_, _1214_, _1213_, _1212_, _1211_, _1210_, _0407_ });
  assign _1208_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13503|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 9'b100000000;
  assign _1209_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13499|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 8'b11111111;
  assign _1210_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13495|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 8'b11111110;
  assign _1211_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13491|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 8'b11111101;
  assign _1212_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13487|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 8'b11111100;
  assign _1213_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13483|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 8'b11111011;
  assign _1214_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13479|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 8'b11111010;
  assign _1215_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13475|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 8'b11111001;
  assign _1216_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13471|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 8'b11111000;
  assign _1217_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13467|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 8'b11110111;
  assign _1218_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13463|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 8'b11110110;
  assign _1219_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13459|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 8'b11110101;
  assign _1220_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13455|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 8'b11110100;
  assign _1221_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13451|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 8'b11110011;
  assign _1222_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13447|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 8'b11110010;
  assign _1223_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13443|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 8'b11110001;
  assign _1224_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13439|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 8'b11110000;
  assign _1225_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13435|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 8'b11101111;
  assign _1226_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13431|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 8'b11101110;
  assign _1227_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13427|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 8'b11101101;
  assign _1228_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13423|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 8'b11101100;
  assign _1229_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13419|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 8'b11101011;
  assign _1230_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13415|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 8'b11101010;
  assign _1231_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13411|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 8'b11101001;
  assign _1232_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13407|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 8'b11101000;
  assign _1233_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13403|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 8'b11100111;
  assign _1234_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13399|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 8'b11100110;
  assign _1235_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13395|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 8'b11100101;
  assign _1236_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13391|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 8'b11100100;
  assign _1237_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13387|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 8'b11100011;
  assign _1238_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13383|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 8'b11100010;
  assign _1239_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13379|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 8'b11100001;
  assign _1240_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13375|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 8'b11100000;
  assign _1241_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13371|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 8'b11011111;
  assign _1242_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13367|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 8'b11011110;
  assign _1243_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13363|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 8'b11011101;
  assign _1244_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13359|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 8'b11011100;
  assign _1245_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13355|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 8'b11011011;
  assign _1246_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13351|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 8'b11011010;
  assign _1247_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13347|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 8'b11011001;
  assign _1248_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13343|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 8'b11011000;
  assign _1249_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13339|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 8'b11010111;
  assign _1250_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13335|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 8'b11010110;
  assign _1251_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13331|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 8'b11010101;
  assign _1252_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13327|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 8'b11010100;
  assign _1253_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13323|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 8'b11010011;
  assign _1254_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13319|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 8'b11010010;
  assign _1255_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13315|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 8'b11010001;
  assign _1256_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13311|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 8'b11010000;
  assign _1257_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13307|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 8'b11001111;
  assign _1258_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13303|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 8'b11001110;
  assign _1259_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13299|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 8'b11001101;
  assign _1260_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13295|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 8'b11001100;
  assign _1261_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13291|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 8'b11001011;
  assign _1262_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13287|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 8'b11001010;
  assign _1263_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13283|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 8'b11001001;
  assign _1264_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13279|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 8'b11001000;
  assign _1265_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13275|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 8'b11000111;
  assign _1266_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13271|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 8'b11000110;
  assign _1267_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13267|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 8'b11000101;
  assign _1268_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13263|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 8'b11000100;
  assign _1269_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13259|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 8'b11000011;
  assign _1270_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13255|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 8'b11000010;
  assign _1271_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13251|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 8'b11000001;
  assign _1272_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13247|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 8'b11000000;
  assign _1273_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13243|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 8'b10111111;
  assign _1274_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13239|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 8'b10111110;
  assign _1275_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13235|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 8'b10111101;
  assign _1276_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13231|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 8'b10111100;
  assign _1277_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13227|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 8'b10111011;
  assign _1278_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13223|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 8'b10111010;
  assign _1279_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13219|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 8'b10111001;
  assign _1280_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13215|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 8'b10111000;
  assign _1281_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13211|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 8'b10110111;
  assign _1282_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13207|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 8'b10110110;
  assign _1283_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13203|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 8'b10110101;
  assign _1284_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13199|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 8'b10110100;
  assign _1285_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13195|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 8'b10110011;
  assign _1286_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13191|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 8'b10110010;
  assign _1287_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13187|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 8'b10110001;
  assign _1288_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13183|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 8'b10110000;
  assign _1289_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13179|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 8'b10101111;
  assign _1290_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13175|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 8'b10101110;
  assign _1291_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13171|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 8'b10101101;
  assign _1292_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13167|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 8'b10101100;
  assign _1293_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13163|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 8'b10101011;
  assign _1294_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13159|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 8'b10101010;
  assign _1295_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13155|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 8'b10101001;
  assign _1296_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13151|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 8'b10101000;
  assign _1297_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13147|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 8'b10100111;
  assign _1298_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13143|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 8'b10100110;
  assign _1299_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13139|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 8'b10100101;
  assign _1300_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13135|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 8'b10100100;
  assign _1301_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13131|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 8'b10100011;
  assign _1302_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13127|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 8'b10100010;
  assign _1303_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13123|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 8'b10100001;
  assign _1304_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13119|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 8'b10100000;
  assign _1305_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13115|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 8'b10011111;
  assign _1306_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13111|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 8'b10011110;
  assign _1307_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13107|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 8'b10011101;
  assign _1308_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13103|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 8'b10011100;
  assign _1309_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13099|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 8'b10011011;
  assign _1310_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13095|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 8'b10011010;
  assign _1311_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13091|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 8'b10011001;
  assign _1312_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13087|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 8'b10011000;
  assign _1313_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13083|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 8'b10010111;
  assign _1314_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13079|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 8'b10010110;
  assign _1315_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13075|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 8'b10010101;
  assign _1316_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13071|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 8'b10010100;
  assign _1317_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13067|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 8'b10010011;
  assign _1318_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13063|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 8'b10010010;
  assign _1319_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13059|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 8'b10010001;
  assign _1320_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13055|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 8'b10010000;
  assign _1321_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13051|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 8'b10001111;
  assign _1322_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13047|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 8'b10001110;
  assign _1323_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13043|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 8'b10001101;
  assign _1324_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13039|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 8'b10001100;
  assign _1325_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13035|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 8'b10001011;
  assign _1326_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13031|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 8'b10001010;
  assign _1327_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13027|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 8'b10001001;
  assign _1328_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13023|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 8'b10001000;
  assign _1329_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13019|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 8'b10000111;
  assign _1330_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13015|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 8'b10000110;
  assign _1331_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13011|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 8'b10000101;
  assign _1332_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13007|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 8'b10000100;
  assign _1333_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13003|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 8'b10000011;
  assign _1334_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12999|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 8'b10000010;
  assign _1335_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12995|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 8'b10000001;
  assign _1336_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12991|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 8'b10000000;
  assign _1337_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12987|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 7'b1111111;
  assign _1338_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12983|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 7'b1111110;
  assign _1339_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12979|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 7'b1111101;
  assign _1340_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12975|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 7'b1111100;
  assign _1341_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12971|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 7'b1111011;
  assign _1342_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12967|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 7'b1111010;
  assign _1343_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12963|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 7'b1111001;
  assign _1344_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12959|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 7'b1111000;
  assign _1345_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12955|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 7'b1110111;
  assign _1346_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12951|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 7'b1110110;
  assign _1347_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12947|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 7'b1110101;
  assign _1348_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12943|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 7'b1110100;
  assign _1349_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12939|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 7'b1110011;
  assign _1350_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12935|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 7'b1110010;
  assign _1351_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12931|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 7'b1110001;
  assign _1352_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12927|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 7'b1110000;
  assign _1353_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12923|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 7'b1101111;
  assign _1354_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12919|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 7'b1101110;
  assign _1355_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12915|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 7'b1101101;
  assign _1356_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12911|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 7'b1101100;
  assign _1357_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12907|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 7'b1101011;
  assign _1358_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12903|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 7'b1101010;
  assign _1359_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12899|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 7'b1101001;
  assign _1360_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12895|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 7'b1101000;
  assign _1361_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12891|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 7'b1100111;
  assign _1362_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12887|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 7'b1100110;
  assign _1363_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12883|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 7'b1100101;
  assign _1364_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12879|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 7'b1100100;
  assign _1365_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12875|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 7'b1100011;
  assign _1366_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12871|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 7'b1100010;
  assign _1367_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12867|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 7'b1100001;
  assign _1368_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12863|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 7'b1100000;
  assign _1369_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12859|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 7'b1011111;
  assign _1370_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12855|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 7'b1011110;
  assign _1371_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12851|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 7'b1011101;
  assign _1372_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12847|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 7'b1011100;
  assign _1373_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12843|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 7'b1011011;
  assign _1374_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12839|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 7'b1011010;
  assign _1375_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12835|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 7'b1011001;
  assign _1376_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12831|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 7'b1011000;
  assign _1377_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12827|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 7'b1010111;
  assign _1378_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12823|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 7'b1010110;
  assign _1379_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12819|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 7'b1010101;
  assign _1380_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12815|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 7'b1010100;
  assign _1381_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12811|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 7'b1010011;
  assign _1382_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12807|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 7'b1010010;
  assign _1383_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12803|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 7'b1010001;
  assign _1384_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12799|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 7'b1010000;
  assign _1385_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12795|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 7'b1001111;
  assign _1386_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12791|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 7'b1001110;
  assign _1387_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12787|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 7'b1001101;
  assign _1388_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12783|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 7'b1001100;
  assign _1389_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12779|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 7'b1001011;
  assign _1390_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12775|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 7'b1001010;
  assign _1391_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12771|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 7'b1001001;
  assign _1392_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12767|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 7'b1001000;
  assign _1393_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12763|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 7'b1000111;
  assign _1394_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12759|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 7'b1000110;
  assign _1395_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12755|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 7'b1000101;
  assign _1396_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12751|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 7'b1000100;
  assign _1397_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12747|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 7'b1000011;
  assign _1398_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12743|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 7'b1000010;
  assign _1399_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12739|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 7'b1000001;
  assign _1400_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12735|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 7'b1000000;
  assign _1401_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12731|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 6'b111111;
  assign _1402_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12727|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 6'b111110;
  assign _1403_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12723|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 6'b111101;
  assign _1404_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12719|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 6'b111100;
  assign _1405_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12715|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 6'b111011;
  assign _1406_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12711|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 6'b111010;
  assign _1407_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12707|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 6'b111001;
  assign _1408_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12703|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 6'b111000;
  assign _1409_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12699|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 6'b110111;
  assign _1410_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12695|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 6'b110110;
  assign _1411_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12691|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 6'b110101;
  assign _1412_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12687|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 6'b110100;
  assign _1413_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12683|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 6'b110011;
  assign _1414_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12679|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 6'b110010;
  assign _1415_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12675|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 6'b110001;
  assign _1416_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12671|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 6'b110000;
  assign _1417_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12667|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 6'b101111;
  assign _1418_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12663|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 6'b101110;
  assign _1419_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12659|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 6'b101101;
  assign _1420_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12655|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 6'b101100;
  assign _1421_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12651|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 6'b101011;
  assign _1422_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12647|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 6'b101010;
  assign _1423_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12643|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 6'b101001;
  assign _1424_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12639|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 6'b101000;
  assign _1425_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12635|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 6'b100111;
  assign _1426_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12631|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 6'b100110;
  assign _1427_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12627|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 6'b100101;
  assign _1428_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12623|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 6'b100100;
  assign _1429_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12619|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 6'b100011;
  assign _1430_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12615|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 6'b100010;
  assign _1431_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12611|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 6'b100001;
  assign _1432_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12607|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 6'b100000;
  assign _1433_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12603|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 5'b11111;
  assign _1434_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12599|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 5'b11110;
  assign _1435_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12595|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 5'b11101;
  assign _1436_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12591|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 5'b11100;
  assign _1437_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12587|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 5'b11011;
  assign _1438_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12583|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 5'b11010;
  assign _1439_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12579|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 5'b11001;
  assign _1440_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12575|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 5'b11000;
  assign _1441_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12571|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 5'b10111;
  assign _1442_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12567|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 5'b10110;
  assign _1443_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12563|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 5'b10101;
  assign _1444_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12559|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 5'b10100;
  assign _1445_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12555|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 5'b10011;
  assign _1446_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12551|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 5'b10010;
  assign _1447_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12547|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 5'b10001;
  assign _1448_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12543|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 5'b10000;
  assign _1449_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12539|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 4'b1111;
  assign _1450_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12535|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 4'b1110;
  assign _1451_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12531|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 4'b1101;
  assign _1452_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12527|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 4'b1100;
  assign _1453_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12523|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 4'b1011;
  assign _1454_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12519|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 4'b1010;
  assign _1455_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12515|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 4'b1001;
  assign _1456_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12511|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 4'b1000;
  assign _1457_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12507|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 3'b111;
  assign _1458_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12503|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 3'b110;
  assign _1459_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12499|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 3'b101;
  assign _1460_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12495|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 3'b100;
  assign _1461_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12491|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 2'b11;
  assign _1462_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12487|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 2'b10;
  assign _1463_ = dp2lut_Y_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12483|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) 1'b1;
  assign _1464_ = ! (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12479|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *) dp2lut_Y_entry_5;
  assign _1465_ = dp2lut_Yinfo_5[17] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12474" *) density_reg256 : _1207_;
  assign _1466_ = dp2lut_Yinfo_5[16] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12471" *) density_reg0 : _1465_;
  assign _0296_ = _0388_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12470" *) _1466_ : lut_Y_data_51;
  function [15:0] _5315_;
    input [15:0] a;
    input [4095:0] b;
    input [255:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:13503|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12478" *)
    (* parallel_case *)
    casez (s)
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1:
        _5315_ = b[15:0];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?:
        _5315_ = b[31:16];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??:
        _5315_ = b[47:32];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???:
        _5315_ = b[63:48];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????:
        _5315_ = b[79:64];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????:
        _5315_ = b[95:80];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????:
        _5315_ = b[111:96];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????:
        _5315_ = b[127:112];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????:
        _5315_ = b[143:128];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????:
        _5315_ = b[159:144];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????:
        _5315_ = b[175:160];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????:
        _5315_ = b[191:176];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????:
        _5315_ = b[207:192];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????:
        _5315_ = b[223:208];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????:
        _5315_ = b[239:224];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????:
        _5315_ = b[255:240];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????:
        _5315_ = b[271:256];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????:
        _5315_ = b[287:272];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????:
        _5315_ = b[303:288];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????:
        _5315_ = b[319:304];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????:
        _5315_ = b[335:320];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????:
        _5315_ = b[351:336];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????:
        _5315_ = b[367:352];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????:
        _5315_ = b[383:368];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????:
        _5315_ = b[399:384];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????:
        _5315_ = b[415:400];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????:
        _5315_ = b[431:416];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????:
        _5315_ = b[447:432];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????:
        _5315_ = b[463:448];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????:
        _5315_ = b[479:464];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????:
        _5315_ = b[495:480];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????:
        _5315_ = b[511:496];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????:
        _5315_ = b[527:512];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????:
        _5315_ = b[543:528];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????:
        _5315_ = b[559:544];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????:
        _5315_ = b[575:560];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????:
        _5315_ = b[591:576];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????:
        _5315_ = b[607:592];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????:
        _5315_ = b[623:608];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????:
        _5315_ = b[639:624];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????:
        _5315_ = b[655:640];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????:
        _5315_ = b[671:656];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????:
        _5315_ = b[687:672];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????:
        _5315_ = b[703:688];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????:
        _5315_ = b[719:704];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????:
        _5315_ = b[735:720];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????:
        _5315_ = b[751:736];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????:
        _5315_ = b[767:752];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????:
        _5315_ = b[783:768];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????:
        _5315_ = b[799:784];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????:
        _5315_ = b[815:800];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????:
        _5315_ = b[831:816];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????:
        _5315_ = b[847:832];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????:
        _5315_ = b[863:848];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????:
        _5315_ = b[879:864];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????:
        _5315_ = b[895:880];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????:
        _5315_ = b[911:896];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????:
        _5315_ = b[927:912];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????:
        _5315_ = b[943:928];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????:
        _5315_ = b[959:944];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????:
        _5315_ = b[975:960];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????:
        _5315_ = b[991:976];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????:
        _5315_ = b[1007:992];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????:
        _5315_ = b[1023:1008];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????:
        _5315_ = b[1039:1024];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????:
        _5315_ = b[1055:1040];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????:
        _5315_ = b[1071:1056];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????:
        _5315_ = b[1087:1072];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????:
        _5315_ = b[1103:1088];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????:
        _5315_ = b[1119:1104];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????:
        _5315_ = b[1135:1120];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????:
        _5315_ = b[1151:1136];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????:
        _5315_ = b[1167:1152];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????:
        _5315_ = b[1183:1168];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????:
        _5315_ = b[1199:1184];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????:
        _5315_ = b[1215:1200];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????:
        _5315_ = b[1231:1216];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????:
        _5315_ = b[1247:1232];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????:
        _5315_ = b[1263:1248];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????:
        _5315_ = b[1279:1264];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????:
        _5315_ = b[1295:1280];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????:
        _5315_ = b[1311:1296];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????:
        _5315_ = b[1327:1312];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????:
        _5315_ = b[1343:1328];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????:
        _5315_ = b[1359:1344];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????:
        _5315_ = b[1375:1360];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????:
        _5315_ = b[1391:1376];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????:
        _5315_ = b[1407:1392];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????:
        _5315_ = b[1423:1408];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????:
        _5315_ = b[1439:1424];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????:
        _5315_ = b[1455:1440];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????:
        _5315_ = b[1471:1456];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????:
        _5315_ = b[1487:1472];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????:
        _5315_ = b[1503:1488];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????:
        _5315_ = b[1519:1504];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????:
        _5315_ = b[1535:1520];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????:
        _5315_ = b[1551:1536];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????:
        _5315_ = b[1567:1552];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????:
        _5315_ = b[1583:1568];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????:
        _5315_ = b[1599:1584];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5315_ = b[1615:1600];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5315_ = b[1631:1616];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5315_ = b[1647:1632];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5315_ = b[1663:1648];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5315_ = b[1679:1664];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5315_ = b[1695:1680];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5315_ = b[1711:1696];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5315_ = b[1727:1712];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5315_ = b[1743:1728];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5315_ = b[1759:1744];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5315_ = b[1775:1760];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5315_ = b[1791:1776];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5315_ = b[1807:1792];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5315_ = b[1823:1808];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5315_ = b[1839:1824];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5315_ = b[1855:1840];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5315_ = b[1871:1856];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5315_ = b[1887:1872];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5315_ = b[1903:1888];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5315_ = b[1919:1904];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5315_ = b[1935:1920];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5315_ = b[1951:1936];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5315_ = b[1967:1952];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5315_ = b[1983:1968];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5315_ = b[1999:1984];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5315_ = b[2015:2000];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5315_ = b[2031:2016];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5315_ = b[2047:2032];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5315_ = b[2063:2048];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5315_ = b[2079:2064];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5315_ = b[2095:2080];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5315_ = b[2111:2096];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5315_ = b[2127:2112];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5315_ = b[2143:2128];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5315_ = b[2159:2144];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5315_ = b[2175:2160];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5315_ = b[2191:2176];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5315_ = b[2207:2192];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5315_ = b[2223:2208];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5315_ = b[2239:2224];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5315_ = b[2255:2240];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5315_ = b[2271:2256];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5315_ = b[2287:2272];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5315_ = b[2303:2288];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5315_ = b[2319:2304];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5315_ = b[2335:2320];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5315_ = b[2351:2336];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5315_ = b[2367:2352];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5315_ = b[2383:2368];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5315_ = b[2399:2384];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5315_ = b[2415:2400];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5315_ = b[2431:2416];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5315_ = b[2447:2432];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5315_ = b[2463:2448];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5315_ = b[2479:2464];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5315_ = b[2495:2480];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5315_ = b[2511:2496];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5315_ = b[2527:2512];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5315_ = b[2543:2528];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5315_ = b[2559:2544];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5315_ = b[2575:2560];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5315_ = b[2591:2576];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5315_ = b[2607:2592];
      256'b????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5315_ = b[2623:2608];
      256'b???????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5315_ = b[2639:2624];
      256'b??????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5315_ = b[2655:2640];
      256'b?????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5315_ = b[2671:2656];
      256'b????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5315_ = b[2687:2672];
      256'b???????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5315_ = b[2703:2688];
      256'b??????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5315_ = b[2719:2704];
      256'b?????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5315_ = b[2735:2720];
      256'b????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5315_ = b[2751:2736];
      256'b???????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5315_ = b[2767:2752];
      256'b??????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5315_ = b[2783:2768];
      256'b?????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5315_ = b[2799:2784];
      256'b????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5315_ = b[2815:2800];
      256'b???????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5315_ = b[2831:2816];
      256'b??????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5315_ = b[2847:2832];
      256'b?????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5315_ = b[2863:2848];
      256'b????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5315_ = b[2879:2864];
      256'b???????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5315_ = b[2895:2880];
      256'b??????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5315_ = b[2911:2896];
      256'b?????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5315_ = b[2927:2912];
      256'b????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5315_ = b[2943:2928];
      256'b???????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5315_ = b[2959:2944];
      256'b??????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5315_ = b[2975:2960];
      256'b?????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5315_ = b[2991:2976];
      256'b????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5315_ = b[3007:2992];
      256'b???????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5315_ = b[3023:3008];
      256'b??????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5315_ = b[3039:3024];
      256'b?????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5315_ = b[3055:3040];
      256'b????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5315_ = b[3071:3056];
      256'b???????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5315_ = b[3087:3072];
      256'b??????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5315_ = b[3103:3088];
      256'b?????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5315_ = b[3119:3104];
      256'b????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5315_ = b[3135:3120];
      256'b???????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5315_ = b[3151:3136];
      256'b??????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5315_ = b[3167:3152];
      256'b?????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5315_ = b[3183:3168];
      256'b????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5315_ = b[3199:3184];
      256'b???????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5315_ = b[3215:3200];
      256'b??????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5315_ = b[3231:3216];
      256'b?????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5315_ = b[3247:3232];
      256'b????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5315_ = b[3263:3248];
      256'b???????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5315_ = b[3279:3264];
      256'b??????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5315_ = b[3295:3280];
      256'b?????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5315_ = b[3311:3296];
      256'b????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5315_ = b[3327:3312];
      256'b???????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5315_ = b[3343:3328];
      256'b??????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5315_ = b[3359:3344];
      256'b?????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5315_ = b[3375:3360];
      256'b????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5315_ = b[3391:3376];
      256'b???????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5315_ = b[3407:3392];
      256'b??????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5315_ = b[3423:3408];
      256'b?????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5315_ = b[3439:3424];
      256'b????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5315_ = b[3455:3440];
      256'b???????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5315_ = b[3471:3456];
      256'b??????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5315_ = b[3487:3472];
      256'b?????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5315_ = b[3503:3488];
      256'b????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5315_ = b[3519:3504];
      256'b???????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5315_ = b[3535:3520];
      256'b??????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5315_ = b[3551:3536];
      256'b?????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5315_ = b[3567:3552];
      256'b????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5315_ = b[3583:3568];
      256'b???????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5315_ = b[3599:3584];
      256'b??????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5315_ = b[3615:3600];
      256'b?????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5315_ = b[3631:3616];
      256'b????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5315_ = b[3647:3632];
      256'b???????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5315_ = b[3663:3648];
      256'b??????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5315_ = b[3679:3664];
      256'b?????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5315_ = b[3695:3680];
      256'b????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5315_ = b[3711:3696];
      256'b???????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5315_ = b[3727:3712];
      256'b??????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5315_ = b[3743:3728];
      256'b?????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5315_ = b[3759:3744];
      256'b????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5315_ = b[3775:3760];
      256'b???????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5315_ = b[3791:3776];
      256'b??????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5315_ = b[3807:3792];
      256'b?????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5315_ = b[3823:3808];
      256'b????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5315_ = b[3839:3824];
      256'b???????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5315_ = b[3855:3840];
      256'b??????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5315_ = b[3871:3856];
      256'b?????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5315_ = b[3887:3872];
      256'b????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5315_ = b[3903:3888];
      256'b???????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5315_ = b[3919:3904];
      256'b??????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5315_ = b[3935:3920];
      256'b?????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5315_ = b[3951:3936];
      256'b????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5315_ = b[3967:3952];
      256'b???????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5315_ = b[3983:3968];
      256'b??????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5315_ = b[3999:3984];
      256'b?????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5315_ = b[4015:4000];
      256'b????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5315_ = b[4031:4016];
      256'b???1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5315_ = b[4047:4032];
      256'b??1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5315_ = b[4063:4048];
      256'b?1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5315_ = b[4079:4064];
      256'b1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5315_ = b[4095:4080];
      default:
        _5315_ = a;
    endcase
  endfunction
  assign _1467_ = _5315_(density_reg0, { density_reg1, density_reg2, density_reg3, density_reg4, density_reg5, density_reg6, density_reg7, density_reg8, density_reg9, density_reg10, density_reg11, density_reg12, density_reg13, density_reg14, density_reg15, density_reg16, density_reg17, density_reg18, density_reg19, density_reg20, density_reg21, density_reg22, density_reg23, density_reg24, density_reg25, density_reg26, density_reg27, density_reg28, density_reg29, density_reg30, density_reg31, density_reg32, density_reg33, density_reg34, density_reg35, density_reg36, density_reg37, density_reg38, density_reg39, density_reg40, density_reg41, density_reg42, density_reg43, density_reg44, density_reg45, density_reg46, density_reg47, density_reg48, density_reg49, density_reg50, density_reg51, density_reg52, density_reg53, density_reg54, density_reg55, density_reg56, density_reg57, density_reg58, density_reg59, density_reg60, density_reg61, density_reg62, density_reg63, density_reg64, density_reg65, density_reg66, density_reg67, density_reg68, density_reg69, density_reg70, density_reg71, density_reg72, density_reg73, density_reg74, density_reg75, density_reg76, density_reg77, density_reg78, density_reg79, density_reg80, density_reg81, density_reg82, density_reg83, density_reg84, density_reg85, density_reg86, density_reg87, density_reg88, density_reg89, density_reg90, density_reg91, density_reg92, density_reg93, density_reg94, density_reg95, density_reg96, density_reg97, density_reg98, density_reg99, density_reg100, density_reg101, density_reg102, density_reg103, density_reg104, density_reg105, density_reg106, density_reg107, density_reg108, density_reg109, density_reg110, density_reg111, density_reg112, density_reg113, density_reg114, density_reg115, density_reg116, density_reg117, density_reg118, density_reg119, density_reg120, density_reg121, density_reg122, density_reg123, density_reg124, density_reg125, density_reg126, density_reg127, density_reg128, density_reg129, density_reg130, density_reg131, density_reg132, density_reg133, density_reg134, density_reg135, density_reg136, density_reg137, density_reg138, density_reg139, density_reg140, density_reg141, density_reg142, density_reg143, density_reg144, density_reg145, density_reg146, density_reg147, density_reg148, density_reg149, density_reg150, density_reg151, density_reg152, density_reg153, density_reg154, density_reg155, density_reg156, density_reg157, density_reg158, density_reg159, density_reg160, density_reg161, density_reg162, density_reg163, density_reg164, density_reg165, density_reg166, density_reg167, density_reg168, density_reg169, density_reg170, density_reg171, density_reg172, density_reg173, density_reg174, density_reg175, density_reg176, density_reg177, density_reg178, density_reg179, density_reg180, density_reg181, density_reg182, density_reg183, density_reg184, density_reg185, density_reg186, density_reg187, density_reg188, density_reg189, density_reg190, density_reg191, density_reg192, density_reg193, density_reg194, density_reg195, density_reg196, density_reg197, density_reg198, density_reg199, density_reg200, density_reg201, density_reg202, density_reg203, density_reg204, density_reg205, density_reg206, density_reg207, density_reg208, density_reg209, density_reg210, density_reg211, density_reg212, density_reg213, density_reg214, density_reg215, density_reg216, density_reg217, density_reg218, density_reg219, density_reg220, density_reg221, density_reg222, density_reg223, density_reg224, density_reg225, density_reg226, density_reg227, density_reg228, density_reg229, density_reg230, density_reg231, density_reg232, density_reg233, density_reg234, density_reg235, density_reg236, density_reg237, density_reg238, density_reg239, density_reg240, density_reg241, density_reg242, density_reg243, density_reg244, density_reg245, density_reg246, density_reg247, density_reg248, density_reg249, density_reg250, density_reg251, density_reg252, density_reg253, density_reg254, density_reg255, density_reg256 }, { _1463_, _1462_, _1461_, _1460_, _1459_, _1458_, _1457_, _1456_, _1455_, _1454_, _1453_, _1452_, _1451_, _1450_, _1449_, _1448_, _1447_, _1446_, _1445_, _1444_, _1443_, _1442_, _1441_, _1440_, _1439_, _1438_, _1437_, _1436_, _1435_, _1434_, _1433_, _1432_, _1431_, _1430_, _1429_, _1428_, _1427_, _1426_, _1425_, _1424_, _1423_, _1422_, _1421_, _1420_, _1419_, _1418_, _1417_, _1416_, _1415_, _1414_, _1413_, _1412_, _1411_, _1410_, _1409_, _1408_, _1407_, _1406_, _1405_, _1404_, _1403_, _1402_, _1401_, _1400_, _1399_, _1398_, _1397_, _1396_, _1395_, _1394_, _1393_, _1392_, _1391_, _1390_, _1389_, _1388_, _1387_, _1386_, _1385_, _1384_, _1383_, _1382_, _1381_, _1380_, _1379_, _1378_, _1377_, _1376_, _1375_, _1374_, _1373_, _1372_, _1371_, _1370_, _1369_, _1368_, _1367_, _1366_, _1365_, _1364_, _1363_, _1362_, _1361_, _1360_, _1359_, _1358_, _1357_, _1356_, _1355_, _1354_, _1353_, _1352_, _1351_, _1350_, _1349_, _1348_, _1347_, _1346_, _1345_, _1344_, _1343_, _1342_, _1341_, _1340_, _1339_, _1338_, _1337_, _1336_, _1335_, _1334_, _1333_, _1332_, _1331_, _1330_, _1329_, _1328_, _1327_, _1326_, _1325_, _1324_, _1323_, _1322_, _1321_, _1320_, _1319_, _1318_, _1317_, _1316_, _1315_, _1314_, _1313_, _1312_, _1311_, _1310_, _1309_, _1308_, _1307_, _1306_, _1305_, _1304_, _1303_, _1302_, _1301_, _1300_, _1299_, _1298_, _1297_, _1296_, _1295_, _1294_, _1293_, _1292_, _1291_, _1290_, _1289_, _1288_, _1287_, _1286_, _1285_, _1284_, _1283_, _1282_, _1281_, _1280_, _1279_, _1278_, _1277_, _1276_, _1275_, _1274_, _1273_, _1272_, _1271_, _1270_, _1269_, _1268_, _1267_, _1266_, _1265_, _1264_, _1263_, _1262_, _1261_, _1260_, _1259_, _1258_, _1257_, _1256_, _1255_, _1254_, _1253_, _1252_, _1251_, _1250_, _1249_, _1248_, _1247_, _1246_, _1245_, _1244_, _1243_, _1242_, _1241_, _1240_, _1239_, _1238_, _1237_, _1236_, _1235_, _1234_, _1233_, _1232_, _1231_, _1230_, _1229_, _1228_, _1227_, _1226_, _1225_, _1224_, _1223_, _1222_, _1221_, _1220_, _1219_, _1218_, _1217_, _1216_, _1215_, _1214_, _1213_, _1212_, _1211_, _1210_, _1209_, _1208_ });
  assign _1468_ = dp2lut_Yinfo_5[17] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12474" *) density_reg256 : _1467_;
  assign _1469_ = dp2lut_Yinfo_5[16] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12471" *) density_reg0 : _1468_;
  assign _0295_ = _0388_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12470" *) _1469_ : lut_Y_data_50;
  function [15:0] _5319_;
    input [15:0] a;
    input [4095:0] b;
    input [255:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12452|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *)
    (* parallel_case *)
    casez (s)
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1:
        _5319_ = b[15:0];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?:
        _5319_ = b[31:16];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??:
        _5319_ = b[47:32];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???:
        _5319_ = b[63:48];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????:
        _5319_ = b[79:64];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????:
        _5319_ = b[95:80];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????:
        _5319_ = b[111:96];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????:
        _5319_ = b[127:112];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????:
        _5319_ = b[143:128];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????:
        _5319_ = b[159:144];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????:
        _5319_ = b[175:160];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????:
        _5319_ = b[191:176];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????:
        _5319_ = b[207:192];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????:
        _5319_ = b[223:208];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????:
        _5319_ = b[239:224];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????:
        _5319_ = b[255:240];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????:
        _5319_ = b[271:256];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????:
        _5319_ = b[287:272];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????:
        _5319_ = b[303:288];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????:
        _5319_ = b[319:304];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????:
        _5319_ = b[335:320];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????:
        _5319_ = b[351:336];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????:
        _5319_ = b[367:352];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????:
        _5319_ = b[383:368];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????:
        _5319_ = b[399:384];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????:
        _5319_ = b[415:400];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????:
        _5319_ = b[431:416];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????:
        _5319_ = b[447:432];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????:
        _5319_ = b[463:448];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????:
        _5319_ = b[479:464];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????:
        _5319_ = b[495:480];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????:
        _5319_ = b[511:496];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????:
        _5319_ = b[527:512];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????:
        _5319_ = b[543:528];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????:
        _5319_ = b[559:544];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????:
        _5319_ = b[575:560];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????:
        _5319_ = b[591:576];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????:
        _5319_ = b[607:592];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????:
        _5319_ = b[623:608];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????:
        _5319_ = b[639:624];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????:
        _5319_ = b[655:640];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????:
        _5319_ = b[671:656];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????:
        _5319_ = b[687:672];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????:
        _5319_ = b[703:688];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????:
        _5319_ = b[719:704];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????:
        _5319_ = b[735:720];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????:
        _5319_ = b[751:736];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????:
        _5319_ = b[767:752];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????:
        _5319_ = b[783:768];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????:
        _5319_ = b[799:784];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????:
        _5319_ = b[815:800];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????:
        _5319_ = b[831:816];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????:
        _5319_ = b[847:832];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????:
        _5319_ = b[863:848];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????:
        _5319_ = b[879:864];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????:
        _5319_ = b[895:880];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????:
        _5319_ = b[911:896];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????:
        _5319_ = b[927:912];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????:
        _5319_ = b[943:928];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????:
        _5319_ = b[959:944];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????:
        _5319_ = b[975:960];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????:
        _5319_ = b[991:976];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????:
        _5319_ = b[1007:992];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????:
        _5319_ = b[1023:1008];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????:
        _5319_ = b[1039:1024];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????:
        _5319_ = b[1055:1040];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????:
        _5319_ = b[1071:1056];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????:
        _5319_ = b[1087:1072];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????:
        _5319_ = b[1103:1088];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????:
        _5319_ = b[1119:1104];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????:
        _5319_ = b[1135:1120];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????:
        _5319_ = b[1151:1136];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????:
        _5319_ = b[1167:1152];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????:
        _5319_ = b[1183:1168];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????:
        _5319_ = b[1199:1184];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????:
        _5319_ = b[1215:1200];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????:
        _5319_ = b[1231:1216];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????:
        _5319_ = b[1247:1232];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????:
        _5319_ = b[1263:1248];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????:
        _5319_ = b[1279:1264];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????:
        _5319_ = b[1295:1280];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????:
        _5319_ = b[1311:1296];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????:
        _5319_ = b[1327:1312];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????:
        _5319_ = b[1343:1328];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????:
        _5319_ = b[1359:1344];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????:
        _5319_ = b[1375:1360];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????:
        _5319_ = b[1391:1376];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????:
        _5319_ = b[1407:1392];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????:
        _5319_ = b[1423:1408];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????:
        _5319_ = b[1439:1424];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????:
        _5319_ = b[1455:1440];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????:
        _5319_ = b[1471:1456];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????:
        _5319_ = b[1487:1472];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????:
        _5319_ = b[1503:1488];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????:
        _5319_ = b[1519:1504];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????:
        _5319_ = b[1535:1520];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????:
        _5319_ = b[1551:1536];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????:
        _5319_ = b[1567:1552];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????:
        _5319_ = b[1583:1568];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????:
        _5319_ = b[1599:1584];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5319_ = b[1615:1600];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5319_ = b[1631:1616];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5319_ = b[1647:1632];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5319_ = b[1663:1648];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5319_ = b[1679:1664];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5319_ = b[1695:1680];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5319_ = b[1711:1696];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5319_ = b[1727:1712];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5319_ = b[1743:1728];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5319_ = b[1759:1744];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5319_ = b[1775:1760];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5319_ = b[1791:1776];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5319_ = b[1807:1792];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5319_ = b[1823:1808];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5319_ = b[1839:1824];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5319_ = b[1855:1840];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5319_ = b[1871:1856];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5319_ = b[1887:1872];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5319_ = b[1903:1888];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5319_ = b[1919:1904];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5319_ = b[1935:1920];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5319_ = b[1951:1936];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5319_ = b[1967:1952];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5319_ = b[1983:1968];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5319_ = b[1999:1984];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5319_ = b[2015:2000];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5319_ = b[2031:2016];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5319_ = b[2047:2032];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5319_ = b[2063:2048];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5319_ = b[2079:2064];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5319_ = b[2095:2080];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5319_ = b[2111:2096];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5319_ = b[2127:2112];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5319_ = b[2143:2128];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5319_ = b[2159:2144];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5319_ = b[2175:2160];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5319_ = b[2191:2176];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5319_ = b[2207:2192];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5319_ = b[2223:2208];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5319_ = b[2239:2224];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5319_ = b[2255:2240];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5319_ = b[2271:2256];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5319_ = b[2287:2272];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5319_ = b[2303:2288];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5319_ = b[2319:2304];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5319_ = b[2335:2320];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5319_ = b[2351:2336];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5319_ = b[2367:2352];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5319_ = b[2383:2368];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5319_ = b[2399:2384];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5319_ = b[2415:2400];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5319_ = b[2431:2416];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5319_ = b[2447:2432];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5319_ = b[2463:2448];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5319_ = b[2479:2464];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5319_ = b[2495:2480];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5319_ = b[2511:2496];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5319_ = b[2527:2512];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5319_ = b[2543:2528];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5319_ = b[2559:2544];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5319_ = b[2575:2560];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5319_ = b[2591:2576];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5319_ = b[2607:2592];
      256'b????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5319_ = b[2623:2608];
      256'b???????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5319_ = b[2639:2624];
      256'b??????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5319_ = b[2655:2640];
      256'b?????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5319_ = b[2671:2656];
      256'b????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5319_ = b[2687:2672];
      256'b???????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5319_ = b[2703:2688];
      256'b??????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5319_ = b[2719:2704];
      256'b?????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5319_ = b[2735:2720];
      256'b????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5319_ = b[2751:2736];
      256'b???????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5319_ = b[2767:2752];
      256'b??????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5319_ = b[2783:2768];
      256'b?????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5319_ = b[2799:2784];
      256'b????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5319_ = b[2815:2800];
      256'b???????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5319_ = b[2831:2816];
      256'b??????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5319_ = b[2847:2832];
      256'b?????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5319_ = b[2863:2848];
      256'b????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5319_ = b[2879:2864];
      256'b???????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5319_ = b[2895:2880];
      256'b??????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5319_ = b[2911:2896];
      256'b?????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5319_ = b[2927:2912];
      256'b????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5319_ = b[2943:2928];
      256'b???????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5319_ = b[2959:2944];
      256'b??????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5319_ = b[2975:2960];
      256'b?????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5319_ = b[2991:2976];
      256'b????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5319_ = b[3007:2992];
      256'b???????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5319_ = b[3023:3008];
      256'b??????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5319_ = b[3039:3024];
      256'b?????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5319_ = b[3055:3040];
      256'b????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5319_ = b[3071:3056];
      256'b???????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5319_ = b[3087:3072];
      256'b??????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5319_ = b[3103:3088];
      256'b?????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5319_ = b[3119:3104];
      256'b????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5319_ = b[3135:3120];
      256'b???????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5319_ = b[3151:3136];
      256'b??????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5319_ = b[3167:3152];
      256'b?????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5319_ = b[3183:3168];
      256'b????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5319_ = b[3199:3184];
      256'b???????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5319_ = b[3215:3200];
      256'b??????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5319_ = b[3231:3216];
      256'b?????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5319_ = b[3247:3232];
      256'b????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5319_ = b[3263:3248];
      256'b???????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5319_ = b[3279:3264];
      256'b??????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5319_ = b[3295:3280];
      256'b?????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5319_ = b[3311:3296];
      256'b????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5319_ = b[3327:3312];
      256'b???????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5319_ = b[3343:3328];
      256'b??????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5319_ = b[3359:3344];
      256'b?????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5319_ = b[3375:3360];
      256'b????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5319_ = b[3391:3376];
      256'b???????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5319_ = b[3407:3392];
      256'b??????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5319_ = b[3423:3408];
      256'b?????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5319_ = b[3439:3424];
      256'b????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5319_ = b[3455:3440];
      256'b???????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5319_ = b[3471:3456];
      256'b??????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5319_ = b[3487:3472];
      256'b?????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5319_ = b[3503:3488];
      256'b????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5319_ = b[3519:3504];
      256'b???????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5319_ = b[3535:3520];
      256'b??????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5319_ = b[3551:3536];
      256'b?????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5319_ = b[3567:3552];
      256'b????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5319_ = b[3583:3568];
      256'b???????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5319_ = b[3599:3584];
      256'b??????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5319_ = b[3615:3600];
      256'b?????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5319_ = b[3631:3616];
      256'b????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5319_ = b[3647:3632];
      256'b???????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5319_ = b[3663:3648];
      256'b??????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5319_ = b[3679:3664];
      256'b?????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5319_ = b[3695:3680];
      256'b????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5319_ = b[3711:3696];
      256'b???????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5319_ = b[3727:3712];
      256'b??????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5319_ = b[3743:3728];
      256'b?????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5319_ = b[3759:3744];
      256'b????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5319_ = b[3775:3760];
      256'b???????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5319_ = b[3791:3776];
      256'b??????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5319_ = b[3807:3792];
      256'b?????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5319_ = b[3823:3808];
      256'b????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5319_ = b[3839:3824];
      256'b???????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5319_ = b[3855:3840];
      256'b??????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5319_ = b[3871:3856];
      256'b?????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5319_ = b[3887:3872];
      256'b????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5319_ = b[3903:3888];
      256'b???????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5319_ = b[3919:3904];
      256'b??????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5319_ = b[3935:3920];
      256'b?????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5319_ = b[3951:3936];
      256'b????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5319_ = b[3967:3952];
      256'b???????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5319_ = b[3983:3968];
      256'b??????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5319_ = b[3999:3984];
      256'b?????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5319_ = b[4015:4000];
      256'b????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5319_ = b[4031:4016];
      256'b???1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5319_ = b[4047:4032];
      256'b??1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5319_ = b[4063:4048];
      256'b?1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5319_ = b[4079:4064];
      256'b1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5319_ = b[4095:4080];
      default:
        _5319_ = a;
    endcase
  endfunction
  assign _1470_ = _5319_(density_reg0, { density_reg1, density_reg2, density_reg3, density_reg4, density_reg5, density_reg6, density_reg7, density_reg8, density_reg9, density_reg10, density_reg11, density_reg12, density_reg13, density_reg14, density_reg15, density_reg16, density_reg17, density_reg18, density_reg19, density_reg20, density_reg21, density_reg22, density_reg23, density_reg24, density_reg25, density_reg26, density_reg27, density_reg28, density_reg29, density_reg30, density_reg31, density_reg32, density_reg33, density_reg34, density_reg35, density_reg36, density_reg37, density_reg38, density_reg39, density_reg40, density_reg41, density_reg42, density_reg43, density_reg44, density_reg45, density_reg46, density_reg47, density_reg48, density_reg49, density_reg50, density_reg51, density_reg52, density_reg53, density_reg54, density_reg55, density_reg56, density_reg57, density_reg58, density_reg59, density_reg60, density_reg61, density_reg62, density_reg63, density_reg64, density_reg65, density_reg66, density_reg67, density_reg68, density_reg69, density_reg70, density_reg71, density_reg72, density_reg73, density_reg74, density_reg75, density_reg76, density_reg77, density_reg78, density_reg79, density_reg80, density_reg81, density_reg82, density_reg83, density_reg84, density_reg85, density_reg86, density_reg87, density_reg88, density_reg89, density_reg90, density_reg91, density_reg92, density_reg93, density_reg94, density_reg95, density_reg96, density_reg97, density_reg98, density_reg99, density_reg100, density_reg101, density_reg102, density_reg103, density_reg104, density_reg105, density_reg106, density_reg107, density_reg108, density_reg109, density_reg110, density_reg111, density_reg112, density_reg113, density_reg114, density_reg115, density_reg116, density_reg117, density_reg118, density_reg119, density_reg120, density_reg121, density_reg122, density_reg123, density_reg124, density_reg125, density_reg126, density_reg127, density_reg128, density_reg129, density_reg130, density_reg131, density_reg132, density_reg133, density_reg134, density_reg135, density_reg136, density_reg137, density_reg138, density_reg139, density_reg140, density_reg141, density_reg142, density_reg143, density_reg144, density_reg145, density_reg146, density_reg147, density_reg148, density_reg149, density_reg150, density_reg151, density_reg152, density_reg153, density_reg154, density_reg155, density_reg156, density_reg157, density_reg158, density_reg159, density_reg160, density_reg161, density_reg162, density_reg163, density_reg164, density_reg165, density_reg166, density_reg167, density_reg168, density_reg169, density_reg170, density_reg171, density_reg172, density_reg173, density_reg174, density_reg175, density_reg176, density_reg177, density_reg178, density_reg179, density_reg180, density_reg181, density_reg182, density_reg183, density_reg184, density_reg185, density_reg186, density_reg187, density_reg188, density_reg189, density_reg190, density_reg191, density_reg192, density_reg193, density_reg194, density_reg195, density_reg196, density_reg197, density_reg198, density_reg199, density_reg200, density_reg201, density_reg202, density_reg203, density_reg204, density_reg205, density_reg206, density_reg207, density_reg208, density_reg209, density_reg210, density_reg211, density_reg212, density_reg213, density_reg214, density_reg215, density_reg216, density_reg217, density_reg218, density_reg219, density_reg220, density_reg221, density_reg222, density_reg223, density_reg224, density_reg225, density_reg226, density_reg227, density_reg228, density_reg229, density_reg230, density_reg231, density_reg232, density_reg233, density_reg234, density_reg235, density_reg236, density_reg237, density_reg238, density_reg239, density_reg240, density_reg241, density_reg242, density_reg243, density_reg244, density_reg245, density_reg246, density_reg247, density_reg248, density_reg249, density_reg250, density_reg251, density_reg252, density_reg253, density_reg254, density_reg255, density_reg256 }, { _1727_, _1726_, _1725_, _1724_, _1723_, _1722_, _1721_, _1720_, _1719_, _1718_, _1717_, _1716_, _1715_, _1714_, _1713_, _1712_, _1711_, _1710_, _1709_, _1708_, _1707_, _1706_, _1705_, _1704_, _1703_, _1702_, _1701_, _1700_, _1699_, _1698_, _1697_, _1696_, _1695_, _1694_, _1693_, _1692_, _1691_, _1690_, _1689_, _1688_, _1687_, _1686_, _1685_, _1684_, _1683_, _1682_, _1681_, _1680_, _1679_, _1678_, _1677_, _1676_, _1675_, _1674_, _1673_, _1672_, _1671_, _1670_, _1669_, _1668_, _1667_, _1666_, _1665_, _1664_, _1663_, _1662_, _1661_, _1660_, _1659_, _1658_, _1657_, _1656_, _1655_, _1654_, _1653_, _1652_, _1651_, _1650_, _1649_, _1648_, _1647_, _1646_, _1645_, _1644_, _1643_, _1642_, _1641_, _1640_, _1639_, _1638_, _1637_, _1636_, _1635_, _1634_, _1633_, _1632_, _1631_, _1630_, _1629_, _1628_, _1627_, _1626_, _1625_, _1624_, _1623_, _1622_, _1621_, _1620_, _1619_, _1618_, _1617_, _1616_, _1615_, _1614_, _1613_, _1612_, _1611_, _1610_, _1609_, _1608_, _1607_, _1606_, _1605_, _1604_, _1603_, _1602_, _1601_, _1600_, _1599_, _1598_, _1597_, _1596_, _1595_, _1594_, _1593_, _1592_, _1591_, _1590_, _1589_, _1588_, _1587_, _1586_, _1585_, _1584_, _1583_, _1582_, _1581_, _1580_, _1579_, _1578_, _1577_, _1576_, _1575_, _1574_, _1573_, _1572_, _1571_, _1570_, _1569_, _1568_, _1567_, _1566_, _1565_, _1564_, _1563_, _1562_, _1561_, _1560_, _1559_, _1558_, _1557_, _1556_, _1555_, _1554_, _1553_, _1552_, _1551_, _1550_, _1549_, _1548_, _1547_, _1546_, _1545_, _1544_, _1543_, _1542_, _1541_, _1540_, _1539_, _1538_, _1537_, _1536_, _1535_, _1534_, _1533_, _1532_, _1531_, _1530_, _1529_, _1528_, _1527_, _1526_, _1525_, _1524_, _1523_, _1522_, _1521_, _1520_, _1519_, _1518_, _1517_, _1516_, _1515_, _1514_, _1513_, _1512_, _1511_, _1510_, _1509_, _1508_, _1507_, _1506_, _1505_, _1504_, _1503_, _1502_, _1501_, _1500_, _1499_, _1498_, _1497_, _1496_, _1495_, _1494_, _1493_, _1492_, _1491_, _1490_, _1489_, _1488_, _1487_, _1486_, _1485_, _1484_, _1483_, _1482_, _1481_, _1480_, _1479_, _1478_, _1477_, _1476_, _1475_, _1474_, _1473_, _0414_ });
  assign _1471_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12452|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 9'b100000000;
  assign _1472_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12448|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 8'b11111111;
  assign _1473_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12444|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 8'b11111110;
  assign _1474_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12440|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 8'b11111101;
  assign _1475_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12436|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 8'b11111100;
  assign _1476_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12432|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 8'b11111011;
  assign _1477_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12428|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 8'b11111010;
  assign _1478_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12424|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 8'b11111001;
  assign _1479_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12420|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 8'b11111000;
  assign _1480_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12416|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 8'b11110111;
  assign _1481_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12412|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 8'b11110110;
  assign _1482_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12408|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 8'b11110101;
  assign _1483_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12404|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 8'b11110100;
  assign _1484_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12400|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 8'b11110011;
  assign _1485_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12396|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 8'b11110010;
  assign _1486_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12392|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 8'b11110001;
  assign _1487_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12388|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 8'b11110000;
  assign _1488_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12384|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 8'b11101111;
  assign _1489_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12380|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 8'b11101110;
  assign _1490_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12376|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 8'b11101101;
  assign _1491_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12372|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 8'b11101100;
  assign _1492_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12368|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 8'b11101011;
  assign _1493_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12364|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 8'b11101010;
  assign _1494_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12360|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 8'b11101001;
  assign _1495_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12356|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 8'b11101000;
  assign _1496_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12352|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 8'b11100111;
  assign _1497_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12348|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 8'b11100110;
  assign _1498_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12344|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 8'b11100101;
  assign _1499_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12340|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 8'b11100100;
  assign _1500_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12336|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 8'b11100011;
  assign _1501_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12332|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 8'b11100010;
  assign _1502_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12328|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 8'b11100001;
  assign _1503_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12324|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 8'b11100000;
  assign _1504_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12320|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 8'b11011111;
  assign _1505_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12316|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 8'b11011110;
  assign _1506_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12312|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 8'b11011101;
  assign _1507_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12308|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 8'b11011100;
  assign _1508_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12304|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 8'b11011011;
  assign _1509_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12300|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 8'b11011010;
  assign _1510_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12296|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 8'b11011001;
  assign _1511_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12292|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 8'b11011000;
  assign _1512_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12288|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 8'b11010111;
  assign _1513_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12284|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 8'b11010110;
  assign _1514_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12280|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 8'b11010101;
  assign _1515_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12276|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 8'b11010100;
  assign _1516_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12272|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 8'b11010011;
  assign _1517_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12268|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 8'b11010010;
  assign _1518_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12264|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 8'b11010001;
  assign _1519_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12260|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 8'b11010000;
  assign _1520_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12256|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 8'b11001111;
  assign _1521_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12252|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 8'b11001110;
  assign _1522_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12248|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 8'b11001101;
  assign _1523_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12244|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 8'b11001100;
  assign _1524_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12240|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 8'b11001011;
  assign _1525_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12236|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 8'b11001010;
  assign _1526_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12232|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 8'b11001001;
  assign _1527_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12228|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 8'b11001000;
  assign _1528_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12224|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 8'b11000111;
  assign _1529_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12220|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 8'b11000110;
  assign _1530_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12216|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 8'b11000101;
  assign _1531_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12212|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 8'b11000100;
  assign _1532_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12208|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 8'b11000011;
  assign _1533_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12204|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 8'b11000010;
  assign _1534_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12200|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 8'b11000001;
  assign _1535_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12196|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 8'b11000000;
  assign _1536_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12192|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 8'b10111111;
  assign _1537_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12188|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 8'b10111110;
  assign _1538_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12184|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 8'b10111101;
  assign _1539_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12180|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 8'b10111100;
  assign _1540_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12176|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 8'b10111011;
  assign _1541_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12172|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 8'b10111010;
  assign _1542_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12168|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 8'b10111001;
  assign _1543_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12164|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 8'b10111000;
  assign _1544_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12160|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 8'b10110111;
  assign _1545_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12156|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 8'b10110110;
  assign _1546_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12152|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 8'b10110101;
  assign _1547_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12148|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 8'b10110100;
  assign _1548_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12144|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 8'b10110011;
  assign _1549_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12140|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 8'b10110010;
  assign _1550_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12136|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 8'b10110001;
  assign _1551_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12132|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 8'b10110000;
  assign _1552_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12128|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 8'b10101111;
  assign _1553_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12124|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 8'b10101110;
  assign _1554_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12120|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 8'b10101101;
  assign _1555_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12116|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 8'b10101100;
  assign _1556_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12112|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 8'b10101011;
  assign _1557_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12108|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 8'b10101010;
  assign _1558_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12104|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 8'b10101001;
  assign _1559_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12100|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 8'b10101000;
  assign _1560_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12096|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 8'b10100111;
  assign _1561_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12092|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 8'b10100110;
  assign _1562_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12088|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 8'b10100101;
  assign _1563_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12084|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 8'b10100100;
  assign _1564_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12080|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 8'b10100011;
  assign _1565_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12076|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 8'b10100010;
  assign _1566_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12072|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 8'b10100001;
  assign _1567_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12068|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 8'b10100000;
  assign _1568_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12064|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 8'b10011111;
  assign _1569_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12060|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 8'b10011110;
  assign _1570_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12056|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 8'b10011101;
  assign _1571_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12052|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 8'b10011100;
  assign _1572_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12048|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 8'b10011011;
  assign _1573_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12044|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 8'b10011010;
  assign _1574_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12040|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 8'b10011001;
  assign _1575_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12036|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 8'b10011000;
  assign _1576_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12032|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 8'b10010111;
  assign _1577_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12028|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 8'b10010110;
  assign _1578_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12024|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 8'b10010101;
  assign _1579_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12020|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 8'b10010100;
  assign _1580_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12016|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 8'b10010011;
  assign _1581_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12012|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 8'b10010010;
  assign _1582_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12008|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 8'b10010001;
  assign _1583_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12004|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 8'b10010000;
  assign _1584_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12000|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 8'b10001111;
  assign _1585_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11996|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 8'b10001110;
  assign _1586_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11992|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 8'b10001101;
  assign _1587_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11988|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 8'b10001100;
  assign _1588_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11984|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 8'b10001011;
  assign _1589_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11980|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 8'b10001010;
  assign _1590_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11976|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 8'b10001001;
  assign _1591_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11972|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 8'b10001000;
  assign _1592_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11968|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 8'b10000111;
  assign _1593_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11964|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 8'b10000110;
  assign _1594_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11960|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 8'b10000101;
  assign _1595_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11956|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 8'b10000100;
  assign _1596_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11952|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 8'b10000011;
  assign _1597_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11948|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 8'b10000010;
  assign _1598_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11944|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 8'b10000001;
  assign _1599_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11940|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 8'b10000000;
  assign _1600_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11936|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 7'b1111111;
  assign _1601_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11932|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 7'b1111110;
  assign _1602_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11928|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 7'b1111101;
  assign _1603_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11924|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 7'b1111100;
  assign _1604_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11920|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 7'b1111011;
  assign _1605_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11916|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 7'b1111010;
  assign _1606_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11912|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 7'b1111001;
  assign _1607_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11908|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 7'b1111000;
  assign _1608_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11904|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 7'b1110111;
  assign _1609_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11900|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 7'b1110110;
  assign _1610_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11896|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 7'b1110101;
  assign _1611_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11892|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 7'b1110100;
  assign _1612_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11888|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 7'b1110011;
  assign _1613_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11884|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 7'b1110010;
  assign _1614_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11880|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 7'b1110001;
  assign _1615_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11876|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 7'b1110000;
  assign _1616_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11872|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 7'b1101111;
  assign _1617_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11868|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 7'b1101110;
  assign _1618_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11864|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 7'b1101101;
  assign _1619_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11860|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 7'b1101100;
  assign _1620_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11856|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 7'b1101011;
  assign _1621_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11852|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 7'b1101010;
  assign _1622_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11848|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 7'b1101001;
  assign _1623_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11844|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 7'b1101000;
  assign _1624_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11840|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 7'b1100111;
  assign _1625_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11836|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 7'b1100110;
  assign _1626_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11832|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 7'b1100101;
  assign _1627_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11828|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 7'b1100100;
  assign _1628_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11824|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 7'b1100011;
  assign _1629_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11820|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 7'b1100010;
  assign _1630_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11816|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 7'b1100001;
  assign _1631_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11812|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 7'b1100000;
  assign _1632_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11808|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 7'b1011111;
  assign _1633_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11804|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 7'b1011110;
  assign _1634_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11800|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 7'b1011101;
  assign _1635_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11796|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 7'b1011100;
  assign _1636_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11792|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 7'b1011011;
  assign _1637_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11788|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 7'b1011010;
  assign _1638_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11784|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 7'b1011001;
  assign _1639_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11780|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 7'b1011000;
  assign _1640_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11776|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 7'b1010111;
  assign _1641_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11772|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 7'b1010110;
  assign _1642_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11768|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 7'b1010101;
  assign _1643_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11764|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 7'b1010100;
  assign _1644_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11760|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 7'b1010011;
  assign _1645_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11756|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 7'b1010010;
  assign _1646_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11752|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 7'b1010001;
  assign _1647_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11748|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 7'b1010000;
  assign _1648_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11744|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 7'b1001111;
  assign _1649_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11740|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 7'b1001110;
  assign _1650_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11736|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 7'b1001101;
  assign _1651_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11732|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 7'b1001100;
  assign _1652_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11728|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 7'b1001011;
  assign _1653_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11724|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 7'b1001010;
  assign _1654_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11720|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 7'b1001001;
  assign _1655_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11716|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 7'b1001000;
  assign _1656_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11712|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 7'b1000111;
  assign _1657_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11708|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 7'b1000110;
  assign _1658_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11704|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 7'b1000101;
  assign _1659_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11700|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 7'b1000100;
  assign _1660_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11696|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 7'b1000011;
  assign _1661_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11692|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 7'b1000010;
  assign _1662_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11688|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 7'b1000001;
  assign _1663_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11684|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 7'b1000000;
  assign _1664_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11680|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 6'b111111;
  assign _1665_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11676|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 6'b111110;
  assign _1666_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11672|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 6'b111101;
  assign _1667_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11668|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 6'b111100;
  assign _1668_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11664|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 6'b111011;
  assign _1669_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11660|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 6'b111010;
  assign _1670_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11656|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 6'b111001;
  assign _1671_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11652|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 6'b111000;
  assign _1672_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11648|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 6'b110111;
  assign _1673_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11644|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 6'b110110;
  assign _1674_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11640|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 6'b110101;
  assign _1675_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11636|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 6'b110100;
  assign _1676_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11632|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 6'b110011;
  assign _1677_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11628|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 6'b110010;
  assign _1678_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11624|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 6'b110001;
  assign _1679_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11620|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 6'b110000;
  assign _1680_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11616|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 6'b101111;
  assign _1681_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11612|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 6'b101110;
  assign _1682_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11608|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 6'b101101;
  assign _1683_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11604|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 6'b101100;
  assign _1684_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11600|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 6'b101011;
  assign _1685_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11596|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 6'b101010;
  assign _1686_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11592|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 6'b101001;
  assign _1687_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11588|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 6'b101000;
  assign _1688_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11584|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 6'b100111;
  assign _1689_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11580|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 6'b100110;
  assign _1690_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11576|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 6'b100101;
  assign _1691_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11572|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 6'b100100;
  assign _1692_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11568|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 6'b100011;
  assign _1693_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11564|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 6'b100010;
  assign _1694_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11560|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 6'b100001;
  assign _1695_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11556|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 6'b100000;
  assign _1696_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11552|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 5'b11111;
  assign _1697_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11548|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 5'b11110;
  assign _1698_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11544|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 5'b11101;
  assign _1699_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11540|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 5'b11100;
  assign _1700_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11536|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 5'b11011;
  assign _1701_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11532|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 5'b11010;
  assign _1702_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11528|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 5'b11001;
  assign _1703_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11524|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 5'b11000;
  assign _1704_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11520|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 5'b10111;
  assign _1705_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11516|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 5'b10110;
  assign _1706_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11512|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 5'b10101;
  assign _1707_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11508|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 5'b10100;
  assign _1708_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11504|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 5'b10011;
  assign _1709_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11500|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 5'b10010;
  assign _1710_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11496|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 5'b10001;
  assign _1711_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11492|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 5'b10000;
  assign _1712_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11488|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 4'b1111;
  assign _1713_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11484|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 4'b1110;
  assign _1714_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11480|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 4'b1101;
  assign _1715_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11476|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 4'b1100;
  assign _1716_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11472|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 4'b1011;
  assign _1717_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11468|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 4'b1010;
  assign _1718_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11464|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 4'b1001;
  assign _1719_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11460|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 4'b1000;
  assign _1720_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11456|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 3'b111;
  assign _1721_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11452|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 3'b110;
  assign _1722_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11448|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 3'b101;
  assign _1723_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11444|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 3'b100;
  assign _1724_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11440|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 2'b11;
  assign _1725_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11436|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 2'b10;
  assign _1726_ = dp2lut_Y_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11432|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) 1'b1;
  assign _1727_ = ! (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11428|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *) dp2lut_Y_entry_4;
  assign _1728_ = dp2lut_Yinfo_4[17] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11423" *) density_reg256 : _1470_;
  assign _1729_ = dp2lut_Yinfo_4[16] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11420" *) density_reg0 : _1728_;
  assign _0294_ = _0387_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11419" *) _1729_ : lut_Y_data_41;
  function [15:0] _5580_;
    input [15:0] a;
    input [4095:0] b;
    input [255:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:12452|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11427" *)
    (* parallel_case *)
    casez (s)
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1:
        _5580_ = b[15:0];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?:
        _5580_ = b[31:16];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??:
        _5580_ = b[47:32];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???:
        _5580_ = b[63:48];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????:
        _5580_ = b[79:64];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????:
        _5580_ = b[95:80];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????:
        _5580_ = b[111:96];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????:
        _5580_ = b[127:112];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????:
        _5580_ = b[143:128];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????:
        _5580_ = b[159:144];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????:
        _5580_ = b[175:160];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????:
        _5580_ = b[191:176];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????:
        _5580_ = b[207:192];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????:
        _5580_ = b[223:208];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????:
        _5580_ = b[239:224];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????:
        _5580_ = b[255:240];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????:
        _5580_ = b[271:256];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????:
        _5580_ = b[287:272];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????:
        _5580_ = b[303:288];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????:
        _5580_ = b[319:304];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????:
        _5580_ = b[335:320];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????:
        _5580_ = b[351:336];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????:
        _5580_ = b[367:352];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????:
        _5580_ = b[383:368];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????:
        _5580_ = b[399:384];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????:
        _5580_ = b[415:400];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????:
        _5580_ = b[431:416];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????:
        _5580_ = b[447:432];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????:
        _5580_ = b[463:448];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????:
        _5580_ = b[479:464];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????:
        _5580_ = b[495:480];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????:
        _5580_ = b[511:496];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????:
        _5580_ = b[527:512];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????:
        _5580_ = b[543:528];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????:
        _5580_ = b[559:544];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????:
        _5580_ = b[575:560];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????:
        _5580_ = b[591:576];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????:
        _5580_ = b[607:592];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????:
        _5580_ = b[623:608];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????:
        _5580_ = b[639:624];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????:
        _5580_ = b[655:640];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????:
        _5580_ = b[671:656];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????:
        _5580_ = b[687:672];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????:
        _5580_ = b[703:688];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????:
        _5580_ = b[719:704];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????:
        _5580_ = b[735:720];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????:
        _5580_ = b[751:736];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????:
        _5580_ = b[767:752];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????:
        _5580_ = b[783:768];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????:
        _5580_ = b[799:784];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????:
        _5580_ = b[815:800];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????:
        _5580_ = b[831:816];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????:
        _5580_ = b[847:832];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????:
        _5580_ = b[863:848];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????:
        _5580_ = b[879:864];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????:
        _5580_ = b[895:880];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????:
        _5580_ = b[911:896];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????:
        _5580_ = b[927:912];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????:
        _5580_ = b[943:928];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????:
        _5580_ = b[959:944];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????:
        _5580_ = b[975:960];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????:
        _5580_ = b[991:976];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????:
        _5580_ = b[1007:992];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????:
        _5580_ = b[1023:1008];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????:
        _5580_ = b[1039:1024];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????:
        _5580_ = b[1055:1040];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????:
        _5580_ = b[1071:1056];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????:
        _5580_ = b[1087:1072];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????:
        _5580_ = b[1103:1088];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????:
        _5580_ = b[1119:1104];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????:
        _5580_ = b[1135:1120];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????:
        _5580_ = b[1151:1136];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????:
        _5580_ = b[1167:1152];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????:
        _5580_ = b[1183:1168];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????:
        _5580_ = b[1199:1184];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????:
        _5580_ = b[1215:1200];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????:
        _5580_ = b[1231:1216];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????:
        _5580_ = b[1247:1232];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????:
        _5580_ = b[1263:1248];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????:
        _5580_ = b[1279:1264];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????:
        _5580_ = b[1295:1280];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????:
        _5580_ = b[1311:1296];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????:
        _5580_ = b[1327:1312];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????:
        _5580_ = b[1343:1328];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????:
        _5580_ = b[1359:1344];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????:
        _5580_ = b[1375:1360];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????:
        _5580_ = b[1391:1376];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????:
        _5580_ = b[1407:1392];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????:
        _5580_ = b[1423:1408];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????:
        _5580_ = b[1439:1424];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????:
        _5580_ = b[1455:1440];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????:
        _5580_ = b[1471:1456];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????:
        _5580_ = b[1487:1472];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????:
        _5580_ = b[1503:1488];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????:
        _5580_ = b[1519:1504];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????:
        _5580_ = b[1535:1520];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????:
        _5580_ = b[1551:1536];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????:
        _5580_ = b[1567:1552];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????:
        _5580_ = b[1583:1568];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????:
        _5580_ = b[1599:1584];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5580_ = b[1615:1600];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5580_ = b[1631:1616];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5580_ = b[1647:1632];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5580_ = b[1663:1648];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5580_ = b[1679:1664];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5580_ = b[1695:1680];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5580_ = b[1711:1696];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5580_ = b[1727:1712];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5580_ = b[1743:1728];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5580_ = b[1759:1744];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5580_ = b[1775:1760];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5580_ = b[1791:1776];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5580_ = b[1807:1792];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5580_ = b[1823:1808];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5580_ = b[1839:1824];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5580_ = b[1855:1840];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5580_ = b[1871:1856];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5580_ = b[1887:1872];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5580_ = b[1903:1888];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5580_ = b[1919:1904];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5580_ = b[1935:1920];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5580_ = b[1951:1936];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5580_ = b[1967:1952];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5580_ = b[1983:1968];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5580_ = b[1999:1984];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5580_ = b[2015:2000];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5580_ = b[2031:2016];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5580_ = b[2047:2032];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5580_ = b[2063:2048];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5580_ = b[2079:2064];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5580_ = b[2095:2080];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5580_ = b[2111:2096];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5580_ = b[2127:2112];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5580_ = b[2143:2128];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5580_ = b[2159:2144];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5580_ = b[2175:2160];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5580_ = b[2191:2176];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5580_ = b[2207:2192];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5580_ = b[2223:2208];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5580_ = b[2239:2224];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5580_ = b[2255:2240];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5580_ = b[2271:2256];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5580_ = b[2287:2272];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5580_ = b[2303:2288];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5580_ = b[2319:2304];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5580_ = b[2335:2320];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5580_ = b[2351:2336];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5580_ = b[2367:2352];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5580_ = b[2383:2368];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5580_ = b[2399:2384];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5580_ = b[2415:2400];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5580_ = b[2431:2416];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5580_ = b[2447:2432];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5580_ = b[2463:2448];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5580_ = b[2479:2464];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5580_ = b[2495:2480];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5580_ = b[2511:2496];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5580_ = b[2527:2512];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5580_ = b[2543:2528];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5580_ = b[2559:2544];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5580_ = b[2575:2560];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5580_ = b[2591:2576];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5580_ = b[2607:2592];
      256'b????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5580_ = b[2623:2608];
      256'b???????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5580_ = b[2639:2624];
      256'b??????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5580_ = b[2655:2640];
      256'b?????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5580_ = b[2671:2656];
      256'b????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5580_ = b[2687:2672];
      256'b???????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5580_ = b[2703:2688];
      256'b??????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5580_ = b[2719:2704];
      256'b?????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5580_ = b[2735:2720];
      256'b????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5580_ = b[2751:2736];
      256'b???????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5580_ = b[2767:2752];
      256'b??????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5580_ = b[2783:2768];
      256'b?????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5580_ = b[2799:2784];
      256'b????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5580_ = b[2815:2800];
      256'b???????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5580_ = b[2831:2816];
      256'b??????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5580_ = b[2847:2832];
      256'b?????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5580_ = b[2863:2848];
      256'b????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5580_ = b[2879:2864];
      256'b???????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5580_ = b[2895:2880];
      256'b??????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5580_ = b[2911:2896];
      256'b?????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5580_ = b[2927:2912];
      256'b????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5580_ = b[2943:2928];
      256'b???????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5580_ = b[2959:2944];
      256'b??????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5580_ = b[2975:2960];
      256'b?????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5580_ = b[2991:2976];
      256'b????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5580_ = b[3007:2992];
      256'b???????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5580_ = b[3023:3008];
      256'b??????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5580_ = b[3039:3024];
      256'b?????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5580_ = b[3055:3040];
      256'b????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5580_ = b[3071:3056];
      256'b???????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5580_ = b[3087:3072];
      256'b??????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5580_ = b[3103:3088];
      256'b?????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5580_ = b[3119:3104];
      256'b????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5580_ = b[3135:3120];
      256'b???????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5580_ = b[3151:3136];
      256'b??????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5580_ = b[3167:3152];
      256'b?????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5580_ = b[3183:3168];
      256'b????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5580_ = b[3199:3184];
      256'b???????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5580_ = b[3215:3200];
      256'b??????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5580_ = b[3231:3216];
      256'b?????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5580_ = b[3247:3232];
      256'b????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5580_ = b[3263:3248];
      256'b???????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5580_ = b[3279:3264];
      256'b??????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5580_ = b[3295:3280];
      256'b?????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5580_ = b[3311:3296];
      256'b????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5580_ = b[3327:3312];
      256'b???????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5580_ = b[3343:3328];
      256'b??????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5580_ = b[3359:3344];
      256'b?????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5580_ = b[3375:3360];
      256'b????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5580_ = b[3391:3376];
      256'b???????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5580_ = b[3407:3392];
      256'b??????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5580_ = b[3423:3408];
      256'b?????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5580_ = b[3439:3424];
      256'b????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5580_ = b[3455:3440];
      256'b???????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5580_ = b[3471:3456];
      256'b??????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5580_ = b[3487:3472];
      256'b?????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5580_ = b[3503:3488];
      256'b????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5580_ = b[3519:3504];
      256'b???????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5580_ = b[3535:3520];
      256'b??????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5580_ = b[3551:3536];
      256'b?????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5580_ = b[3567:3552];
      256'b????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5580_ = b[3583:3568];
      256'b???????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5580_ = b[3599:3584];
      256'b??????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5580_ = b[3615:3600];
      256'b?????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5580_ = b[3631:3616];
      256'b????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5580_ = b[3647:3632];
      256'b???????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5580_ = b[3663:3648];
      256'b??????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5580_ = b[3679:3664];
      256'b?????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5580_ = b[3695:3680];
      256'b????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5580_ = b[3711:3696];
      256'b???????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5580_ = b[3727:3712];
      256'b??????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5580_ = b[3743:3728];
      256'b?????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5580_ = b[3759:3744];
      256'b????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5580_ = b[3775:3760];
      256'b???????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5580_ = b[3791:3776];
      256'b??????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5580_ = b[3807:3792];
      256'b?????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5580_ = b[3823:3808];
      256'b????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5580_ = b[3839:3824];
      256'b???????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5580_ = b[3855:3840];
      256'b??????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5580_ = b[3871:3856];
      256'b?????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5580_ = b[3887:3872];
      256'b????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5580_ = b[3903:3888];
      256'b???????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5580_ = b[3919:3904];
      256'b??????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5580_ = b[3935:3920];
      256'b?????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5580_ = b[3951:3936];
      256'b????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5580_ = b[3967:3952];
      256'b???????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5580_ = b[3983:3968];
      256'b??????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5580_ = b[3999:3984];
      256'b?????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5580_ = b[4015:4000];
      256'b????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5580_ = b[4031:4016];
      256'b???1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5580_ = b[4047:4032];
      256'b??1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5580_ = b[4063:4048];
      256'b?1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5580_ = b[4079:4064];
      256'b1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5580_ = b[4095:4080];
      default:
        _5580_ = a;
    endcase
  endfunction
  assign _1730_ = _5580_(density_reg0, { density_reg1, density_reg2, density_reg3, density_reg4, density_reg5, density_reg6, density_reg7, density_reg8, density_reg9, density_reg10, density_reg11, density_reg12, density_reg13, density_reg14, density_reg15, density_reg16, density_reg17, density_reg18, density_reg19, density_reg20, density_reg21, density_reg22, density_reg23, density_reg24, density_reg25, density_reg26, density_reg27, density_reg28, density_reg29, density_reg30, density_reg31, density_reg32, density_reg33, density_reg34, density_reg35, density_reg36, density_reg37, density_reg38, density_reg39, density_reg40, density_reg41, density_reg42, density_reg43, density_reg44, density_reg45, density_reg46, density_reg47, density_reg48, density_reg49, density_reg50, density_reg51, density_reg52, density_reg53, density_reg54, density_reg55, density_reg56, density_reg57, density_reg58, density_reg59, density_reg60, density_reg61, density_reg62, density_reg63, density_reg64, density_reg65, density_reg66, density_reg67, density_reg68, density_reg69, density_reg70, density_reg71, density_reg72, density_reg73, density_reg74, density_reg75, density_reg76, density_reg77, density_reg78, density_reg79, density_reg80, density_reg81, density_reg82, density_reg83, density_reg84, density_reg85, density_reg86, density_reg87, density_reg88, density_reg89, density_reg90, density_reg91, density_reg92, density_reg93, density_reg94, density_reg95, density_reg96, density_reg97, density_reg98, density_reg99, density_reg100, density_reg101, density_reg102, density_reg103, density_reg104, density_reg105, density_reg106, density_reg107, density_reg108, density_reg109, density_reg110, density_reg111, density_reg112, density_reg113, density_reg114, density_reg115, density_reg116, density_reg117, density_reg118, density_reg119, density_reg120, density_reg121, density_reg122, density_reg123, density_reg124, density_reg125, density_reg126, density_reg127, density_reg128, density_reg129, density_reg130, density_reg131, density_reg132, density_reg133, density_reg134, density_reg135, density_reg136, density_reg137, density_reg138, density_reg139, density_reg140, density_reg141, density_reg142, density_reg143, density_reg144, density_reg145, density_reg146, density_reg147, density_reg148, density_reg149, density_reg150, density_reg151, density_reg152, density_reg153, density_reg154, density_reg155, density_reg156, density_reg157, density_reg158, density_reg159, density_reg160, density_reg161, density_reg162, density_reg163, density_reg164, density_reg165, density_reg166, density_reg167, density_reg168, density_reg169, density_reg170, density_reg171, density_reg172, density_reg173, density_reg174, density_reg175, density_reg176, density_reg177, density_reg178, density_reg179, density_reg180, density_reg181, density_reg182, density_reg183, density_reg184, density_reg185, density_reg186, density_reg187, density_reg188, density_reg189, density_reg190, density_reg191, density_reg192, density_reg193, density_reg194, density_reg195, density_reg196, density_reg197, density_reg198, density_reg199, density_reg200, density_reg201, density_reg202, density_reg203, density_reg204, density_reg205, density_reg206, density_reg207, density_reg208, density_reg209, density_reg210, density_reg211, density_reg212, density_reg213, density_reg214, density_reg215, density_reg216, density_reg217, density_reg218, density_reg219, density_reg220, density_reg221, density_reg222, density_reg223, density_reg224, density_reg225, density_reg226, density_reg227, density_reg228, density_reg229, density_reg230, density_reg231, density_reg232, density_reg233, density_reg234, density_reg235, density_reg236, density_reg237, density_reg238, density_reg239, density_reg240, density_reg241, density_reg242, density_reg243, density_reg244, density_reg245, density_reg246, density_reg247, density_reg248, density_reg249, density_reg250, density_reg251, density_reg252, density_reg253, density_reg254, density_reg255, density_reg256 }, { _1726_, _1725_, _1724_, _1723_, _1722_, _1721_, _1720_, _1719_, _1718_, _1717_, _1716_, _1715_, _1714_, _1713_, _1712_, _1711_, _1710_, _1709_, _1708_, _1707_, _1706_, _1705_, _1704_, _1703_, _1702_, _1701_, _1700_, _1699_, _1698_, _1697_, _1696_, _1695_, _1694_, _1693_, _1692_, _1691_, _1690_, _1689_, _1688_, _1687_, _1686_, _1685_, _1684_, _1683_, _1682_, _1681_, _1680_, _1679_, _1678_, _1677_, _1676_, _1675_, _1674_, _1673_, _1672_, _1671_, _1670_, _1669_, _1668_, _1667_, _1666_, _1665_, _1664_, _1663_, _1662_, _1661_, _1660_, _1659_, _1658_, _1657_, _1656_, _1655_, _1654_, _1653_, _1652_, _1651_, _1650_, _1649_, _1648_, _1647_, _1646_, _1645_, _1644_, _1643_, _1642_, _1641_, _1640_, _1639_, _1638_, _1637_, _1636_, _1635_, _1634_, _1633_, _1632_, _1631_, _1630_, _1629_, _1628_, _1627_, _1626_, _1625_, _1624_, _1623_, _1622_, _1621_, _1620_, _1619_, _1618_, _1617_, _1616_, _1615_, _1614_, _1613_, _1612_, _1611_, _1610_, _1609_, _1608_, _1607_, _1606_, _1605_, _1604_, _1603_, _1602_, _1601_, _1600_, _1599_, _1598_, _1597_, _1596_, _1595_, _1594_, _1593_, _1592_, _1591_, _1590_, _1589_, _1588_, _1587_, _1586_, _1585_, _1584_, _1583_, _1582_, _1581_, _1580_, _1579_, _1578_, _1577_, _1576_, _1575_, _1574_, _1573_, _1572_, _1571_, _1570_, _1569_, _1568_, _1567_, _1566_, _1565_, _1564_, _1563_, _1562_, _1561_, _1560_, _1559_, _1558_, _1557_, _1556_, _1555_, _1554_, _1553_, _1552_, _1551_, _1550_, _1549_, _1548_, _1547_, _1546_, _1545_, _1544_, _1543_, _1542_, _1541_, _1540_, _1539_, _1538_, _1537_, _1536_, _1535_, _1534_, _1533_, _1532_, _1531_, _1530_, _1529_, _1528_, _1527_, _1526_, _1525_, _1524_, _1523_, _1522_, _1521_, _1520_, _1519_, _1518_, _1517_, _1516_, _1515_, _1514_, _1513_, _1512_, _1511_, _1510_, _1509_, _1508_, _1507_, _1506_, _1505_, _1504_, _1503_, _1502_, _1501_, _1500_, _1499_, _1498_, _1497_, _1496_, _1495_, _1494_, _1493_, _1492_, _1491_, _1490_, _1489_, _1488_, _1487_, _1486_, _1485_, _1484_, _1483_, _1482_, _1481_, _1480_, _1479_, _1478_, _1477_, _1476_, _1475_, _1474_, _1473_, _1472_, _1471_ });
  assign _1731_ = dp2lut_Yinfo_4[17] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11423" *) density_reg256 : _1730_;
  assign _1732_ = dp2lut_Yinfo_4[16] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11420" *) density_reg0 : _1731_;
  assign _0293_ = _0387_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11419" *) _1732_ : lut_Y_data_40;
  function [15:0] _5584_;
    input [15:0] a;
    input [4095:0] b;
    input [255:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11401|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *)
    (* parallel_case *)
    casez (s)
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1:
        _5584_ = b[15:0];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?:
        _5584_ = b[31:16];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??:
        _5584_ = b[47:32];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???:
        _5584_ = b[63:48];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????:
        _5584_ = b[79:64];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????:
        _5584_ = b[95:80];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????:
        _5584_ = b[111:96];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????:
        _5584_ = b[127:112];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????:
        _5584_ = b[143:128];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????:
        _5584_ = b[159:144];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????:
        _5584_ = b[175:160];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????:
        _5584_ = b[191:176];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????:
        _5584_ = b[207:192];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????:
        _5584_ = b[223:208];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????:
        _5584_ = b[239:224];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????:
        _5584_ = b[255:240];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????:
        _5584_ = b[271:256];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????:
        _5584_ = b[287:272];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????:
        _5584_ = b[303:288];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????:
        _5584_ = b[319:304];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????:
        _5584_ = b[335:320];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????:
        _5584_ = b[351:336];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????:
        _5584_ = b[367:352];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????:
        _5584_ = b[383:368];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????:
        _5584_ = b[399:384];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????:
        _5584_ = b[415:400];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????:
        _5584_ = b[431:416];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????:
        _5584_ = b[447:432];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????:
        _5584_ = b[463:448];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????:
        _5584_ = b[479:464];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????:
        _5584_ = b[495:480];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????:
        _5584_ = b[511:496];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????:
        _5584_ = b[527:512];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????:
        _5584_ = b[543:528];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????:
        _5584_ = b[559:544];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????:
        _5584_ = b[575:560];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????:
        _5584_ = b[591:576];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????:
        _5584_ = b[607:592];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????:
        _5584_ = b[623:608];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????:
        _5584_ = b[639:624];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????:
        _5584_ = b[655:640];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????:
        _5584_ = b[671:656];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????:
        _5584_ = b[687:672];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????:
        _5584_ = b[703:688];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????:
        _5584_ = b[719:704];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????:
        _5584_ = b[735:720];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????:
        _5584_ = b[751:736];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????:
        _5584_ = b[767:752];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????:
        _5584_ = b[783:768];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????:
        _5584_ = b[799:784];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????:
        _5584_ = b[815:800];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????:
        _5584_ = b[831:816];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????:
        _5584_ = b[847:832];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????:
        _5584_ = b[863:848];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????:
        _5584_ = b[879:864];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????:
        _5584_ = b[895:880];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????:
        _5584_ = b[911:896];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????:
        _5584_ = b[927:912];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????:
        _5584_ = b[943:928];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????:
        _5584_ = b[959:944];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????:
        _5584_ = b[975:960];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????:
        _5584_ = b[991:976];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????:
        _5584_ = b[1007:992];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????:
        _5584_ = b[1023:1008];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????:
        _5584_ = b[1039:1024];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????:
        _5584_ = b[1055:1040];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????:
        _5584_ = b[1071:1056];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????:
        _5584_ = b[1087:1072];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????:
        _5584_ = b[1103:1088];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????:
        _5584_ = b[1119:1104];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????:
        _5584_ = b[1135:1120];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????:
        _5584_ = b[1151:1136];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????:
        _5584_ = b[1167:1152];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????:
        _5584_ = b[1183:1168];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????:
        _5584_ = b[1199:1184];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????:
        _5584_ = b[1215:1200];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????:
        _5584_ = b[1231:1216];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????:
        _5584_ = b[1247:1232];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????:
        _5584_ = b[1263:1248];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????:
        _5584_ = b[1279:1264];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????:
        _5584_ = b[1295:1280];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????:
        _5584_ = b[1311:1296];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????:
        _5584_ = b[1327:1312];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????:
        _5584_ = b[1343:1328];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????:
        _5584_ = b[1359:1344];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????:
        _5584_ = b[1375:1360];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????:
        _5584_ = b[1391:1376];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????:
        _5584_ = b[1407:1392];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????:
        _5584_ = b[1423:1408];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????:
        _5584_ = b[1439:1424];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????:
        _5584_ = b[1455:1440];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????:
        _5584_ = b[1471:1456];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????:
        _5584_ = b[1487:1472];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????:
        _5584_ = b[1503:1488];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????:
        _5584_ = b[1519:1504];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????:
        _5584_ = b[1535:1520];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????:
        _5584_ = b[1551:1536];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????:
        _5584_ = b[1567:1552];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????:
        _5584_ = b[1583:1568];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????:
        _5584_ = b[1599:1584];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5584_ = b[1615:1600];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5584_ = b[1631:1616];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5584_ = b[1647:1632];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5584_ = b[1663:1648];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5584_ = b[1679:1664];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5584_ = b[1695:1680];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5584_ = b[1711:1696];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5584_ = b[1727:1712];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5584_ = b[1743:1728];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5584_ = b[1759:1744];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5584_ = b[1775:1760];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5584_ = b[1791:1776];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5584_ = b[1807:1792];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5584_ = b[1823:1808];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5584_ = b[1839:1824];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5584_ = b[1855:1840];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5584_ = b[1871:1856];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5584_ = b[1887:1872];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5584_ = b[1903:1888];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5584_ = b[1919:1904];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5584_ = b[1935:1920];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5584_ = b[1951:1936];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5584_ = b[1967:1952];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5584_ = b[1983:1968];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5584_ = b[1999:1984];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5584_ = b[2015:2000];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5584_ = b[2031:2016];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5584_ = b[2047:2032];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5584_ = b[2063:2048];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5584_ = b[2079:2064];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5584_ = b[2095:2080];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5584_ = b[2111:2096];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5584_ = b[2127:2112];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5584_ = b[2143:2128];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5584_ = b[2159:2144];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5584_ = b[2175:2160];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5584_ = b[2191:2176];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5584_ = b[2207:2192];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5584_ = b[2223:2208];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5584_ = b[2239:2224];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5584_ = b[2255:2240];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5584_ = b[2271:2256];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5584_ = b[2287:2272];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5584_ = b[2303:2288];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5584_ = b[2319:2304];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5584_ = b[2335:2320];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5584_ = b[2351:2336];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5584_ = b[2367:2352];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5584_ = b[2383:2368];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5584_ = b[2399:2384];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5584_ = b[2415:2400];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5584_ = b[2431:2416];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5584_ = b[2447:2432];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5584_ = b[2463:2448];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5584_ = b[2479:2464];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5584_ = b[2495:2480];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5584_ = b[2511:2496];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5584_ = b[2527:2512];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5584_ = b[2543:2528];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5584_ = b[2559:2544];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5584_ = b[2575:2560];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5584_ = b[2591:2576];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5584_ = b[2607:2592];
      256'b????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5584_ = b[2623:2608];
      256'b???????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5584_ = b[2639:2624];
      256'b??????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5584_ = b[2655:2640];
      256'b?????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5584_ = b[2671:2656];
      256'b????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5584_ = b[2687:2672];
      256'b???????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5584_ = b[2703:2688];
      256'b??????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5584_ = b[2719:2704];
      256'b?????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5584_ = b[2735:2720];
      256'b????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5584_ = b[2751:2736];
      256'b???????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5584_ = b[2767:2752];
      256'b??????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5584_ = b[2783:2768];
      256'b?????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5584_ = b[2799:2784];
      256'b????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5584_ = b[2815:2800];
      256'b???????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5584_ = b[2831:2816];
      256'b??????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5584_ = b[2847:2832];
      256'b?????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5584_ = b[2863:2848];
      256'b????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5584_ = b[2879:2864];
      256'b???????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5584_ = b[2895:2880];
      256'b??????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5584_ = b[2911:2896];
      256'b?????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5584_ = b[2927:2912];
      256'b????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5584_ = b[2943:2928];
      256'b???????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5584_ = b[2959:2944];
      256'b??????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5584_ = b[2975:2960];
      256'b?????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5584_ = b[2991:2976];
      256'b????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5584_ = b[3007:2992];
      256'b???????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5584_ = b[3023:3008];
      256'b??????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5584_ = b[3039:3024];
      256'b?????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5584_ = b[3055:3040];
      256'b????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5584_ = b[3071:3056];
      256'b???????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5584_ = b[3087:3072];
      256'b??????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5584_ = b[3103:3088];
      256'b?????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5584_ = b[3119:3104];
      256'b????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5584_ = b[3135:3120];
      256'b???????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5584_ = b[3151:3136];
      256'b??????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5584_ = b[3167:3152];
      256'b?????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5584_ = b[3183:3168];
      256'b????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5584_ = b[3199:3184];
      256'b???????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5584_ = b[3215:3200];
      256'b??????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5584_ = b[3231:3216];
      256'b?????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5584_ = b[3247:3232];
      256'b????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5584_ = b[3263:3248];
      256'b???????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5584_ = b[3279:3264];
      256'b??????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5584_ = b[3295:3280];
      256'b?????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5584_ = b[3311:3296];
      256'b????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5584_ = b[3327:3312];
      256'b???????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5584_ = b[3343:3328];
      256'b??????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5584_ = b[3359:3344];
      256'b?????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5584_ = b[3375:3360];
      256'b????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5584_ = b[3391:3376];
      256'b???????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5584_ = b[3407:3392];
      256'b??????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5584_ = b[3423:3408];
      256'b?????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5584_ = b[3439:3424];
      256'b????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5584_ = b[3455:3440];
      256'b???????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5584_ = b[3471:3456];
      256'b??????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5584_ = b[3487:3472];
      256'b?????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5584_ = b[3503:3488];
      256'b????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5584_ = b[3519:3504];
      256'b???????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5584_ = b[3535:3520];
      256'b??????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5584_ = b[3551:3536];
      256'b?????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5584_ = b[3567:3552];
      256'b????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5584_ = b[3583:3568];
      256'b???????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5584_ = b[3599:3584];
      256'b??????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5584_ = b[3615:3600];
      256'b?????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5584_ = b[3631:3616];
      256'b????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5584_ = b[3647:3632];
      256'b???????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5584_ = b[3663:3648];
      256'b??????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5584_ = b[3679:3664];
      256'b?????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5584_ = b[3695:3680];
      256'b????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5584_ = b[3711:3696];
      256'b???????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5584_ = b[3727:3712];
      256'b??????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5584_ = b[3743:3728];
      256'b?????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5584_ = b[3759:3744];
      256'b????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5584_ = b[3775:3760];
      256'b???????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5584_ = b[3791:3776];
      256'b??????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5584_ = b[3807:3792];
      256'b?????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5584_ = b[3823:3808];
      256'b????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5584_ = b[3839:3824];
      256'b???????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5584_ = b[3855:3840];
      256'b??????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5584_ = b[3871:3856];
      256'b?????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5584_ = b[3887:3872];
      256'b????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5584_ = b[3903:3888];
      256'b???????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5584_ = b[3919:3904];
      256'b??????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5584_ = b[3935:3920];
      256'b?????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5584_ = b[3951:3936];
      256'b????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5584_ = b[3967:3952];
      256'b???????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5584_ = b[3983:3968];
      256'b??????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5584_ = b[3999:3984];
      256'b?????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5584_ = b[4015:4000];
      256'b????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5584_ = b[4031:4016];
      256'b???1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5584_ = b[4047:4032];
      256'b??1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5584_ = b[4063:4048];
      256'b?1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5584_ = b[4079:4064];
      256'b1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5584_ = b[4095:4080];
      default:
        _5584_ = a;
    endcase
  endfunction
  assign _1733_ = _5584_(density_reg0, { density_reg1, density_reg2, density_reg3, density_reg4, density_reg5, density_reg6, density_reg7, density_reg8, density_reg9, density_reg10, density_reg11, density_reg12, density_reg13, density_reg14, density_reg15, density_reg16, density_reg17, density_reg18, density_reg19, density_reg20, density_reg21, density_reg22, density_reg23, density_reg24, density_reg25, density_reg26, density_reg27, density_reg28, density_reg29, density_reg30, density_reg31, density_reg32, density_reg33, density_reg34, density_reg35, density_reg36, density_reg37, density_reg38, density_reg39, density_reg40, density_reg41, density_reg42, density_reg43, density_reg44, density_reg45, density_reg46, density_reg47, density_reg48, density_reg49, density_reg50, density_reg51, density_reg52, density_reg53, density_reg54, density_reg55, density_reg56, density_reg57, density_reg58, density_reg59, density_reg60, density_reg61, density_reg62, density_reg63, density_reg64, density_reg65, density_reg66, density_reg67, density_reg68, density_reg69, density_reg70, density_reg71, density_reg72, density_reg73, density_reg74, density_reg75, density_reg76, density_reg77, density_reg78, density_reg79, density_reg80, density_reg81, density_reg82, density_reg83, density_reg84, density_reg85, density_reg86, density_reg87, density_reg88, density_reg89, density_reg90, density_reg91, density_reg92, density_reg93, density_reg94, density_reg95, density_reg96, density_reg97, density_reg98, density_reg99, density_reg100, density_reg101, density_reg102, density_reg103, density_reg104, density_reg105, density_reg106, density_reg107, density_reg108, density_reg109, density_reg110, density_reg111, density_reg112, density_reg113, density_reg114, density_reg115, density_reg116, density_reg117, density_reg118, density_reg119, density_reg120, density_reg121, density_reg122, density_reg123, density_reg124, density_reg125, density_reg126, density_reg127, density_reg128, density_reg129, density_reg130, density_reg131, density_reg132, density_reg133, density_reg134, density_reg135, density_reg136, density_reg137, density_reg138, density_reg139, density_reg140, density_reg141, density_reg142, density_reg143, density_reg144, density_reg145, density_reg146, density_reg147, density_reg148, density_reg149, density_reg150, density_reg151, density_reg152, density_reg153, density_reg154, density_reg155, density_reg156, density_reg157, density_reg158, density_reg159, density_reg160, density_reg161, density_reg162, density_reg163, density_reg164, density_reg165, density_reg166, density_reg167, density_reg168, density_reg169, density_reg170, density_reg171, density_reg172, density_reg173, density_reg174, density_reg175, density_reg176, density_reg177, density_reg178, density_reg179, density_reg180, density_reg181, density_reg182, density_reg183, density_reg184, density_reg185, density_reg186, density_reg187, density_reg188, density_reg189, density_reg190, density_reg191, density_reg192, density_reg193, density_reg194, density_reg195, density_reg196, density_reg197, density_reg198, density_reg199, density_reg200, density_reg201, density_reg202, density_reg203, density_reg204, density_reg205, density_reg206, density_reg207, density_reg208, density_reg209, density_reg210, density_reg211, density_reg212, density_reg213, density_reg214, density_reg215, density_reg216, density_reg217, density_reg218, density_reg219, density_reg220, density_reg221, density_reg222, density_reg223, density_reg224, density_reg225, density_reg226, density_reg227, density_reg228, density_reg229, density_reg230, density_reg231, density_reg232, density_reg233, density_reg234, density_reg235, density_reg236, density_reg237, density_reg238, density_reg239, density_reg240, density_reg241, density_reg242, density_reg243, density_reg244, density_reg245, density_reg246, density_reg247, density_reg248, density_reg249, density_reg250, density_reg251, density_reg252, density_reg253, density_reg254, density_reg255, density_reg256 }, { _1990_, _1989_, _1988_, _1987_, _1986_, _1985_, _1984_, _1983_, _1982_, _1981_, _1980_, _1979_, _1978_, _1977_, _1976_, _1975_, _1974_, _1973_, _1972_, _1971_, _1970_, _1969_, _1968_, _1967_, _1966_, _1965_, _1964_, _1963_, _1962_, _1961_, _1960_, _1959_, _1958_, _1957_, _1956_, _1955_, _1954_, _1953_, _1952_, _1951_, _1950_, _1949_, _1948_, _1947_, _1946_, _1945_, _1944_, _1943_, _1942_, _1941_, _1940_, _1939_, _1938_, _1937_, _1936_, _1935_, _1934_, _1933_, _1932_, _1931_, _1930_, _1929_, _1928_, _1927_, _1926_, _1925_, _1924_, _1923_, _1922_, _1921_, _1920_, _1919_, _1918_, _1917_, _1916_, _1915_, _1914_, _1913_, _1912_, _1911_, _1910_, _1909_, _1908_, _1907_, _1906_, _1905_, _1904_, _1903_, _1902_, _1901_, _1900_, _1899_, _1898_, _1897_, _1896_, _1895_, _1894_, _1893_, _1892_, _1891_, _1890_, _1889_, _1888_, _1887_, _1886_, _1885_, _1884_, _1883_, _1882_, _1881_, _1880_, _1879_, _1878_, _1877_, _1876_, _1875_, _1874_, _1873_, _1872_, _1871_, _1870_, _1869_, _1868_, _1867_, _1866_, _1865_, _1864_, _1863_, _1862_, _1861_, _1860_, _1859_, _1858_, _1857_, _1856_, _1855_, _1854_, _1853_, _1852_, _1851_, _1850_, _1849_, _1848_, _1847_, _1846_, _1845_, _1844_, _1843_, _1842_, _1841_, _1840_, _1839_, _1838_, _1837_, _1836_, _1835_, _1834_, _1833_, _1832_, _1831_, _1830_, _1829_, _1828_, _1827_, _1826_, _1825_, _1824_, _1823_, _1822_, _1821_, _1820_, _1819_, _1818_, _1817_, _1816_, _1815_, _1814_, _1813_, _1812_, _1811_, _1810_, _1809_, _1808_, _1807_, _1806_, _1805_, _1804_, _1803_, _1802_, _1801_, _1800_, _1799_, _1798_, _1797_, _1796_, _1795_, _1794_, _1793_, _1792_, _1791_, _1790_, _1789_, _1788_, _1787_, _1786_, _1785_, _1784_, _1783_, _1782_, _1781_, _1780_, _1779_, _1778_, _1777_, _1776_, _1775_, _1774_, _1773_, _1772_, _1771_, _1770_, _1769_, _1768_, _1767_, _1766_, _1765_, _1764_, _1763_, _1762_, _1761_, _1760_, _1759_, _1758_, _1757_, _1756_, _1755_, _1754_, _1753_, _1752_, _1751_, _1750_, _1749_, _1748_, _1747_, _1746_, _1745_, _1744_, _1743_, _1742_, _1741_, _1740_, _1739_, _1738_, _1737_, _1736_, _0418_ });
  assign _1734_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11401|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 9'b100000000;
  assign _1735_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11397|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 8'b11111111;
  assign _1736_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11393|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 8'b11111110;
  assign _1737_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11389|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 8'b11111101;
  assign _1738_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11385|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 8'b11111100;
  assign _1739_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11381|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 8'b11111011;
  assign _1740_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11377|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 8'b11111010;
  assign _1741_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11373|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 8'b11111001;
  assign _1742_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11369|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 8'b11111000;
  assign _1743_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11365|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 8'b11110111;
  assign _1744_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11361|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 8'b11110110;
  assign _1745_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11357|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 8'b11110101;
  assign _1746_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11353|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 8'b11110100;
  assign _1747_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11349|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 8'b11110011;
  assign _1748_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11345|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 8'b11110010;
  assign _1749_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11341|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 8'b11110001;
  assign _1750_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11337|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 8'b11110000;
  assign _1751_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11333|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 8'b11101111;
  assign _1752_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11329|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 8'b11101110;
  assign _1753_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11325|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 8'b11101101;
  assign _1754_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11321|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 8'b11101100;
  assign _1755_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11317|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 8'b11101011;
  assign _1756_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11313|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 8'b11101010;
  assign _1757_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11309|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 8'b11101001;
  assign _1758_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11305|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 8'b11101000;
  assign _1759_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11301|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 8'b11100111;
  assign _1760_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11297|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 8'b11100110;
  assign _1761_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11293|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 8'b11100101;
  assign _1762_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11289|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 8'b11100100;
  assign _1763_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11285|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 8'b11100011;
  assign _1764_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11281|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 8'b11100010;
  assign _1765_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11277|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 8'b11100001;
  assign _1766_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11273|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 8'b11100000;
  assign _1767_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11269|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 8'b11011111;
  assign _1768_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11265|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 8'b11011110;
  assign _1769_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11261|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 8'b11011101;
  assign _1770_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11257|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 8'b11011100;
  assign _1771_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11253|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 8'b11011011;
  assign _1772_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11249|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 8'b11011010;
  assign _1773_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11245|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 8'b11011001;
  assign _1774_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11241|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 8'b11011000;
  assign _1775_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11237|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 8'b11010111;
  assign _1776_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11233|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 8'b11010110;
  assign _1777_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11229|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 8'b11010101;
  assign _1778_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11225|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 8'b11010100;
  assign _1779_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11221|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 8'b11010011;
  assign _1780_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11217|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 8'b11010010;
  assign _1781_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11213|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 8'b11010001;
  assign _1782_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11209|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 8'b11010000;
  assign _1783_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11205|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 8'b11001111;
  assign _1784_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11201|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 8'b11001110;
  assign _1785_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11197|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 8'b11001101;
  assign _1786_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11193|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 8'b11001100;
  assign _1787_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11189|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 8'b11001011;
  assign _1788_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11185|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 8'b11001010;
  assign _1789_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11181|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 8'b11001001;
  assign _1790_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11177|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 8'b11001000;
  assign _1791_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11173|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 8'b11000111;
  assign _1792_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11169|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 8'b11000110;
  assign _1793_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11165|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 8'b11000101;
  assign _1794_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11161|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 8'b11000100;
  assign _1795_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11157|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 8'b11000011;
  assign _1796_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11153|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 8'b11000010;
  assign _1797_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11149|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 8'b11000001;
  assign _1798_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11145|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 8'b11000000;
  assign _1799_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11141|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 8'b10111111;
  assign _1800_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11137|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 8'b10111110;
  assign _1801_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11133|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 8'b10111101;
  assign _1802_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11129|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 8'b10111100;
  assign _1803_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11125|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 8'b10111011;
  assign _1804_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11121|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 8'b10111010;
  assign _1805_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11117|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 8'b10111001;
  assign _1806_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11113|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 8'b10111000;
  assign _1807_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11109|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 8'b10110111;
  assign _1808_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11105|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 8'b10110110;
  assign _1809_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11101|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 8'b10110101;
  assign _1810_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11097|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 8'b10110100;
  assign _1811_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11093|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 8'b10110011;
  assign _1812_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11089|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 8'b10110010;
  assign _1813_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11085|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 8'b10110001;
  assign _1814_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11081|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 8'b10110000;
  assign _1815_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11077|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 8'b10101111;
  assign _1816_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11073|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 8'b10101110;
  assign _1817_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11069|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 8'b10101101;
  assign _1818_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11065|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 8'b10101100;
  assign _1819_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11061|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 8'b10101011;
  assign _1820_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11057|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 8'b10101010;
  assign _1821_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11053|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 8'b10101001;
  assign _1822_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11049|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 8'b10101000;
  assign _1823_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11045|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 8'b10100111;
  assign _1824_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11041|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 8'b10100110;
  assign _1825_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11037|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 8'b10100101;
  assign _1826_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11033|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 8'b10100100;
  assign _1827_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11029|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 8'b10100011;
  assign _1828_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11025|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 8'b10100010;
  assign _1829_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11021|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 8'b10100001;
  assign _1830_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11017|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 8'b10100000;
  assign _1831_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11013|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 8'b10011111;
  assign _1832_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11009|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 8'b10011110;
  assign _1833_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11005|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 8'b10011101;
  assign _1834_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11001|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 8'b10011100;
  assign _1835_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10997|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 8'b10011011;
  assign _1836_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10993|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 8'b10011010;
  assign _1837_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10989|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 8'b10011001;
  assign _1838_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10985|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 8'b10011000;
  assign _1839_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10981|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 8'b10010111;
  assign _1840_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10977|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 8'b10010110;
  assign _1841_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10973|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 8'b10010101;
  assign _1842_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10969|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 8'b10010100;
  assign _1843_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10965|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 8'b10010011;
  assign _1844_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10961|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 8'b10010010;
  assign _1845_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10957|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 8'b10010001;
  assign _1846_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10953|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 8'b10010000;
  assign _1847_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10949|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 8'b10001111;
  assign _1848_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10945|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 8'b10001110;
  assign _1849_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10941|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 8'b10001101;
  assign _1850_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10937|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 8'b10001100;
  assign _1851_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10933|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 8'b10001011;
  assign _1852_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10929|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 8'b10001010;
  assign _1853_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10925|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 8'b10001001;
  assign _1854_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10921|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 8'b10001000;
  assign _1855_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10917|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 8'b10000111;
  assign _1856_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10913|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 8'b10000110;
  assign _1857_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10909|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 8'b10000101;
  assign _1858_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10905|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 8'b10000100;
  assign _1859_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10901|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 8'b10000011;
  assign _1860_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10897|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 8'b10000010;
  assign _1861_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10893|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 8'b10000001;
  assign _1862_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10889|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 8'b10000000;
  assign _1863_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10885|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 7'b1111111;
  assign _1864_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10881|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 7'b1111110;
  assign _1865_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10877|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 7'b1111101;
  assign _1866_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10873|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 7'b1111100;
  assign _1867_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10869|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 7'b1111011;
  assign _1868_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10865|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 7'b1111010;
  assign _1869_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10861|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 7'b1111001;
  assign _1870_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10857|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 7'b1111000;
  assign _1871_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10853|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 7'b1110111;
  assign _1872_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10849|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 7'b1110110;
  assign _1873_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10845|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 7'b1110101;
  assign _1874_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10841|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 7'b1110100;
  assign _1875_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10837|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 7'b1110011;
  assign _1876_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10833|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 7'b1110010;
  assign _1877_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10829|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 7'b1110001;
  assign _1878_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10825|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 7'b1110000;
  assign _1879_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10821|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 7'b1101111;
  assign _1880_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10817|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 7'b1101110;
  assign _1881_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10813|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 7'b1101101;
  assign _1882_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10809|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 7'b1101100;
  assign _1883_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10805|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 7'b1101011;
  assign _1884_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10801|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 7'b1101010;
  assign _1885_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10797|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 7'b1101001;
  assign _1886_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10793|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 7'b1101000;
  assign _1887_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10789|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 7'b1100111;
  assign _1888_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10785|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 7'b1100110;
  assign _1889_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10781|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 7'b1100101;
  assign _1890_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10777|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 7'b1100100;
  assign _1891_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10773|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 7'b1100011;
  assign _1892_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10769|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 7'b1100010;
  assign _1893_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10765|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 7'b1100001;
  assign _1894_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10761|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 7'b1100000;
  assign _1895_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10757|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 7'b1011111;
  assign _1896_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10753|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 7'b1011110;
  assign _1897_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10749|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 7'b1011101;
  assign _1898_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10745|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 7'b1011100;
  assign _1899_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10741|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 7'b1011011;
  assign _1900_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10737|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 7'b1011010;
  assign _1901_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10733|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 7'b1011001;
  assign _1902_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10729|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 7'b1011000;
  assign _1903_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10725|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 7'b1010111;
  assign _1904_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10721|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 7'b1010110;
  assign _1905_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10717|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 7'b1010101;
  assign _1906_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10713|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 7'b1010100;
  assign _1907_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10709|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 7'b1010011;
  assign _1908_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10705|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 7'b1010010;
  assign _1909_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10701|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 7'b1010001;
  assign _1910_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10697|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 7'b1010000;
  assign _1911_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10693|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 7'b1001111;
  assign _1912_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10689|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 7'b1001110;
  assign _1913_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10685|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 7'b1001101;
  assign _1914_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10681|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 7'b1001100;
  assign _1915_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10677|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 7'b1001011;
  assign _1916_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10673|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 7'b1001010;
  assign _1917_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10669|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 7'b1001001;
  assign _1918_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10665|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 7'b1001000;
  assign _1919_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10661|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 7'b1000111;
  assign _1920_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10657|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 7'b1000110;
  assign _1921_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10653|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 7'b1000101;
  assign _1922_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10649|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 7'b1000100;
  assign _1923_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10645|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 7'b1000011;
  assign _1924_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10641|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 7'b1000010;
  assign _1925_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10637|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 7'b1000001;
  assign _1926_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10633|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 7'b1000000;
  assign _1927_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10629|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 6'b111111;
  assign _1928_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10625|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 6'b111110;
  assign _1929_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10621|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 6'b111101;
  assign _1930_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10617|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 6'b111100;
  assign _1931_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10613|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 6'b111011;
  assign _1932_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10609|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 6'b111010;
  assign _1933_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10605|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 6'b111001;
  assign _1934_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10601|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 6'b111000;
  assign _1935_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10597|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 6'b110111;
  assign _1936_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10593|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 6'b110110;
  assign _1937_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10589|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 6'b110101;
  assign _1938_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10585|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 6'b110100;
  assign _1939_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10581|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 6'b110011;
  assign _1940_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10577|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 6'b110010;
  assign _1941_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10573|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 6'b110001;
  assign _1942_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10569|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 6'b110000;
  assign _1943_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10565|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 6'b101111;
  assign _1944_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10561|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 6'b101110;
  assign _1945_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10557|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 6'b101101;
  assign _1946_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10553|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 6'b101100;
  assign _1947_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10549|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 6'b101011;
  assign _1948_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10545|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 6'b101010;
  assign _1949_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10541|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 6'b101001;
  assign _1950_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10537|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 6'b101000;
  assign _1951_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10533|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 6'b100111;
  assign _1952_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10529|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 6'b100110;
  assign _1953_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10525|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 6'b100101;
  assign _1954_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10521|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 6'b100100;
  assign _1955_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10517|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 6'b100011;
  assign _1956_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10513|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 6'b100010;
  assign _1957_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10509|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 6'b100001;
  assign _1958_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10505|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 6'b100000;
  assign _1959_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10501|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 5'b11111;
  assign _1960_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10497|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 5'b11110;
  assign _1961_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10493|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 5'b11101;
  assign _1962_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10489|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 5'b11100;
  assign _1963_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10485|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 5'b11011;
  assign _1964_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10481|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 5'b11010;
  assign _1965_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10477|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 5'b11001;
  assign _1966_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10473|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 5'b11000;
  assign _1967_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10469|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 5'b10111;
  assign _1968_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10465|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 5'b10110;
  assign _1969_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10461|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 5'b10101;
  assign _1970_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10457|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 5'b10100;
  assign _1971_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10453|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 5'b10011;
  assign _1972_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10449|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 5'b10010;
  assign _1973_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10445|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 5'b10001;
  assign _1974_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10441|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 5'b10000;
  assign _1975_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10437|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 4'b1111;
  assign _1976_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10433|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 4'b1110;
  assign _1977_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10429|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 4'b1101;
  assign _1978_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10425|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 4'b1100;
  assign _1979_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10421|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 4'b1011;
  assign _1980_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10417|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 4'b1010;
  assign _1981_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10413|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 4'b1001;
  assign _1982_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10409|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 4'b1000;
  assign _1983_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10405|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 3'b111;
  assign _1984_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10401|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 3'b110;
  assign _1985_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10397|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 3'b101;
  assign _1986_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10393|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 3'b100;
  assign _1987_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10389|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 2'b11;
  assign _1988_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10385|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 2'b10;
  assign _1989_ = dp2lut_Y_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10381|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) 1'b1;
  assign _1990_ = ! (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10377|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *) dp2lut_Y_entry_3;
  assign _1991_ = dp2lut_Yinfo_3[17] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10372" *) density_reg256 : _1733_;
  assign _1992_ = dp2lut_Yinfo_3[16] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10369" *) density_reg0 : _1991_;
  assign _0292_ = _0385_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10368" *) _1992_ : lut_Y_data_31;
  function [15:0] _5845_;
    input [15:0] a;
    input [4095:0] b;
    input [255:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:11401|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10376" *)
    (* parallel_case *)
    casez (s)
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1:
        _5845_ = b[15:0];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?:
        _5845_ = b[31:16];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??:
        _5845_ = b[47:32];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???:
        _5845_ = b[63:48];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????:
        _5845_ = b[79:64];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????:
        _5845_ = b[95:80];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????:
        _5845_ = b[111:96];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????:
        _5845_ = b[127:112];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????:
        _5845_ = b[143:128];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????:
        _5845_ = b[159:144];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????:
        _5845_ = b[175:160];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????:
        _5845_ = b[191:176];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????:
        _5845_ = b[207:192];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????:
        _5845_ = b[223:208];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????:
        _5845_ = b[239:224];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????:
        _5845_ = b[255:240];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????:
        _5845_ = b[271:256];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????:
        _5845_ = b[287:272];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????:
        _5845_ = b[303:288];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????:
        _5845_ = b[319:304];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????:
        _5845_ = b[335:320];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????:
        _5845_ = b[351:336];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????:
        _5845_ = b[367:352];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????:
        _5845_ = b[383:368];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????:
        _5845_ = b[399:384];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????:
        _5845_ = b[415:400];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????:
        _5845_ = b[431:416];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????:
        _5845_ = b[447:432];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????:
        _5845_ = b[463:448];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????:
        _5845_ = b[479:464];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????:
        _5845_ = b[495:480];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????:
        _5845_ = b[511:496];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????:
        _5845_ = b[527:512];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????:
        _5845_ = b[543:528];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????:
        _5845_ = b[559:544];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????:
        _5845_ = b[575:560];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????:
        _5845_ = b[591:576];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????:
        _5845_ = b[607:592];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????:
        _5845_ = b[623:608];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????:
        _5845_ = b[639:624];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????:
        _5845_ = b[655:640];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????:
        _5845_ = b[671:656];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????:
        _5845_ = b[687:672];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????:
        _5845_ = b[703:688];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????:
        _5845_ = b[719:704];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????:
        _5845_ = b[735:720];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????:
        _5845_ = b[751:736];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????:
        _5845_ = b[767:752];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????:
        _5845_ = b[783:768];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????:
        _5845_ = b[799:784];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????:
        _5845_ = b[815:800];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????:
        _5845_ = b[831:816];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????:
        _5845_ = b[847:832];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????:
        _5845_ = b[863:848];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????:
        _5845_ = b[879:864];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????:
        _5845_ = b[895:880];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????:
        _5845_ = b[911:896];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????:
        _5845_ = b[927:912];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????:
        _5845_ = b[943:928];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????:
        _5845_ = b[959:944];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????:
        _5845_ = b[975:960];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????:
        _5845_ = b[991:976];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????:
        _5845_ = b[1007:992];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????:
        _5845_ = b[1023:1008];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????:
        _5845_ = b[1039:1024];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????:
        _5845_ = b[1055:1040];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????:
        _5845_ = b[1071:1056];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????:
        _5845_ = b[1087:1072];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????:
        _5845_ = b[1103:1088];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????:
        _5845_ = b[1119:1104];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????:
        _5845_ = b[1135:1120];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????:
        _5845_ = b[1151:1136];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????:
        _5845_ = b[1167:1152];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????:
        _5845_ = b[1183:1168];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????:
        _5845_ = b[1199:1184];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????:
        _5845_ = b[1215:1200];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????:
        _5845_ = b[1231:1216];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????:
        _5845_ = b[1247:1232];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????:
        _5845_ = b[1263:1248];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????:
        _5845_ = b[1279:1264];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????:
        _5845_ = b[1295:1280];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????:
        _5845_ = b[1311:1296];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????:
        _5845_ = b[1327:1312];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????:
        _5845_ = b[1343:1328];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????:
        _5845_ = b[1359:1344];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????:
        _5845_ = b[1375:1360];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????:
        _5845_ = b[1391:1376];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????:
        _5845_ = b[1407:1392];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????:
        _5845_ = b[1423:1408];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????:
        _5845_ = b[1439:1424];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????:
        _5845_ = b[1455:1440];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????:
        _5845_ = b[1471:1456];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????:
        _5845_ = b[1487:1472];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????:
        _5845_ = b[1503:1488];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????:
        _5845_ = b[1519:1504];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????:
        _5845_ = b[1535:1520];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????:
        _5845_ = b[1551:1536];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????:
        _5845_ = b[1567:1552];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????:
        _5845_ = b[1583:1568];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????:
        _5845_ = b[1599:1584];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5845_ = b[1615:1600];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5845_ = b[1631:1616];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5845_ = b[1647:1632];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5845_ = b[1663:1648];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5845_ = b[1679:1664];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5845_ = b[1695:1680];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5845_ = b[1711:1696];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5845_ = b[1727:1712];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5845_ = b[1743:1728];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5845_ = b[1759:1744];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5845_ = b[1775:1760];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5845_ = b[1791:1776];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5845_ = b[1807:1792];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5845_ = b[1823:1808];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5845_ = b[1839:1824];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5845_ = b[1855:1840];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5845_ = b[1871:1856];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5845_ = b[1887:1872];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5845_ = b[1903:1888];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5845_ = b[1919:1904];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5845_ = b[1935:1920];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5845_ = b[1951:1936];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5845_ = b[1967:1952];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5845_ = b[1983:1968];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5845_ = b[1999:1984];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5845_ = b[2015:2000];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5845_ = b[2031:2016];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5845_ = b[2047:2032];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5845_ = b[2063:2048];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5845_ = b[2079:2064];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5845_ = b[2095:2080];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5845_ = b[2111:2096];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5845_ = b[2127:2112];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5845_ = b[2143:2128];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5845_ = b[2159:2144];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5845_ = b[2175:2160];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5845_ = b[2191:2176];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5845_ = b[2207:2192];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5845_ = b[2223:2208];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5845_ = b[2239:2224];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5845_ = b[2255:2240];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5845_ = b[2271:2256];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5845_ = b[2287:2272];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5845_ = b[2303:2288];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5845_ = b[2319:2304];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5845_ = b[2335:2320];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5845_ = b[2351:2336];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5845_ = b[2367:2352];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5845_ = b[2383:2368];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5845_ = b[2399:2384];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5845_ = b[2415:2400];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5845_ = b[2431:2416];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5845_ = b[2447:2432];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5845_ = b[2463:2448];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5845_ = b[2479:2464];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5845_ = b[2495:2480];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5845_ = b[2511:2496];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5845_ = b[2527:2512];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5845_ = b[2543:2528];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5845_ = b[2559:2544];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5845_ = b[2575:2560];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5845_ = b[2591:2576];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5845_ = b[2607:2592];
      256'b????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5845_ = b[2623:2608];
      256'b???????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5845_ = b[2639:2624];
      256'b??????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5845_ = b[2655:2640];
      256'b?????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5845_ = b[2671:2656];
      256'b????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5845_ = b[2687:2672];
      256'b???????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5845_ = b[2703:2688];
      256'b??????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5845_ = b[2719:2704];
      256'b?????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5845_ = b[2735:2720];
      256'b????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5845_ = b[2751:2736];
      256'b???????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5845_ = b[2767:2752];
      256'b??????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5845_ = b[2783:2768];
      256'b?????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5845_ = b[2799:2784];
      256'b????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5845_ = b[2815:2800];
      256'b???????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5845_ = b[2831:2816];
      256'b??????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5845_ = b[2847:2832];
      256'b?????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5845_ = b[2863:2848];
      256'b????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5845_ = b[2879:2864];
      256'b???????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5845_ = b[2895:2880];
      256'b??????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5845_ = b[2911:2896];
      256'b?????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5845_ = b[2927:2912];
      256'b????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5845_ = b[2943:2928];
      256'b???????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5845_ = b[2959:2944];
      256'b??????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5845_ = b[2975:2960];
      256'b?????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5845_ = b[2991:2976];
      256'b????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5845_ = b[3007:2992];
      256'b???????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5845_ = b[3023:3008];
      256'b??????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5845_ = b[3039:3024];
      256'b?????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5845_ = b[3055:3040];
      256'b????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5845_ = b[3071:3056];
      256'b???????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5845_ = b[3087:3072];
      256'b??????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5845_ = b[3103:3088];
      256'b?????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5845_ = b[3119:3104];
      256'b????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5845_ = b[3135:3120];
      256'b???????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5845_ = b[3151:3136];
      256'b??????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5845_ = b[3167:3152];
      256'b?????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5845_ = b[3183:3168];
      256'b????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5845_ = b[3199:3184];
      256'b???????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5845_ = b[3215:3200];
      256'b??????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5845_ = b[3231:3216];
      256'b?????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5845_ = b[3247:3232];
      256'b????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5845_ = b[3263:3248];
      256'b???????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5845_ = b[3279:3264];
      256'b??????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5845_ = b[3295:3280];
      256'b?????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5845_ = b[3311:3296];
      256'b????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5845_ = b[3327:3312];
      256'b???????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5845_ = b[3343:3328];
      256'b??????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5845_ = b[3359:3344];
      256'b?????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5845_ = b[3375:3360];
      256'b????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5845_ = b[3391:3376];
      256'b???????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5845_ = b[3407:3392];
      256'b??????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5845_ = b[3423:3408];
      256'b?????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5845_ = b[3439:3424];
      256'b????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5845_ = b[3455:3440];
      256'b???????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5845_ = b[3471:3456];
      256'b??????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5845_ = b[3487:3472];
      256'b?????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5845_ = b[3503:3488];
      256'b????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5845_ = b[3519:3504];
      256'b???????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5845_ = b[3535:3520];
      256'b??????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5845_ = b[3551:3536];
      256'b?????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5845_ = b[3567:3552];
      256'b????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5845_ = b[3583:3568];
      256'b???????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5845_ = b[3599:3584];
      256'b??????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5845_ = b[3615:3600];
      256'b?????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5845_ = b[3631:3616];
      256'b????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5845_ = b[3647:3632];
      256'b???????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5845_ = b[3663:3648];
      256'b??????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5845_ = b[3679:3664];
      256'b?????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5845_ = b[3695:3680];
      256'b????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5845_ = b[3711:3696];
      256'b???????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5845_ = b[3727:3712];
      256'b??????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5845_ = b[3743:3728];
      256'b?????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5845_ = b[3759:3744];
      256'b????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5845_ = b[3775:3760];
      256'b???????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5845_ = b[3791:3776];
      256'b??????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5845_ = b[3807:3792];
      256'b?????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5845_ = b[3823:3808];
      256'b????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5845_ = b[3839:3824];
      256'b???????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5845_ = b[3855:3840];
      256'b??????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5845_ = b[3871:3856];
      256'b?????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5845_ = b[3887:3872];
      256'b????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5845_ = b[3903:3888];
      256'b???????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5845_ = b[3919:3904];
      256'b??????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5845_ = b[3935:3920];
      256'b?????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5845_ = b[3951:3936];
      256'b????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5845_ = b[3967:3952];
      256'b???????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5845_ = b[3983:3968];
      256'b??????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5845_ = b[3999:3984];
      256'b?????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5845_ = b[4015:4000];
      256'b????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5845_ = b[4031:4016];
      256'b???1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5845_ = b[4047:4032];
      256'b??1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5845_ = b[4063:4048];
      256'b?1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5845_ = b[4079:4064];
      256'b1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5845_ = b[4095:4080];
      default:
        _5845_ = a;
    endcase
  endfunction
  assign _1993_ = _5845_(density_reg0, { density_reg1, density_reg2, density_reg3, density_reg4, density_reg5, density_reg6, density_reg7, density_reg8, density_reg9, density_reg10, density_reg11, density_reg12, density_reg13, density_reg14, density_reg15, density_reg16, density_reg17, density_reg18, density_reg19, density_reg20, density_reg21, density_reg22, density_reg23, density_reg24, density_reg25, density_reg26, density_reg27, density_reg28, density_reg29, density_reg30, density_reg31, density_reg32, density_reg33, density_reg34, density_reg35, density_reg36, density_reg37, density_reg38, density_reg39, density_reg40, density_reg41, density_reg42, density_reg43, density_reg44, density_reg45, density_reg46, density_reg47, density_reg48, density_reg49, density_reg50, density_reg51, density_reg52, density_reg53, density_reg54, density_reg55, density_reg56, density_reg57, density_reg58, density_reg59, density_reg60, density_reg61, density_reg62, density_reg63, density_reg64, density_reg65, density_reg66, density_reg67, density_reg68, density_reg69, density_reg70, density_reg71, density_reg72, density_reg73, density_reg74, density_reg75, density_reg76, density_reg77, density_reg78, density_reg79, density_reg80, density_reg81, density_reg82, density_reg83, density_reg84, density_reg85, density_reg86, density_reg87, density_reg88, density_reg89, density_reg90, density_reg91, density_reg92, density_reg93, density_reg94, density_reg95, density_reg96, density_reg97, density_reg98, density_reg99, density_reg100, density_reg101, density_reg102, density_reg103, density_reg104, density_reg105, density_reg106, density_reg107, density_reg108, density_reg109, density_reg110, density_reg111, density_reg112, density_reg113, density_reg114, density_reg115, density_reg116, density_reg117, density_reg118, density_reg119, density_reg120, density_reg121, density_reg122, density_reg123, density_reg124, density_reg125, density_reg126, density_reg127, density_reg128, density_reg129, density_reg130, density_reg131, density_reg132, density_reg133, density_reg134, density_reg135, density_reg136, density_reg137, density_reg138, density_reg139, density_reg140, density_reg141, density_reg142, density_reg143, density_reg144, density_reg145, density_reg146, density_reg147, density_reg148, density_reg149, density_reg150, density_reg151, density_reg152, density_reg153, density_reg154, density_reg155, density_reg156, density_reg157, density_reg158, density_reg159, density_reg160, density_reg161, density_reg162, density_reg163, density_reg164, density_reg165, density_reg166, density_reg167, density_reg168, density_reg169, density_reg170, density_reg171, density_reg172, density_reg173, density_reg174, density_reg175, density_reg176, density_reg177, density_reg178, density_reg179, density_reg180, density_reg181, density_reg182, density_reg183, density_reg184, density_reg185, density_reg186, density_reg187, density_reg188, density_reg189, density_reg190, density_reg191, density_reg192, density_reg193, density_reg194, density_reg195, density_reg196, density_reg197, density_reg198, density_reg199, density_reg200, density_reg201, density_reg202, density_reg203, density_reg204, density_reg205, density_reg206, density_reg207, density_reg208, density_reg209, density_reg210, density_reg211, density_reg212, density_reg213, density_reg214, density_reg215, density_reg216, density_reg217, density_reg218, density_reg219, density_reg220, density_reg221, density_reg222, density_reg223, density_reg224, density_reg225, density_reg226, density_reg227, density_reg228, density_reg229, density_reg230, density_reg231, density_reg232, density_reg233, density_reg234, density_reg235, density_reg236, density_reg237, density_reg238, density_reg239, density_reg240, density_reg241, density_reg242, density_reg243, density_reg244, density_reg245, density_reg246, density_reg247, density_reg248, density_reg249, density_reg250, density_reg251, density_reg252, density_reg253, density_reg254, density_reg255, density_reg256 }, { _1989_, _1988_, _1987_, _1986_, _1985_, _1984_, _1983_, _1982_, _1981_, _1980_, _1979_, _1978_, _1977_, _1976_, _1975_, _1974_, _1973_, _1972_, _1971_, _1970_, _1969_, _1968_, _1967_, _1966_, _1965_, _1964_, _1963_, _1962_, _1961_, _1960_, _1959_, _1958_, _1957_, _1956_, _1955_, _1954_, _1953_, _1952_, _1951_, _1950_, _1949_, _1948_, _1947_, _1946_, _1945_, _1944_, _1943_, _1942_, _1941_, _1940_, _1939_, _1938_, _1937_, _1936_, _1935_, _1934_, _1933_, _1932_, _1931_, _1930_, _1929_, _1928_, _1927_, _1926_, _1925_, _1924_, _1923_, _1922_, _1921_, _1920_, _1919_, _1918_, _1917_, _1916_, _1915_, _1914_, _1913_, _1912_, _1911_, _1910_, _1909_, _1908_, _1907_, _1906_, _1905_, _1904_, _1903_, _1902_, _1901_, _1900_, _1899_, _1898_, _1897_, _1896_, _1895_, _1894_, _1893_, _1892_, _1891_, _1890_, _1889_, _1888_, _1887_, _1886_, _1885_, _1884_, _1883_, _1882_, _1881_, _1880_, _1879_, _1878_, _1877_, _1876_, _1875_, _1874_, _1873_, _1872_, _1871_, _1870_, _1869_, _1868_, _1867_, _1866_, _1865_, _1864_, _1863_, _1862_, _1861_, _1860_, _1859_, _1858_, _1857_, _1856_, _1855_, _1854_, _1853_, _1852_, _1851_, _1850_, _1849_, _1848_, _1847_, _1846_, _1845_, _1844_, _1843_, _1842_, _1841_, _1840_, _1839_, _1838_, _1837_, _1836_, _1835_, _1834_, _1833_, _1832_, _1831_, _1830_, _1829_, _1828_, _1827_, _1826_, _1825_, _1824_, _1823_, _1822_, _1821_, _1820_, _1819_, _1818_, _1817_, _1816_, _1815_, _1814_, _1813_, _1812_, _1811_, _1810_, _1809_, _1808_, _1807_, _1806_, _1805_, _1804_, _1803_, _1802_, _1801_, _1800_, _1799_, _1798_, _1797_, _1796_, _1795_, _1794_, _1793_, _1792_, _1791_, _1790_, _1789_, _1788_, _1787_, _1786_, _1785_, _1784_, _1783_, _1782_, _1781_, _1780_, _1779_, _1778_, _1777_, _1776_, _1775_, _1774_, _1773_, _1772_, _1771_, _1770_, _1769_, _1768_, _1767_, _1766_, _1765_, _1764_, _1763_, _1762_, _1761_, _1760_, _1759_, _1758_, _1757_, _1756_, _1755_, _1754_, _1753_, _1752_, _1751_, _1750_, _1749_, _1748_, _1747_, _1746_, _1745_, _1744_, _1743_, _1742_, _1741_, _1740_, _1739_, _1738_, _1737_, _1736_, _1735_, _1734_ });
  assign _1994_ = dp2lut_Yinfo_3[17] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10372" *) density_reg256 : _1993_;
  assign _1995_ = dp2lut_Yinfo_3[16] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10369" *) density_reg0 : _1994_;
  assign _0291_ = _0385_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10368" *) _1995_ : lut_Y_data_30;
  function [15:0] _5849_;
    input [15:0] a;
    input [4095:0] b;
    input [255:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10350|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *)
    (* parallel_case *)
    casez (s)
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1:
        _5849_ = b[15:0];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?:
        _5849_ = b[31:16];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??:
        _5849_ = b[47:32];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???:
        _5849_ = b[63:48];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????:
        _5849_ = b[79:64];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????:
        _5849_ = b[95:80];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????:
        _5849_ = b[111:96];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????:
        _5849_ = b[127:112];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????:
        _5849_ = b[143:128];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????:
        _5849_ = b[159:144];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????:
        _5849_ = b[175:160];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????:
        _5849_ = b[191:176];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????:
        _5849_ = b[207:192];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????:
        _5849_ = b[223:208];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????:
        _5849_ = b[239:224];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????:
        _5849_ = b[255:240];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????:
        _5849_ = b[271:256];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????:
        _5849_ = b[287:272];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????:
        _5849_ = b[303:288];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????:
        _5849_ = b[319:304];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????:
        _5849_ = b[335:320];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????:
        _5849_ = b[351:336];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????:
        _5849_ = b[367:352];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????:
        _5849_ = b[383:368];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????:
        _5849_ = b[399:384];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????:
        _5849_ = b[415:400];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????:
        _5849_ = b[431:416];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????:
        _5849_ = b[447:432];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????:
        _5849_ = b[463:448];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????:
        _5849_ = b[479:464];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????:
        _5849_ = b[495:480];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????:
        _5849_ = b[511:496];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????:
        _5849_ = b[527:512];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????:
        _5849_ = b[543:528];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????:
        _5849_ = b[559:544];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????:
        _5849_ = b[575:560];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????:
        _5849_ = b[591:576];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????:
        _5849_ = b[607:592];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????:
        _5849_ = b[623:608];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????:
        _5849_ = b[639:624];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????:
        _5849_ = b[655:640];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????:
        _5849_ = b[671:656];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????:
        _5849_ = b[687:672];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????:
        _5849_ = b[703:688];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????:
        _5849_ = b[719:704];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????:
        _5849_ = b[735:720];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????:
        _5849_ = b[751:736];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????:
        _5849_ = b[767:752];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????:
        _5849_ = b[783:768];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????:
        _5849_ = b[799:784];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????:
        _5849_ = b[815:800];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????:
        _5849_ = b[831:816];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????:
        _5849_ = b[847:832];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????:
        _5849_ = b[863:848];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????:
        _5849_ = b[879:864];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????:
        _5849_ = b[895:880];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????:
        _5849_ = b[911:896];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????:
        _5849_ = b[927:912];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????:
        _5849_ = b[943:928];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????:
        _5849_ = b[959:944];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????:
        _5849_ = b[975:960];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????:
        _5849_ = b[991:976];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????:
        _5849_ = b[1007:992];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????:
        _5849_ = b[1023:1008];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????:
        _5849_ = b[1039:1024];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????:
        _5849_ = b[1055:1040];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????:
        _5849_ = b[1071:1056];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????:
        _5849_ = b[1087:1072];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????:
        _5849_ = b[1103:1088];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????:
        _5849_ = b[1119:1104];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????:
        _5849_ = b[1135:1120];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????:
        _5849_ = b[1151:1136];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????:
        _5849_ = b[1167:1152];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????:
        _5849_ = b[1183:1168];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????:
        _5849_ = b[1199:1184];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????:
        _5849_ = b[1215:1200];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????:
        _5849_ = b[1231:1216];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????:
        _5849_ = b[1247:1232];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????:
        _5849_ = b[1263:1248];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????:
        _5849_ = b[1279:1264];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????:
        _5849_ = b[1295:1280];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????:
        _5849_ = b[1311:1296];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????:
        _5849_ = b[1327:1312];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????:
        _5849_ = b[1343:1328];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????:
        _5849_ = b[1359:1344];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????:
        _5849_ = b[1375:1360];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????:
        _5849_ = b[1391:1376];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????:
        _5849_ = b[1407:1392];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????:
        _5849_ = b[1423:1408];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????:
        _5849_ = b[1439:1424];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????:
        _5849_ = b[1455:1440];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????:
        _5849_ = b[1471:1456];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????:
        _5849_ = b[1487:1472];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????:
        _5849_ = b[1503:1488];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????:
        _5849_ = b[1519:1504];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????:
        _5849_ = b[1535:1520];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????:
        _5849_ = b[1551:1536];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????:
        _5849_ = b[1567:1552];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????:
        _5849_ = b[1583:1568];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????:
        _5849_ = b[1599:1584];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5849_ = b[1615:1600];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5849_ = b[1631:1616];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5849_ = b[1647:1632];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5849_ = b[1663:1648];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5849_ = b[1679:1664];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5849_ = b[1695:1680];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5849_ = b[1711:1696];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5849_ = b[1727:1712];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5849_ = b[1743:1728];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5849_ = b[1759:1744];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5849_ = b[1775:1760];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5849_ = b[1791:1776];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5849_ = b[1807:1792];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5849_ = b[1823:1808];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5849_ = b[1839:1824];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5849_ = b[1855:1840];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5849_ = b[1871:1856];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5849_ = b[1887:1872];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5849_ = b[1903:1888];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5849_ = b[1919:1904];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5849_ = b[1935:1920];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5849_ = b[1951:1936];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5849_ = b[1967:1952];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5849_ = b[1983:1968];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5849_ = b[1999:1984];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5849_ = b[2015:2000];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5849_ = b[2031:2016];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5849_ = b[2047:2032];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5849_ = b[2063:2048];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5849_ = b[2079:2064];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5849_ = b[2095:2080];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5849_ = b[2111:2096];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5849_ = b[2127:2112];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5849_ = b[2143:2128];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5849_ = b[2159:2144];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5849_ = b[2175:2160];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5849_ = b[2191:2176];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5849_ = b[2207:2192];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5849_ = b[2223:2208];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5849_ = b[2239:2224];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5849_ = b[2255:2240];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5849_ = b[2271:2256];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5849_ = b[2287:2272];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5849_ = b[2303:2288];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5849_ = b[2319:2304];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5849_ = b[2335:2320];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5849_ = b[2351:2336];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5849_ = b[2367:2352];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5849_ = b[2383:2368];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5849_ = b[2399:2384];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5849_ = b[2415:2400];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5849_ = b[2431:2416];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5849_ = b[2447:2432];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5849_ = b[2463:2448];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5849_ = b[2479:2464];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5849_ = b[2495:2480];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5849_ = b[2511:2496];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5849_ = b[2527:2512];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5849_ = b[2543:2528];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5849_ = b[2559:2544];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5849_ = b[2575:2560];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5849_ = b[2591:2576];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5849_ = b[2607:2592];
      256'b????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5849_ = b[2623:2608];
      256'b???????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5849_ = b[2639:2624];
      256'b??????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5849_ = b[2655:2640];
      256'b?????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5849_ = b[2671:2656];
      256'b????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5849_ = b[2687:2672];
      256'b???????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5849_ = b[2703:2688];
      256'b??????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5849_ = b[2719:2704];
      256'b?????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5849_ = b[2735:2720];
      256'b????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5849_ = b[2751:2736];
      256'b???????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5849_ = b[2767:2752];
      256'b??????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5849_ = b[2783:2768];
      256'b?????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5849_ = b[2799:2784];
      256'b????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5849_ = b[2815:2800];
      256'b???????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5849_ = b[2831:2816];
      256'b??????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5849_ = b[2847:2832];
      256'b?????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5849_ = b[2863:2848];
      256'b????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5849_ = b[2879:2864];
      256'b???????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5849_ = b[2895:2880];
      256'b??????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5849_ = b[2911:2896];
      256'b?????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5849_ = b[2927:2912];
      256'b????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5849_ = b[2943:2928];
      256'b???????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5849_ = b[2959:2944];
      256'b??????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5849_ = b[2975:2960];
      256'b?????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5849_ = b[2991:2976];
      256'b????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5849_ = b[3007:2992];
      256'b???????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5849_ = b[3023:3008];
      256'b??????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5849_ = b[3039:3024];
      256'b?????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5849_ = b[3055:3040];
      256'b????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5849_ = b[3071:3056];
      256'b???????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5849_ = b[3087:3072];
      256'b??????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5849_ = b[3103:3088];
      256'b?????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5849_ = b[3119:3104];
      256'b????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5849_ = b[3135:3120];
      256'b???????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5849_ = b[3151:3136];
      256'b??????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5849_ = b[3167:3152];
      256'b?????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5849_ = b[3183:3168];
      256'b????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5849_ = b[3199:3184];
      256'b???????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5849_ = b[3215:3200];
      256'b??????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5849_ = b[3231:3216];
      256'b?????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5849_ = b[3247:3232];
      256'b????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5849_ = b[3263:3248];
      256'b???????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5849_ = b[3279:3264];
      256'b??????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5849_ = b[3295:3280];
      256'b?????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5849_ = b[3311:3296];
      256'b????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5849_ = b[3327:3312];
      256'b???????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5849_ = b[3343:3328];
      256'b??????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5849_ = b[3359:3344];
      256'b?????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5849_ = b[3375:3360];
      256'b????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5849_ = b[3391:3376];
      256'b???????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5849_ = b[3407:3392];
      256'b??????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5849_ = b[3423:3408];
      256'b?????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5849_ = b[3439:3424];
      256'b????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5849_ = b[3455:3440];
      256'b???????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5849_ = b[3471:3456];
      256'b??????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5849_ = b[3487:3472];
      256'b?????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5849_ = b[3503:3488];
      256'b????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5849_ = b[3519:3504];
      256'b???????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5849_ = b[3535:3520];
      256'b??????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5849_ = b[3551:3536];
      256'b?????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5849_ = b[3567:3552];
      256'b????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5849_ = b[3583:3568];
      256'b???????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5849_ = b[3599:3584];
      256'b??????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5849_ = b[3615:3600];
      256'b?????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5849_ = b[3631:3616];
      256'b????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5849_ = b[3647:3632];
      256'b???????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5849_ = b[3663:3648];
      256'b??????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5849_ = b[3679:3664];
      256'b?????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5849_ = b[3695:3680];
      256'b????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5849_ = b[3711:3696];
      256'b???????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5849_ = b[3727:3712];
      256'b??????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5849_ = b[3743:3728];
      256'b?????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5849_ = b[3759:3744];
      256'b????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5849_ = b[3775:3760];
      256'b???????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5849_ = b[3791:3776];
      256'b??????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5849_ = b[3807:3792];
      256'b?????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5849_ = b[3823:3808];
      256'b????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5849_ = b[3839:3824];
      256'b???????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5849_ = b[3855:3840];
      256'b??????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5849_ = b[3871:3856];
      256'b?????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5849_ = b[3887:3872];
      256'b????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5849_ = b[3903:3888];
      256'b???????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5849_ = b[3919:3904];
      256'b??????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5849_ = b[3935:3920];
      256'b?????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5849_ = b[3951:3936];
      256'b????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5849_ = b[3967:3952];
      256'b???????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5849_ = b[3983:3968];
      256'b??????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5849_ = b[3999:3984];
      256'b?????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5849_ = b[4015:4000];
      256'b????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5849_ = b[4031:4016];
      256'b???1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5849_ = b[4047:4032];
      256'b??1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5849_ = b[4063:4048];
      256'b?1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5849_ = b[4079:4064];
      256'b1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _5849_ = b[4095:4080];
      default:
        _5849_ = a;
    endcase
  endfunction
  assign _1996_ = _5849_(density_reg0, { density_reg1, density_reg2, density_reg3, density_reg4, density_reg5, density_reg6, density_reg7, density_reg8, density_reg9, density_reg10, density_reg11, density_reg12, density_reg13, density_reg14, density_reg15, density_reg16, density_reg17, density_reg18, density_reg19, density_reg20, density_reg21, density_reg22, density_reg23, density_reg24, density_reg25, density_reg26, density_reg27, density_reg28, density_reg29, density_reg30, density_reg31, density_reg32, density_reg33, density_reg34, density_reg35, density_reg36, density_reg37, density_reg38, density_reg39, density_reg40, density_reg41, density_reg42, density_reg43, density_reg44, density_reg45, density_reg46, density_reg47, density_reg48, density_reg49, density_reg50, density_reg51, density_reg52, density_reg53, density_reg54, density_reg55, density_reg56, density_reg57, density_reg58, density_reg59, density_reg60, density_reg61, density_reg62, density_reg63, density_reg64, density_reg65, density_reg66, density_reg67, density_reg68, density_reg69, density_reg70, density_reg71, density_reg72, density_reg73, density_reg74, density_reg75, density_reg76, density_reg77, density_reg78, density_reg79, density_reg80, density_reg81, density_reg82, density_reg83, density_reg84, density_reg85, density_reg86, density_reg87, density_reg88, density_reg89, density_reg90, density_reg91, density_reg92, density_reg93, density_reg94, density_reg95, density_reg96, density_reg97, density_reg98, density_reg99, density_reg100, density_reg101, density_reg102, density_reg103, density_reg104, density_reg105, density_reg106, density_reg107, density_reg108, density_reg109, density_reg110, density_reg111, density_reg112, density_reg113, density_reg114, density_reg115, density_reg116, density_reg117, density_reg118, density_reg119, density_reg120, density_reg121, density_reg122, density_reg123, density_reg124, density_reg125, density_reg126, density_reg127, density_reg128, density_reg129, density_reg130, density_reg131, density_reg132, density_reg133, density_reg134, density_reg135, density_reg136, density_reg137, density_reg138, density_reg139, density_reg140, density_reg141, density_reg142, density_reg143, density_reg144, density_reg145, density_reg146, density_reg147, density_reg148, density_reg149, density_reg150, density_reg151, density_reg152, density_reg153, density_reg154, density_reg155, density_reg156, density_reg157, density_reg158, density_reg159, density_reg160, density_reg161, density_reg162, density_reg163, density_reg164, density_reg165, density_reg166, density_reg167, density_reg168, density_reg169, density_reg170, density_reg171, density_reg172, density_reg173, density_reg174, density_reg175, density_reg176, density_reg177, density_reg178, density_reg179, density_reg180, density_reg181, density_reg182, density_reg183, density_reg184, density_reg185, density_reg186, density_reg187, density_reg188, density_reg189, density_reg190, density_reg191, density_reg192, density_reg193, density_reg194, density_reg195, density_reg196, density_reg197, density_reg198, density_reg199, density_reg200, density_reg201, density_reg202, density_reg203, density_reg204, density_reg205, density_reg206, density_reg207, density_reg208, density_reg209, density_reg210, density_reg211, density_reg212, density_reg213, density_reg214, density_reg215, density_reg216, density_reg217, density_reg218, density_reg219, density_reg220, density_reg221, density_reg222, density_reg223, density_reg224, density_reg225, density_reg226, density_reg227, density_reg228, density_reg229, density_reg230, density_reg231, density_reg232, density_reg233, density_reg234, density_reg235, density_reg236, density_reg237, density_reg238, density_reg239, density_reg240, density_reg241, density_reg242, density_reg243, density_reg244, density_reg245, density_reg246, density_reg247, density_reg248, density_reg249, density_reg250, density_reg251, density_reg252, density_reg253, density_reg254, density_reg255, density_reg256 }, { _2253_, _2252_, _2251_, _2250_, _2249_, _2248_, _2247_, _2246_, _2245_, _2244_, _2243_, _2242_, _2241_, _2240_, _2239_, _2238_, _2237_, _2236_, _2235_, _2234_, _2233_, _2232_, _2231_, _2230_, _2229_, _2228_, _2227_, _2226_, _2225_, _2224_, _2223_, _2222_, _2221_, _2220_, _2219_, _2218_, _2217_, _2216_, _2215_, _2214_, _2213_, _2212_, _2211_, _2210_, _2209_, _2208_, _2207_, _2206_, _2205_, _2204_, _2203_, _2202_, _2201_, _2200_, _2199_, _2198_, _2197_, _2196_, _2195_, _2194_, _2193_, _2192_, _2191_, _2190_, _2189_, _2188_, _2187_, _2186_, _2185_, _2184_, _2183_, _2182_, _2181_, _2180_, _2179_, _2178_, _2177_, _2176_, _2175_, _2174_, _2173_, _2172_, _2171_, _2170_, _2169_, _2168_, _2167_, _2166_, _2165_, _2164_, _2163_, _2162_, _2161_, _2160_, _2159_, _2158_, _2157_, _2156_, _2155_, _2154_, _2153_, _2152_, _2151_, _2150_, _2149_, _2148_, _2147_, _2146_, _2145_, _2144_, _2143_, _2142_, _2141_, _2140_, _2139_, _2138_, _2137_, _2136_, _2135_, _2134_, _2133_, _2132_, _2131_, _2130_, _2129_, _2128_, _2127_, _2126_, _2125_, _2124_, _2123_, _2122_, _2121_, _2120_, _2119_, _2118_, _2117_, _2116_, _2115_, _2114_, _2113_, _2112_, _2111_, _2110_, _2109_, _2108_, _2107_, _2106_, _2105_, _2104_, _2103_, _2102_, _2101_, _2100_, _2099_, _2098_, _2097_, _2096_, _2095_, _2094_, _2093_, _2092_, _2091_, _2090_, _2089_, _2088_, _2087_, _2086_, _2085_, _2084_, _2083_, _2082_, _2081_, _2080_, _2079_, _2078_, _2077_, _2076_, _2075_, _2074_, _2073_, _2072_, _2071_, _2070_, _2069_, _2068_, _2067_, _2066_, _2065_, _2064_, _2063_, _2062_, _2061_, _2060_, _2059_, _2058_, _2057_, _2056_, _2055_, _2054_, _2053_, _2052_, _2051_, _2050_, _2049_, _2048_, _2047_, _2046_, _2045_, _2044_, _2043_, _2042_, _2041_, _2040_, _2039_, _2038_, _2037_, _2036_, _2035_, _2034_, _2033_, _2032_, _2031_, _2030_, _2029_, _2028_, _2027_, _2026_, _2025_, _2024_, _2023_, _2022_, _2021_, _2020_, _2019_, _2018_, _2017_, _2016_, _2015_, _2014_, _2013_, _2012_, _2011_, _2010_, _2009_, _2008_, _2007_, _2006_, _2005_, _2004_, _2003_, _2002_, _2001_, _2000_, _1999_, _0404_ });
  assign _1997_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10350|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 9'b100000000;
  assign _1998_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10346|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 8'b11111111;
  assign _1999_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10342|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 8'b11111110;
  assign _2000_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10338|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 8'b11111101;
  assign _2001_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10334|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 8'b11111100;
  assign _2002_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10330|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 8'b11111011;
  assign _2003_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10326|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 8'b11111010;
  assign _2004_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10322|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 8'b11111001;
  assign _2005_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10318|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 8'b11111000;
  assign _2006_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10314|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 8'b11110111;
  assign _2007_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10310|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 8'b11110110;
  assign _2008_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10306|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 8'b11110101;
  assign _2009_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10302|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 8'b11110100;
  assign _2010_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10298|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 8'b11110011;
  assign _2011_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10294|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 8'b11110010;
  assign _2012_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10290|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 8'b11110001;
  assign _2013_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10286|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 8'b11110000;
  assign _2014_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10282|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 8'b11101111;
  assign _2015_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10278|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 8'b11101110;
  assign _2016_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10274|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 8'b11101101;
  assign _2017_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10270|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 8'b11101100;
  assign _2018_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10266|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 8'b11101011;
  assign _2019_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10262|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 8'b11101010;
  assign _2020_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10258|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 8'b11101001;
  assign _2021_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10254|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 8'b11101000;
  assign _2022_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10250|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 8'b11100111;
  assign _2023_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10246|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 8'b11100110;
  assign _2024_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10242|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 8'b11100101;
  assign _2025_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10238|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 8'b11100100;
  assign _2026_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10234|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 8'b11100011;
  assign _2027_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10230|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 8'b11100010;
  assign _2028_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10226|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 8'b11100001;
  assign _2029_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10222|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 8'b11100000;
  assign _2030_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10218|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 8'b11011111;
  assign _2031_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10214|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 8'b11011110;
  assign _2032_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10210|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 8'b11011101;
  assign _2033_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10206|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 8'b11011100;
  assign _2034_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10202|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 8'b11011011;
  assign _2035_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10198|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 8'b11011010;
  assign _2036_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10194|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 8'b11011001;
  assign _2037_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10190|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 8'b11011000;
  assign _2038_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10186|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 8'b11010111;
  assign _2039_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10182|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 8'b11010110;
  assign _2040_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10178|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 8'b11010101;
  assign _2041_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10174|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 8'b11010100;
  assign _2042_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10170|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 8'b11010011;
  assign _2043_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10166|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 8'b11010010;
  assign _2044_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10162|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 8'b11010001;
  assign _2045_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10158|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 8'b11010000;
  assign _2046_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10154|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 8'b11001111;
  assign _2047_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10150|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 8'b11001110;
  assign _2048_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10146|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 8'b11001101;
  assign _2049_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10142|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 8'b11001100;
  assign _2050_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10138|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 8'b11001011;
  assign _2051_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10134|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 8'b11001010;
  assign _2052_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10130|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 8'b11001001;
  assign _2053_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10126|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 8'b11001000;
  assign _2054_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10122|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 8'b11000111;
  assign _2055_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10118|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 8'b11000110;
  assign _2056_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10114|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 8'b11000101;
  assign _2057_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10110|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 8'b11000100;
  assign _2058_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10106|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 8'b11000011;
  assign _2059_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10102|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 8'b11000010;
  assign _2060_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10098|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 8'b11000001;
  assign _2061_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10094|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 8'b11000000;
  assign _2062_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10090|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 8'b10111111;
  assign _2063_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10086|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 8'b10111110;
  assign _2064_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10082|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 8'b10111101;
  assign _2065_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10078|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 8'b10111100;
  assign _2066_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10074|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 8'b10111011;
  assign _2067_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10070|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 8'b10111010;
  assign _2068_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10066|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 8'b10111001;
  assign _2069_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10062|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 8'b10111000;
  assign _2070_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10058|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 8'b10110111;
  assign _2071_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10054|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 8'b10110110;
  assign _2072_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10050|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 8'b10110101;
  assign _2073_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10046|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 8'b10110100;
  assign _2074_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10042|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 8'b10110011;
  assign _2075_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10038|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 8'b10110010;
  assign _2076_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10034|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 8'b10110001;
  assign _2077_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10030|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 8'b10110000;
  assign _2078_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10026|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 8'b10101111;
  assign _2079_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10022|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 8'b10101110;
  assign _2080_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10018|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 8'b10101101;
  assign _2081_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10014|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 8'b10101100;
  assign _2082_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10010|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 8'b10101011;
  assign _2083_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10006|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 8'b10101010;
  assign _2084_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10002|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 8'b10101001;
  assign _2085_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9998|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 8'b10101000;
  assign _2086_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9994|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 8'b10100111;
  assign _2087_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9990|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 8'b10100110;
  assign _2088_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9986|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 8'b10100101;
  assign _2089_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9982|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 8'b10100100;
  assign _2090_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9978|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 8'b10100011;
  assign _2091_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9974|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 8'b10100010;
  assign _2092_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9970|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 8'b10100001;
  assign _2093_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9966|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 8'b10100000;
  assign _2094_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9962|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 8'b10011111;
  assign _2095_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9958|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 8'b10011110;
  assign _2096_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9954|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 8'b10011101;
  assign _2097_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9950|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 8'b10011100;
  assign _2098_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9946|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 8'b10011011;
  assign _2099_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9942|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 8'b10011010;
  assign _2100_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9938|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 8'b10011001;
  assign _2101_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9934|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 8'b10011000;
  assign _2102_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9930|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 8'b10010111;
  assign _2103_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9926|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 8'b10010110;
  assign _2104_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9922|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 8'b10010101;
  assign _2105_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9918|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 8'b10010100;
  assign _2106_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9914|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 8'b10010011;
  assign _2107_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9910|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 8'b10010010;
  assign _2108_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9906|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 8'b10010001;
  assign _2109_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9902|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 8'b10010000;
  assign _2110_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9898|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 8'b10001111;
  assign _2111_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9894|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 8'b10001110;
  assign _2112_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9890|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 8'b10001101;
  assign _2113_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9886|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 8'b10001100;
  assign _2114_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9882|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 8'b10001011;
  assign _2115_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9878|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 8'b10001010;
  assign _2116_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9874|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 8'b10001001;
  assign _2117_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9870|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 8'b10001000;
  assign _2118_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9866|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 8'b10000111;
  assign _2119_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9862|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 8'b10000110;
  assign _2120_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9858|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 8'b10000101;
  assign _2121_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9854|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 8'b10000100;
  assign _2122_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9850|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 8'b10000011;
  assign _2123_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9846|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 8'b10000010;
  assign _2124_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9842|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 8'b10000001;
  assign _2125_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9838|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 8'b10000000;
  assign _2126_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9834|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 7'b1111111;
  assign _2127_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9830|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 7'b1111110;
  assign _2128_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9826|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 7'b1111101;
  assign _2129_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9822|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 7'b1111100;
  assign _2130_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9818|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 7'b1111011;
  assign _2131_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9814|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 7'b1111010;
  assign _2132_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9810|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 7'b1111001;
  assign _2133_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9806|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 7'b1111000;
  assign _2134_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9802|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 7'b1110111;
  assign _2135_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9798|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 7'b1110110;
  assign _2136_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9794|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 7'b1110101;
  assign _2137_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9790|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 7'b1110100;
  assign _2138_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9786|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 7'b1110011;
  assign _2139_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9782|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 7'b1110010;
  assign _2140_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9778|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 7'b1110001;
  assign _2141_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9774|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 7'b1110000;
  assign _2142_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9770|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 7'b1101111;
  assign _2143_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9766|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 7'b1101110;
  assign _2144_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9762|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 7'b1101101;
  assign _2145_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9758|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 7'b1101100;
  assign _2146_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9754|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 7'b1101011;
  assign _2147_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9750|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 7'b1101010;
  assign _2148_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9746|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 7'b1101001;
  assign _2149_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9742|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 7'b1101000;
  assign _2150_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9738|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 7'b1100111;
  assign _2151_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9734|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 7'b1100110;
  assign _2152_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9730|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 7'b1100101;
  assign _2153_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9726|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 7'b1100100;
  assign _2154_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9722|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 7'b1100011;
  assign _2155_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9718|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 7'b1100010;
  assign _2156_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9714|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 7'b1100001;
  assign _2157_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9710|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 7'b1100000;
  assign _2158_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9706|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 7'b1011111;
  assign _2159_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9702|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 7'b1011110;
  assign _2160_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9698|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 7'b1011101;
  assign _2161_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9694|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 7'b1011100;
  assign _2162_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9690|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 7'b1011011;
  assign _2163_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9686|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 7'b1011010;
  assign _2164_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9682|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 7'b1011001;
  assign _2165_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9678|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 7'b1011000;
  assign _2166_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9674|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 7'b1010111;
  assign _2167_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9670|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 7'b1010110;
  assign _2168_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9666|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 7'b1010101;
  assign _2169_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9662|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 7'b1010100;
  assign _2170_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9658|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 7'b1010011;
  assign _2171_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9654|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 7'b1010010;
  assign _2172_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9650|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 7'b1010001;
  assign _2173_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9646|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 7'b1010000;
  assign _2174_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9642|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 7'b1001111;
  assign _2175_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9638|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 7'b1001110;
  assign _2176_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9634|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 7'b1001101;
  assign _2177_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9630|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 7'b1001100;
  assign _2178_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9626|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 7'b1001011;
  assign _2179_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9622|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 7'b1001010;
  assign _2180_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9618|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 7'b1001001;
  assign _2181_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9614|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 7'b1001000;
  assign _2182_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9610|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 7'b1000111;
  assign _2183_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9606|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 7'b1000110;
  assign _2184_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9602|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 7'b1000101;
  assign _2185_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9598|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 7'b1000100;
  assign _2186_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9594|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 7'b1000011;
  assign _2187_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9590|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 7'b1000010;
  assign _2188_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9586|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 7'b1000001;
  assign _2189_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9582|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 7'b1000000;
  assign _2190_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9578|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 6'b111111;
  assign _2191_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9574|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 6'b111110;
  assign _2192_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9570|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 6'b111101;
  assign _2193_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9566|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 6'b111100;
  assign _2194_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9562|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 6'b111011;
  assign _2195_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9558|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 6'b111010;
  assign _2196_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9554|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 6'b111001;
  assign _2197_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9550|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 6'b111000;
  assign _2198_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9546|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 6'b110111;
  assign _2199_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9542|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 6'b110110;
  assign _2200_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9538|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 6'b110101;
  assign _2201_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9534|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 6'b110100;
  assign _2202_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9530|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 6'b110011;
  assign _2203_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9526|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 6'b110010;
  assign _2204_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9522|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 6'b110001;
  assign _2205_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9518|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 6'b110000;
  assign _2206_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9514|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 6'b101111;
  assign _2207_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9510|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 6'b101110;
  assign _2208_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9506|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 6'b101101;
  assign _2209_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9502|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 6'b101100;
  assign _2210_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9498|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 6'b101011;
  assign _2211_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9494|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 6'b101010;
  assign _2212_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9490|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 6'b101001;
  assign _2213_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9486|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 6'b101000;
  assign _2214_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9482|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 6'b100111;
  assign _2215_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9478|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 6'b100110;
  assign _2216_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9474|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 6'b100101;
  assign _2217_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9470|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 6'b100100;
  assign _2218_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9466|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 6'b100011;
  assign _2219_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9462|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 6'b100010;
  assign _2220_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9458|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 6'b100001;
  assign _2221_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9454|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 6'b100000;
  assign _2222_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9450|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 5'b11111;
  assign _2223_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9446|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 5'b11110;
  assign _2224_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9442|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 5'b11101;
  assign _2225_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9438|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 5'b11100;
  assign _2226_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9434|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 5'b11011;
  assign _2227_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9430|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 5'b11010;
  assign _2228_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9426|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 5'b11001;
  assign _2229_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9422|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 5'b11000;
  assign _2230_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9418|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 5'b10111;
  assign _2231_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9414|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 5'b10110;
  assign _2232_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9410|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 5'b10101;
  assign _2233_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9406|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 5'b10100;
  assign _2234_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9402|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 5'b10011;
  assign _2235_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9398|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 5'b10010;
  assign _2236_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9394|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 5'b10001;
  assign _2237_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9390|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 5'b10000;
  assign _2238_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9386|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 4'b1111;
  assign _2239_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9382|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 4'b1110;
  assign _2240_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9378|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 4'b1101;
  assign _2241_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9374|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 4'b1100;
  assign _2242_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9370|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 4'b1011;
  assign _2243_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9366|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 4'b1010;
  assign _2244_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9362|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 4'b1001;
  assign _2245_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9358|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 4'b1000;
  assign _2246_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9354|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 3'b111;
  assign _2247_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9350|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 3'b110;
  assign _2248_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9346|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 3'b101;
  assign _2249_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9342|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 3'b100;
  assign _2250_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9338|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 2'b11;
  assign _2251_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9334|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 2'b10;
  assign _2252_ = dp2lut_Y_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9330|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) 1'b1;
  assign _2253_ = ! (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9326|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *) dp2lut_Y_entry_2;
  assign _2254_ = dp2lut_Yinfo_2[17] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9321" *) density_reg256 : _1996_;
  assign _2255_ = dp2lut_Yinfo_2[16] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9318" *) density_reg0 : _2254_;
  assign _0290_ = _0402_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9317" *) _2255_ : lut_Y_data_21;
  function [15:0] _6110_;
    input [15:0] a;
    input [4095:0] b;
    input [255:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:10350|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9325" *)
    (* parallel_case *)
    casez (s)
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1:
        _6110_ = b[15:0];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?:
        _6110_ = b[31:16];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??:
        _6110_ = b[47:32];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???:
        _6110_ = b[63:48];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????:
        _6110_ = b[79:64];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????:
        _6110_ = b[95:80];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????:
        _6110_ = b[111:96];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????:
        _6110_ = b[127:112];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????:
        _6110_ = b[143:128];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????:
        _6110_ = b[159:144];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????:
        _6110_ = b[175:160];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????:
        _6110_ = b[191:176];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????:
        _6110_ = b[207:192];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????:
        _6110_ = b[223:208];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????:
        _6110_ = b[239:224];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????:
        _6110_ = b[255:240];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????:
        _6110_ = b[271:256];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????:
        _6110_ = b[287:272];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????:
        _6110_ = b[303:288];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????:
        _6110_ = b[319:304];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????:
        _6110_ = b[335:320];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????:
        _6110_ = b[351:336];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????:
        _6110_ = b[367:352];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????:
        _6110_ = b[383:368];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????:
        _6110_ = b[399:384];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????:
        _6110_ = b[415:400];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????:
        _6110_ = b[431:416];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????:
        _6110_ = b[447:432];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????:
        _6110_ = b[463:448];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????:
        _6110_ = b[479:464];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????:
        _6110_ = b[495:480];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????:
        _6110_ = b[511:496];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????:
        _6110_ = b[527:512];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????:
        _6110_ = b[543:528];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????:
        _6110_ = b[559:544];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????:
        _6110_ = b[575:560];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????:
        _6110_ = b[591:576];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????:
        _6110_ = b[607:592];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????:
        _6110_ = b[623:608];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????:
        _6110_ = b[639:624];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????:
        _6110_ = b[655:640];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????:
        _6110_ = b[671:656];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????:
        _6110_ = b[687:672];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????:
        _6110_ = b[703:688];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????:
        _6110_ = b[719:704];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????:
        _6110_ = b[735:720];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????:
        _6110_ = b[751:736];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????:
        _6110_ = b[767:752];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????:
        _6110_ = b[783:768];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????:
        _6110_ = b[799:784];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????:
        _6110_ = b[815:800];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????:
        _6110_ = b[831:816];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????:
        _6110_ = b[847:832];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????:
        _6110_ = b[863:848];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????:
        _6110_ = b[879:864];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????:
        _6110_ = b[895:880];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????:
        _6110_ = b[911:896];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????:
        _6110_ = b[927:912];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????:
        _6110_ = b[943:928];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????:
        _6110_ = b[959:944];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????:
        _6110_ = b[975:960];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????:
        _6110_ = b[991:976];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????:
        _6110_ = b[1007:992];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????:
        _6110_ = b[1023:1008];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????:
        _6110_ = b[1039:1024];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????:
        _6110_ = b[1055:1040];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????:
        _6110_ = b[1071:1056];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????:
        _6110_ = b[1087:1072];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????:
        _6110_ = b[1103:1088];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????:
        _6110_ = b[1119:1104];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????:
        _6110_ = b[1135:1120];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????:
        _6110_ = b[1151:1136];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????:
        _6110_ = b[1167:1152];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????:
        _6110_ = b[1183:1168];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????:
        _6110_ = b[1199:1184];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????:
        _6110_ = b[1215:1200];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????:
        _6110_ = b[1231:1216];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????:
        _6110_ = b[1247:1232];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????:
        _6110_ = b[1263:1248];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????:
        _6110_ = b[1279:1264];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????:
        _6110_ = b[1295:1280];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????:
        _6110_ = b[1311:1296];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????:
        _6110_ = b[1327:1312];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????:
        _6110_ = b[1343:1328];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????:
        _6110_ = b[1359:1344];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????:
        _6110_ = b[1375:1360];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????:
        _6110_ = b[1391:1376];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????:
        _6110_ = b[1407:1392];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????:
        _6110_ = b[1423:1408];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????:
        _6110_ = b[1439:1424];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????:
        _6110_ = b[1455:1440];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????:
        _6110_ = b[1471:1456];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????:
        _6110_ = b[1487:1472];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????:
        _6110_ = b[1503:1488];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????:
        _6110_ = b[1519:1504];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????:
        _6110_ = b[1535:1520];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????:
        _6110_ = b[1551:1536];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????:
        _6110_ = b[1567:1552];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????:
        _6110_ = b[1583:1568];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????:
        _6110_ = b[1599:1584];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6110_ = b[1615:1600];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6110_ = b[1631:1616];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6110_ = b[1647:1632];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6110_ = b[1663:1648];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6110_ = b[1679:1664];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6110_ = b[1695:1680];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6110_ = b[1711:1696];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6110_ = b[1727:1712];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6110_ = b[1743:1728];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6110_ = b[1759:1744];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6110_ = b[1775:1760];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6110_ = b[1791:1776];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6110_ = b[1807:1792];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6110_ = b[1823:1808];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6110_ = b[1839:1824];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6110_ = b[1855:1840];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6110_ = b[1871:1856];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6110_ = b[1887:1872];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6110_ = b[1903:1888];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6110_ = b[1919:1904];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6110_ = b[1935:1920];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6110_ = b[1951:1936];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6110_ = b[1967:1952];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6110_ = b[1983:1968];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6110_ = b[1999:1984];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6110_ = b[2015:2000];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6110_ = b[2031:2016];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6110_ = b[2047:2032];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6110_ = b[2063:2048];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6110_ = b[2079:2064];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6110_ = b[2095:2080];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6110_ = b[2111:2096];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6110_ = b[2127:2112];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6110_ = b[2143:2128];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6110_ = b[2159:2144];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6110_ = b[2175:2160];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6110_ = b[2191:2176];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6110_ = b[2207:2192];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6110_ = b[2223:2208];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6110_ = b[2239:2224];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6110_ = b[2255:2240];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6110_ = b[2271:2256];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6110_ = b[2287:2272];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6110_ = b[2303:2288];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6110_ = b[2319:2304];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6110_ = b[2335:2320];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6110_ = b[2351:2336];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6110_ = b[2367:2352];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6110_ = b[2383:2368];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6110_ = b[2399:2384];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6110_ = b[2415:2400];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6110_ = b[2431:2416];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6110_ = b[2447:2432];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6110_ = b[2463:2448];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6110_ = b[2479:2464];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6110_ = b[2495:2480];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6110_ = b[2511:2496];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6110_ = b[2527:2512];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6110_ = b[2543:2528];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6110_ = b[2559:2544];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6110_ = b[2575:2560];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6110_ = b[2591:2576];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6110_ = b[2607:2592];
      256'b????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6110_ = b[2623:2608];
      256'b???????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6110_ = b[2639:2624];
      256'b??????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6110_ = b[2655:2640];
      256'b?????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6110_ = b[2671:2656];
      256'b????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6110_ = b[2687:2672];
      256'b???????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6110_ = b[2703:2688];
      256'b??????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6110_ = b[2719:2704];
      256'b?????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6110_ = b[2735:2720];
      256'b????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6110_ = b[2751:2736];
      256'b???????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6110_ = b[2767:2752];
      256'b??????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6110_ = b[2783:2768];
      256'b?????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6110_ = b[2799:2784];
      256'b????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6110_ = b[2815:2800];
      256'b???????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6110_ = b[2831:2816];
      256'b??????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6110_ = b[2847:2832];
      256'b?????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6110_ = b[2863:2848];
      256'b????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6110_ = b[2879:2864];
      256'b???????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6110_ = b[2895:2880];
      256'b??????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6110_ = b[2911:2896];
      256'b?????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6110_ = b[2927:2912];
      256'b????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6110_ = b[2943:2928];
      256'b???????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6110_ = b[2959:2944];
      256'b??????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6110_ = b[2975:2960];
      256'b?????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6110_ = b[2991:2976];
      256'b????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6110_ = b[3007:2992];
      256'b???????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6110_ = b[3023:3008];
      256'b??????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6110_ = b[3039:3024];
      256'b?????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6110_ = b[3055:3040];
      256'b????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6110_ = b[3071:3056];
      256'b???????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6110_ = b[3087:3072];
      256'b??????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6110_ = b[3103:3088];
      256'b?????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6110_ = b[3119:3104];
      256'b????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6110_ = b[3135:3120];
      256'b???????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6110_ = b[3151:3136];
      256'b??????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6110_ = b[3167:3152];
      256'b?????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6110_ = b[3183:3168];
      256'b????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6110_ = b[3199:3184];
      256'b???????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6110_ = b[3215:3200];
      256'b??????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6110_ = b[3231:3216];
      256'b?????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6110_ = b[3247:3232];
      256'b????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6110_ = b[3263:3248];
      256'b???????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6110_ = b[3279:3264];
      256'b??????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6110_ = b[3295:3280];
      256'b?????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6110_ = b[3311:3296];
      256'b????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6110_ = b[3327:3312];
      256'b???????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6110_ = b[3343:3328];
      256'b??????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6110_ = b[3359:3344];
      256'b?????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6110_ = b[3375:3360];
      256'b????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6110_ = b[3391:3376];
      256'b???????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6110_ = b[3407:3392];
      256'b??????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6110_ = b[3423:3408];
      256'b?????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6110_ = b[3439:3424];
      256'b????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6110_ = b[3455:3440];
      256'b???????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6110_ = b[3471:3456];
      256'b??????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6110_ = b[3487:3472];
      256'b?????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6110_ = b[3503:3488];
      256'b????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6110_ = b[3519:3504];
      256'b???????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6110_ = b[3535:3520];
      256'b??????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6110_ = b[3551:3536];
      256'b?????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6110_ = b[3567:3552];
      256'b????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6110_ = b[3583:3568];
      256'b???????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6110_ = b[3599:3584];
      256'b??????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6110_ = b[3615:3600];
      256'b?????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6110_ = b[3631:3616];
      256'b????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6110_ = b[3647:3632];
      256'b???????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6110_ = b[3663:3648];
      256'b??????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6110_ = b[3679:3664];
      256'b?????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6110_ = b[3695:3680];
      256'b????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6110_ = b[3711:3696];
      256'b???????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6110_ = b[3727:3712];
      256'b??????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6110_ = b[3743:3728];
      256'b?????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6110_ = b[3759:3744];
      256'b????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6110_ = b[3775:3760];
      256'b???????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6110_ = b[3791:3776];
      256'b??????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6110_ = b[3807:3792];
      256'b?????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6110_ = b[3823:3808];
      256'b????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6110_ = b[3839:3824];
      256'b???????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6110_ = b[3855:3840];
      256'b??????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6110_ = b[3871:3856];
      256'b?????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6110_ = b[3887:3872];
      256'b????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6110_ = b[3903:3888];
      256'b???????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6110_ = b[3919:3904];
      256'b??????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6110_ = b[3935:3920];
      256'b?????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6110_ = b[3951:3936];
      256'b????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6110_ = b[3967:3952];
      256'b???????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6110_ = b[3983:3968];
      256'b??????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6110_ = b[3999:3984];
      256'b?????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6110_ = b[4015:4000];
      256'b????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6110_ = b[4031:4016];
      256'b???1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6110_ = b[4047:4032];
      256'b??1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6110_ = b[4063:4048];
      256'b?1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6110_ = b[4079:4064];
      256'b1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6110_ = b[4095:4080];
      default:
        _6110_ = a;
    endcase
  endfunction
  assign _2256_ = _6110_(density_reg0, { density_reg1, density_reg2, density_reg3, density_reg4, density_reg5, density_reg6, density_reg7, density_reg8, density_reg9, density_reg10, density_reg11, density_reg12, density_reg13, density_reg14, density_reg15, density_reg16, density_reg17, density_reg18, density_reg19, density_reg20, density_reg21, density_reg22, density_reg23, density_reg24, density_reg25, density_reg26, density_reg27, density_reg28, density_reg29, density_reg30, density_reg31, density_reg32, density_reg33, density_reg34, density_reg35, density_reg36, density_reg37, density_reg38, density_reg39, density_reg40, density_reg41, density_reg42, density_reg43, density_reg44, density_reg45, density_reg46, density_reg47, density_reg48, density_reg49, density_reg50, density_reg51, density_reg52, density_reg53, density_reg54, density_reg55, density_reg56, density_reg57, density_reg58, density_reg59, density_reg60, density_reg61, density_reg62, density_reg63, density_reg64, density_reg65, density_reg66, density_reg67, density_reg68, density_reg69, density_reg70, density_reg71, density_reg72, density_reg73, density_reg74, density_reg75, density_reg76, density_reg77, density_reg78, density_reg79, density_reg80, density_reg81, density_reg82, density_reg83, density_reg84, density_reg85, density_reg86, density_reg87, density_reg88, density_reg89, density_reg90, density_reg91, density_reg92, density_reg93, density_reg94, density_reg95, density_reg96, density_reg97, density_reg98, density_reg99, density_reg100, density_reg101, density_reg102, density_reg103, density_reg104, density_reg105, density_reg106, density_reg107, density_reg108, density_reg109, density_reg110, density_reg111, density_reg112, density_reg113, density_reg114, density_reg115, density_reg116, density_reg117, density_reg118, density_reg119, density_reg120, density_reg121, density_reg122, density_reg123, density_reg124, density_reg125, density_reg126, density_reg127, density_reg128, density_reg129, density_reg130, density_reg131, density_reg132, density_reg133, density_reg134, density_reg135, density_reg136, density_reg137, density_reg138, density_reg139, density_reg140, density_reg141, density_reg142, density_reg143, density_reg144, density_reg145, density_reg146, density_reg147, density_reg148, density_reg149, density_reg150, density_reg151, density_reg152, density_reg153, density_reg154, density_reg155, density_reg156, density_reg157, density_reg158, density_reg159, density_reg160, density_reg161, density_reg162, density_reg163, density_reg164, density_reg165, density_reg166, density_reg167, density_reg168, density_reg169, density_reg170, density_reg171, density_reg172, density_reg173, density_reg174, density_reg175, density_reg176, density_reg177, density_reg178, density_reg179, density_reg180, density_reg181, density_reg182, density_reg183, density_reg184, density_reg185, density_reg186, density_reg187, density_reg188, density_reg189, density_reg190, density_reg191, density_reg192, density_reg193, density_reg194, density_reg195, density_reg196, density_reg197, density_reg198, density_reg199, density_reg200, density_reg201, density_reg202, density_reg203, density_reg204, density_reg205, density_reg206, density_reg207, density_reg208, density_reg209, density_reg210, density_reg211, density_reg212, density_reg213, density_reg214, density_reg215, density_reg216, density_reg217, density_reg218, density_reg219, density_reg220, density_reg221, density_reg222, density_reg223, density_reg224, density_reg225, density_reg226, density_reg227, density_reg228, density_reg229, density_reg230, density_reg231, density_reg232, density_reg233, density_reg234, density_reg235, density_reg236, density_reg237, density_reg238, density_reg239, density_reg240, density_reg241, density_reg242, density_reg243, density_reg244, density_reg245, density_reg246, density_reg247, density_reg248, density_reg249, density_reg250, density_reg251, density_reg252, density_reg253, density_reg254, density_reg255, density_reg256 }, { _2252_, _2251_, _2250_, _2249_, _2248_, _2247_, _2246_, _2245_, _2244_, _2243_, _2242_, _2241_, _2240_, _2239_, _2238_, _2237_, _2236_, _2235_, _2234_, _2233_, _2232_, _2231_, _2230_, _2229_, _2228_, _2227_, _2226_, _2225_, _2224_, _2223_, _2222_, _2221_, _2220_, _2219_, _2218_, _2217_, _2216_, _2215_, _2214_, _2213_, _2212_, _2211_, _2210_, _2209_, _2208_, _2207_, _2206_, _2205_, _2204_, _2203_, _2202_, _2201_, _2200_, _2199_, _2198_, _2197_, _2196_, _2195_, _2194_, _2193_, _2192_, _2191_, _2190_, _2189_, _2188_, _2187_, _2186_, _2185_, _2184_, _2183_, _2182_, _2181_, _2180_, _2179_, _2178_, _2177_, _2176_, _2175_, _2174_, _2173_, _2172_, _2171_, _2170_, _2169_, _2168_, _2167_, _2166_, _2165_, _2164_, _2163_, _2162_, _2161_, _2160_, _2159_, _2158_, _2157_, _2156_, _2155_, _2154_, _2153_, _2152_, _2151_, _2150_, _2149_, _2148_, _2147_, _2146_, _2145_, _2144_, _2143_, _2142_, _2141_, _2140_, _2139_, _2138_, _2137_, _2136_, _2135_, _2134_, _2133_, _2132_, _2131_, _2130_, _2129_, _2128_, _2127_, _2126_, _2125_, _2124_, _2123_, _2122_, _2121_, _2120_, _2119_, _2118_, _2117_, _2116_, _2115_, _2114_, _2113_, _2112_, _2111_, _2110_, _2109_, _2108_, _2107_, _2106_, _2105_, _2104_, _2103_, _2102_, _2101_, _2100_, _2099_, _2098_, _2097_, _2096_, _2095_, _2094_, _2093_, _2092_, _2091_, _2090_, _2089_, _2088_, _2087_, _2086_, _2085_, _2084_, _2083_, _2082_, _2081_, _2080_, _2079_, _2078_, _2077_, _2076_, _2075_, _2074_, _2073_, _2072_, _2071_, _2070_, _2069_, _2068_, _2067_, _2066_, _2065_, _2064_, _2063_, _2062_, _2061_, _2060_, _2059_, _2058_, _2057_, _2056_, _2055_, _2054_, _2053_, _2052_, _2051_, _2050_, _2049_, _2048_, _2047_, _2046_, _2045_, _2044_, _2043_, _2042_, _2041_, _2040_, _2039_, _2038_, _2037_, _2036_, _2035_, _2034_, _2033_, _2032_, _2031_, _2030_, _2029_, _2028_, _2027_, _2026_, _2025_, _2024_, _2023_, _2022_, _2021_, _2020_, _2019_, _2018_, _2017_, _2016_, _2015_, _2014_, _2013_, _2012_, _2011_, _2010_, _2009_, _2008_, _2007_, _2006_, _2005_, _2004_, _2003_, _2002_, _2001_, _2000_, _1999_, _1998_, _1997_ });
  assign _2257_ = dp2lut_Yinfo_2[17] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9321" *) density_reg256 : _2256_;
  assign _2258_ = dp2lut_Yinfo_2[16] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9318" *) density_reg0 : _2257_;
  assign _0289_ = _0402_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9317" *) _2258_ : lut_Y_data_20;
  function [15:0] _6114_;
    input [15:0] a;
    input [4095:0] b;
    input [255:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9299|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *)
    (* parallel_case *)
    casez (s)
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1:
        _6114_ = b[15:0];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?:
        _6114_ = b[31:16];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??:
        _6114_ = b[47:32];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???:
        _6114_ = b[63:48];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????:
        _6114_ = b[79:64];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????:
        _6114_ = b[95:80];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????:
        _6114_ = b[111:96];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????:
        _6114_ = b[127:112];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????:
        _6114_ = b[143:128];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????:
        _6114_ = b[159:144];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????:
        _6114_ = b[175:160];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????:
        _6114_ = b[191:176];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????:
        _6114_ = b[207:192];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????:
        _6114_ = b[223:208];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????:
        _6114_ = b[239:224];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????:
        _6114_ = b[255:240];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????:
        _6114_ = b[271:256];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????:
        _6114_ = b[287:272];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????:
        _6114_ = b[303:288];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????:
        _6114_ = b[319:304];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????:
        _6114_ = b[335:320];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????:
        _6114_ = b[351:336];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????:
        _6114_ = b[367:352];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????:
        _6114_ = b[383:368];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????:
        _6114_ = b[399:384];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????:
        _6114_ = b[415:400];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????:
        _6114_ = b[431:416];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????:
        _6114_ = b[447:432];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????:
        _6114_ = b[463:448];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????:
        _6114_ = b[479:464];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????:
        _6114_ = b[495:480];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????:
        _6114_ = b[511:496];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????:
        _6114_ = b[527:512];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????:
        _6114_ = b[543:528];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????:
        _6114_ = b[559:544];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????:
        _6114_ = b[575:560];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????:
        _6114_ = b[591:576];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????:
        _6114_ = b[607:592];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????:
        _6114_ = b[623:608];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????:
        _6114_ = b[639:624];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????:
        _6114_ = b[655:640];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????:
        _6114_ = b[671:656];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????:
        _6114_ = b[687:672];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????:
        _6114_ = b[703:688];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????:
        _6114_ = b[719:704];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????:
        _6114_ = b[735:720];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????:
        _6114_ = b[751:736];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????:
        _6114_ = b[767:752];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????:
        _6114_ = b[783:768];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????:
        _6114_ = b[799:784];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????:
        _6114_ = b[815:800];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????:
        _6114_ = b[831:816];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????:
        _6114_ = b[847:832];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????:
        _6114_ = b[863:848];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????:
        _6114_ = b[879:864];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????:
        _6114_ = b[895:880];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????:
        _6114_ = b[911:896];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????:
        _6114_ = b[927:912];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????:
        _6114_ = b[943:928];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????:
        _6114_ = b[959:944];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????:
        _6114_ = b[975:960];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????:
        _6114_ = b[991:976];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????:
        _6114_ = b[1007:992];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????:
        _6114_ = b[1023:1008];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????:
        _6114_ = b[1039:1024];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????:
        _6114_ = b[1055:1040];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????:
        _6114_ = b[1071:1056];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????:
        _6114_ = b[1087:1072];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????:
        _6114_ = b[1103:1088];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????:
        _6114_ = b[1119:1104];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????:
        _6114_ = b[1135:1120];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????:
        _6114_ = b[1151:1136];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????:
        _6114_ = b[1167:1152];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????:
        _6114_ = b[1183:1168];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????:
        _6114_ = b[1199:1184];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????:
        _6114_ = b[1215:1200];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????:
        _6114_ = b[1231:1216];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????:
        _6114_ = b[1247:1232];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????:
        _6114_ = b[1263:1248];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????:
        _6114_ = b[1279:1264];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????:
        _6114_ = b[1295:1280];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????:
        _6114_ = b[1311:1296];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????:
        _6114_ = b[1327:1312];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????:
        _6114_ = b[1343:1328];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????:
        _6114_ = b[1359:1344];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????:
        _6114_ = b[1375:1360];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????:
        _6114_ = b[1391:1376];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????:
        _6114_ = b[1407:1392];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????:
        _6114_ = b[1423:1408];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????:
        _6114_ = b[1439:1424];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????:
        _6114_ = b[1455:1440];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????:
        _6114_ = b[1471:1456];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????:
        _6114_ = b[1487:1472];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????:
        _6114_ = b[1503:1488];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????:
        _6114_ = b[1519:1504];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????:
        _6114_ = b[1535:1520];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????:
        _6114_ = b[1551:1536];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????:
        _6114_ = b[1567:1552];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????:
        _6114_ = b[1583:1568];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????:
        _6114_ = b[1599:1584];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6114_ = b[1615:1600];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6114_ = b[1631:1616];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6114_ = b[1647:1632];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6114_ = b[1663:1648];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6114_ = b[1679:1664];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6114_ = b[1695:1680];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6114_ = b[1711:1696];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6114_ = b[1727:1712];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6114_ = b[1743:1728];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6114_ = b[1759:1744];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6114_ = b[1775:1760];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6114_ = b[1791:1776];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6114_ = b[1807:1792];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6114_ = b[1823:1808];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6114_ = b[1839:1824];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6114_ = b[1855:1840];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6114_ = b[1871:1856];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6114_ = b[1887:1872];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6114_ = b[1903:1888];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6114_ = b[1919:1904];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6114_ = b[1935:1920];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6114_ = b[1951:1936];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6114_ = b[1967:1952];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6114_ = b[1983:1968];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6114_ = b[1999:1984];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6114_ = b[2015:2000];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6114_ = b[2031:2016];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6114_ = b[2047:2032];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6114_ = b[2063:2048];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6114_ = b[2079:2064];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6114_ = b[2095:2080];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6114_ = b[2111:2096];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6114_ = b[2127:2112];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6114_ = b[2143:2128];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6114_ = b[2159:2144];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6114_ = b[2175:2160];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6114_ = b[2191:2176];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6114_ = b[2207:2192];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6114_ = b[2223:2208];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6114_ = b[2239:2224];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6114_ = b[2255:2240];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6114_ = b[2271:2256];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6114_ = b[2287:2272];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6114_ = b[2303:2288];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6114_ = b[2319:2304];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6114_ = b[2335:2320];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6114_ = b[2351:2336];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6114_ = b[2367:2352];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6114_ = b[2383:2368];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6114_ = b[2399:2384];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6114_ = b[2415:2400];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6114_ = b[2431:2416];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6114_ = b[2447:2432];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6114_ = b[2463:2448];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6114_ = b[2479:2464];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6114_ = b[2495:2480];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6114_ = b[2511:2496];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6114_ = b[2527:2512];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6114_ = b[2543:2528];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6114_ = b[2559:2544];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6114_ = b[2575:2560];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6114_ = b[2591:2576];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6114_ = b[2607:2592];
      256'b????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6114_ = b[2623:2608];
      256'b???????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6114_ = b[2639:2624];
      256'b??????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6114_ = b[2655:2640];
      256'b?????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6114_ = b[2671:2656];
      256'b????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6114_ = b[2687:2672];
      256'b???????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6114_ = b[2703:2688];
      256'b??????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6114_ = b[2719:2704];
      256'b?????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6114_ = b[2735:2720];
      256'b????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6114_ = b[2751:2736];
      256'b???????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6114_ = b[2767:2752];
      256'b??????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6114_ = b[2783:2768];
      256'b?????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6114_ = b[2799:2784];
      256'b????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6114_ = b[2815:2800];
      256'b???????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6114_ = b[2831:2816];
      256'b??????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6114_ = b[2847:2832];
      256'b?????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6114_ = b[2863:2848];
      256'b????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6114_ = b[2879:2864];
      256'b???????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6114_ = b[2895:2880];
      256'b??????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6114_ = b[2911:2896];
      256'b?????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6114_ = b[2927:2912];
      256'b????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6114_ = b[2943:2928];
      256'b???????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6114_ = b[2959:2944];
      256'b??????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6114_ = b[2975:2960];
      256'b?????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6114_ = b[2991:2976];
      256'b????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6114_ = b[3007:2992];
      256'b???????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6114_ = b[3023:3008];
      256'b??????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6114_ = b[3039:3024];
      256'b?????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6114_ = b[3055:3040];
      256'b????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6114_ = b[3071:3056];
      256'b???????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6114_ = b[3087:3072];
      256'b??????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6114_ = b[3103:3088];
      256'b?????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6114_ = b[3119:3104];
      256'b????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6114_ = b[3135:3120];
      256'b???????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6114_ = b[3151:3136];
      256'b??????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6114_ = b[3167:3152];
      256'b?????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6114_ = b[3183:3168];
      256'b????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6114_ = b[3199:3184];
      256'b???????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6114_ = b[3215:3200];
      256'b??????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6114_ = b[3231:3216];
      256'b?????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6114_ = b[3247:3232];
      256'b????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6114_ = b[3263:3248];
      256'b???????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6114_ = b[3279:3264];
      256'b??????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6114_ = b[3295:3280];
      256'b?????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6114_ = b[3311:3296];
      256'b????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6114_ = b[3327:3312];
      256'b???????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6114_ = b[3343:3328];
      256'b??????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6114_ = b[3359:3344];
      256'b?????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6114_ = b[3375:3360];
      256'b????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6114_ = b[3391:3376];
      256'b???????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6114_ = b[3407:3392];
      256'b??????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6114_ = b[3423:3408];
      256'b?????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6114_ = b[3439:3424];
      256'b????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6114_ = b[3455:3440];
      256'b???????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6114_ = b[3471:3456];
      256'b??????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6114_ = b[3487:3472];
      256'b?????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6114_ = b[3503:3488];
      256'b????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6114_ = b[3519:3504];
      256'b???????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6114_ = b[3535:3520];
      256'b??????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6114_ = b[3551:3536];
      256'b?????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6114_ = b[3567:3552];
      256'b????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6114_ = b[3583:3568];
      256'b???????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6114_ = b[3599:3584];
      256'b??????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6114_ = b[3615:3600];
      256'b?????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6114_ = b[3631:3616];
      256'b????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6114_ = b[3647:3632];
      256'b???????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6114_ = b[3663:3648];
      256'b??????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6114_ = b[3679:3664];
      256'b?????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6114_ = b[3695:3680];
      256'b????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6114_ = b[3711:3696];
      256'b???????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6114_ = b[3727:3712];
      256'b??????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6114_ = b[3743:3728];
      256'b?????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6114_ = b[3759:3744];
      256'b????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6114_ = b[3775:3760];
      256'b???????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6114_ = b[3791:3776];
      256'b??????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6114_ = b[3807:3792];
      256'b?????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6114_ = b[3823:3808];
      256'b????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6114_ = b[3839:3824];
      256'b???????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6114_ = b[3855:3840];
      256'b??????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6114_ = b[3871:3856];
      256'b?????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6114_ = b[3887:3872];
      256'b????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6114_ = b[3903:3888];
      256'b???????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6114_ = b[3919:3904];
      256'b??????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6114_ = b[3935:3920];
      256'b?????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6114_ = b[3951:3936];
      256'b????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6114_ = b[3967:3952];
      256'b???????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6114_ = b[3983:3968];
      256'b??????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6114_ = b[3999:3984];
      256'b?????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6114_ = b[4015:4000];
      256'b????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6114_ = b[4031:4016];
      256'b???1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6114_ = b[4047:4032];
      256'b??1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6114_ = b[4063:4048];
      256'b?1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6114_ = b[4079:4064];
      256'b1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6114_ = b[4095:4080];
      default:
        _6114_ = a;
    endcase
  endfunction
  assign _2259_ = _6114_(density_reg0, { density_reg1, density_reg2, density_reg3, density_reg4, density_reg5, density_reg6, density_reg7, density_reg8, density_reg9, density_reg10, density_reg11, density_reg12, density_reg13, density_reg14, density_reg15, density_reg16, density_reg17, density_reg18, density_reg19, density_reg20, density_reg21, density_reg22, density_reg23, density_reg24, density_reg25, density_reg26, density_reg27, density_reg28, density_reg29, density_reg30, density_reg31, density_reg32, density_reg33, density_reg34, density_reg35, density_reg36, density_reg37, density_reg38, density_reg39, density_reg40, density_reg41, density_reg42, density_reg43, density_reg44, density_reg45, density_reg46, density_reg47, density_reg48, density_reg49, density_reg50, density_reg51, density_reg52, density_reg53, density_reg54, density_reg55, density_reg56, density_reg57, density_reg58, density_reg59, density_reg60, density_reg61, density_reg62, density_reg63, density_reg64, density_reg65, density_reg66, density_reg67, density_reg68, density_reg69, density_reg70, density_reg71, density_reg72, density_reg73, density_reg74, density_reg75, density_reg76, density_reg77, density_reg78, density_reg79, density_reg80, density_reg81, density_reg82, density_reg83, density_reg84, density_reg85, density_reg86, density_reg87, density_reg88, density_reg89, density_reg90, density_reg91, density_reg92, density_reg93, density_reg94, density_reg95, density_reg96, density_reg97, density_reg98, density_reg99, density_reg100, density_reg101, density_reg102, density_reg103, density_reg104, density_reg105, density_reg106, density_reg107, density_reg108, density_reg109, density_reg110, density_reg111, density_reg112, density_reg113, density_reg114, density_reg115, density_reg116, density_reg117, density_reg118, density_reg119, density_reg120, density_reg121, density_reg122, density_reg123, density_reg124, density_reg125, density_reg126, density_reg127, density_reg128, density_reg129, density_reg130, density_reg131, density_reg132, density_reg133, density_reg134, density_reg135, density_reg136, density_reg137, density_reg138, density_reg139, density_reg140, density_reg141, density_reg142, density_reg143, density_reg144, density_reg145, density_reg146, density_reg147, density_reg148, density_reg149, density_reg150, density_reg151, density_reg152, density_reg153, density_reg154, density_reg155, density_reg156, density_reg157, density_reg158, density_reg159, density_reg160, density_reg161, density_reg162, density_reg163, density_reg164, density_reg165, density_reg166, density_reg167, density_reg168, density_reg169, density_reg170, density_reg171, density_reg172, density_reg173, density_reg174, density_reg175, density_reg176, density_reg177, density_reg178, density_reg179, density_reg180, density_reg181, density_reg182, density_reg183, density_reg184, density_reg185, density_reg186, density_reg187, density_reg188, density_reg189, density_reg190, density_reg191, density_reg192, density_reg193, density_reg194, density_reg195, density_reg196, density_reg197, density_reg198, density_reg199, density_reg200, density_reg201, density_reg202, density_reg203, density_reg204, density_reg205, density_reg206, density_reg207, density_reg208, density_reg209, density_reg210, density_reg211, density_reg212, density_reg213, density_reg214, density_reg215, density_reg216, density_reg217, density_reg218, density_reg219, density_reg220, density_reg221, density_reg222, density_reg223, density_reg224, density_reg225, density_reg226, density_reg227, density_reg228, density_reg229, density_reg230, density_reg231, density_reg232, density_reg233, density_reg234, density_reg235, density_reg236, density_reg237, density_reg238, density_reg239, density_reg240, density_reg241, density_reg242, density_reg243, density_reg244, density_reg245, density_reg246, density_reg247, density_reg248, density_reg249, density_reg250, density_reg251, density_reg252, density_reg253, density_reg254, density_reg255, density_reg256 }, { _2516_, _2515_, _2514_, _2513_, _2512_, _2511_, _2510_, _2509_, _2508_, _2507_, _2506_, _2505_, _2504_, _2503_, _2502_, _2501_, _2500_, _2499_, _2498_, _2497_, _2496_, _2495_, _2494_, _2493_, _2492_, _2491_, _2490_, _2489_, _2488_, _2487_, _2486_, _2485_, _2484_, _2483_, _2482_, _2481_, _2480_, _2479_, _2478_, _2477_, _2476_, _2475_, _2474_, _2473_, _2472_, _2471_, _2470_, _2469_, _2468_, _2467_, _2466_, _2465_, _2464_, _2463_, _2462_, _2461_, _2460_, _2459_, _2458_, _2457_, _2456_, _2455_, _2454_, _2453_, _2452_, _2451_, _2450_, _2449_, _2448_, _2447_, _2446_, _2445_, _2444_, _2443_, _2442_, _2441_, _2440_, _2439_, _2438_, _2437_, _2436_, _2435_, _2434_, _2433_, _2432_, _2431_, _2430_, _2429_, _2428_, _2427_, _2426_, _2425_, _2424_, _2423_, _2422_, _2421_, _2420_, _2419_, _2418_, _2417_, _2416_, _2415_, _2414_, _2413_, _2412_, _2411_, _2410_, _2409_, _2408_, _2407_, _2406_, _2405_, _2404_, _2403_, _2402_, _2401_, _2400_, _2399_, _2398_, _2397_, _2396_, _2395_, _2394_, _2393_, _2392_, _2391_, _2390_, _2389_, _2388_, _2387_, _2386_, _2385_, _2384_, _2383_, _2382_, _2381_, _2380_, _2379_, _2378_, _2377_, _2376_, _2375_, _2374_, _2373_, _2372_, _2371_, _2370_, _2369_, _2368_, _2367_, _2366_, _2365_, _2364_, _2363_, _2362_, _2361_, _2360_, _2359_, _2358_, _2357_, _2356_, _2355_, _2354_, _2353_, _2352_, _2351_, _2350_, _2349_, _2348_, _2347_, _2346_, _2345_, _2344_, _2343_, _2342_, _2341_, _2340_, _2339_, _2338_, _2337_, _2336_, _2335_, _2334_, _2333_, _2332_, _2331_, _2330_, _2329_, _2328_, _2327_, _2326_, _2325_, _2324_, _2323_, _2322_, _2321_, _2320_, _2319_, _2318_, _2317_, _2316_, _2315_, _2314_, _2313_, _2312_, _2311_, _2310_, _2309_, _2308_, _2307_, _2306_, _2305_, _2304_, _2303_, _2302_, _2301_, _2300_, _2299_, _2298_, _2297_, _2296_, _2295_, _2294_, _2293_, _2292_, _2291_, _2290_, _2289_, _2288_, _2287_, _2286_, _2285_, _2284_, _2283_, _2282_, _2281_, _2280_, _2279_, _2278_, _2277_, _2276_, _2275_, _2274_, _2273_, _2272_, _2271_, _2270_, _2269_, _2268_, _2267_, _2266_, _2265_, _2264_, _2263_, _2262_, _0405_ });
  assign _2260_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9299|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 9'b100000000;
  assign _2261_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9295|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 8'b11111111;
  assign _2262_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9291|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 8'b11111110;
  assign _2263_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9287|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 8'b11111101;
  assign _2264_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9283|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 8'b11111100;
  assign _2265_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9279|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 8'b11111011;
  assign _2266_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9275|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 8'b11111010;
  assign _2267_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9271|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 8'b11111001;
  assign _2268_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9267|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 8'b11111000;
  assign _2269_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9263|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 8'b11110111;
  assign _2270_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9259|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 8'b11110110;
  assign _2271_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9255|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 8'b11110101;
  assign _2272_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9251|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 8'b11110100;
  assign _2273_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9247|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 8'b11110011;
  assign _2274_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9243|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 8'b11110010;
  assign _2275_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9239|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 8'b11110001;
  assign _2276_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9235|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 8'b11110000;
  assign _2277_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9231|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 8'b11101111;
  assign _2278_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9227|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 8'b11101110;
  assign _2279_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9223|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 8'b11101101;
  assign _2280_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9219|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 8'b11101100;
  assign _2281_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9215|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 8'b11101011;
  assign _2282_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9211|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 8'b11101010;
  assign _2283_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9207|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 8'b11101001;
  assign _2284_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9203|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 8'b11101000;
  assign _2285_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9199|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 8'b11100111;
  assign _2286_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9195|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 8'b11100110;
  assign _2287_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9191|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 8'b11100101;
  assign _2288_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9187|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 8'b11100100;
  assign _2289_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9183|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 8'b11100011;
  assign _2290_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9179|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 8'b11100010;
  assign _2291_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9175|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 8'b11100001;
  assign _2292_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9171|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 8'b11100000;
  assign _2293_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9167|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 8'b11011111;
  assign _2294_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9163|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 8'b11011110;
  assign _2295_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9159|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 8'b11011101;
  assign _2296_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9155|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 8'b11011100;
  assign _2297_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9151|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 8'b11011011;
  assign _2298_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9147|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 8'b11011010;
  assign _2299_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9143|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 8'b11011001;
  assign _2300_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9139|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 8'b11011000;
  assign _2301_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9135|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 8'b11010111;
  assign _2302_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9131|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 8'b11010110;
  assign _2303_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9127|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 8'b11010101;
  assign _2304_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9123|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 8'b11010100;
  assign _2305_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9119|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 8'b11010011;
  assign _2306_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9115|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 8'b11010010;
  assign _2307_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9111|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 8'b11010001;
  assign _2308_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9107|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 8'b11010000;
  assign _2309_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9103|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 8'b11001111;
  assign _2310_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9099|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 8'b11001110;
  assign _2311_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9095|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 8'b11001101;
  assign _2312_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9091|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 8'b11001100;
  assign _2313_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9087|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 8'b11001011;
  assign _2314_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9083|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 8'b11001010;
  assign _2315_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9079|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 8'b11001001;
  assign _2316_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9075|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 8'b11001000;
  assign _2317_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9071|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 8'b11000111;
  assign _2318_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9067|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 8'b11000110;
  assign _2319_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9063|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 8'b11000101;
  assign _2320_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9059|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 8'b11000100;
  assign _2321_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9055|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 8'b11000011;
  assign _2322_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9051|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 8'b11000010;
  assign _2323_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9047|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 8'b11000001;
  assign _2324_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9043|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 8'b11000000;
  assign _2325_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9039|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 8'b10111111;
  assign _2326_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9035|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 8'b10111110;
  assign _2327_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9031|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 8'b10111101;
  assign _2328_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9027|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 8'b10111100;
  assign _2329_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9023|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 8'b10111011;
  assign _2330_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9019|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 8'b10111010;
  assign _2331_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9015|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 8'b10111001;
  assign _2332_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9011|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 8'b10111000;
  assign _2333_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9007|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 8'b10110111;
  assign _2334_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9003|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 8'b10110110;
  assign _2335_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8999|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 8'b10110101;
  assign _2336_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8995|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 8'b10110100;
  assign _2337_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8991|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 8'b10110011;
  assign _2338_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8987|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 8'b10110010;
  assign _2339_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8983|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 8'b10110001;
  assign _2340_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8979|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 8'b10110000;
  assign _2341_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8975|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 8'b10101111;
  assign _2342_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8971|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 8'b10101110;
  assign _2343_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8967|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 8'b10101101;
  assign _2344_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8963|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 8'b10101100;
  assign _2345_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8959|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 8'b10101011;
  assign _2346_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8955|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 8'b10101010;
  assign _2347_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8951|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 8'b10101001;
  assign _2348_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8947|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 8'b10101000;
  assign _2349_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8943|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 8'b10100111;
  assign _2350_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8939|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 8'b10100110;
  assign _2351_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8935|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 8'b10100101;
  assign _2352_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8931|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 8'b10100100;
  assign _2353_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8927|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 8'b10100011;
  assign _2354_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8923|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 8'b10100010;
  assign _2355_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8919|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 8'b10100001;
  assign _2356_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8915|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 8'b10100000;
  assign _2357_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8911|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 8'b10011111;
  assign _2358_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8907|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 8'b10011110;
  assign _2359_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8903|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 8'b10011101;
  assign _2360_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8899|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 8'b10011100;
  assign _2361_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8895|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 8'b10011011;
  assign _2362_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8891|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 8'b10011010;
  assign _2363_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8887|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 8'b10011001;
  assign _2364_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8883|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 8'b10011000;
  assign _2365_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8879|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 8'b10010111;
  assign _2366_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8875|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 8'b10010110;
  assign _2367_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8871|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 8'b10010101;
  assign _2368_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8867|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 8'b10010100;
  assign _2369_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8863|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 8'b10010011;
  assign _2370_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8859|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 8'b10010010;
  assign _2371_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8855|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 8'b10010001;
  assign _2372_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8851|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 8'b10010000;
  assign _2373_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8847|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 8'b10001111;
  assign _2374_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8843|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 8'b10001110;
  assign _2375_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8839|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 8'b10001101;
  assign _2376_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8835|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 8'b10001100;
  assign _2377_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8831|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 8'b10001011;
  assign _2378_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8827|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 8'b10001010;
  assign _2379_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8823|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 8'b10001001;
  assign _2380_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8819|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 8'b10001000;
  assign _2381_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8815|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 8'b10000111;
  assign _2382_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8811|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 8'b10000110;
  assign _2383_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8807|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 8'b10000101;
  assign _2384_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8803|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 8'b10000100;
  assign _2385_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8799|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 8'b10000011;
  assign _2386_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8795|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 8'b10000010;
  assign _2387_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8791|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 8'b10000001;
  assign _2388_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8787|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 8'b10000000;
  assign _2389_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8783|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 7'b1111111;
  assign _2390_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8779|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 7'b1111110;
  assign _2391_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8775|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 7'b1111101;
  assign _2392_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8771|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 7'b1111100;
  assign _2393_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8767|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 7'b1111011;
  assign _2394_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8763|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 7'b1111010;
  assign _2395_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8759|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 7'b1111001;
  assign _2396_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8755|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 7'b1111000;
  assign _2397_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8751|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 7'b1110111;
  assign _2398_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8747|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 7'b1110110;
  assign _2399_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8743|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 7'b1110101;
  assign _2400_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8739|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 7'b1110100;
  assign _2401_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8735|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 7'b1110011;
  assign _2402_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8731|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 7'b1110010;
  assign _2403_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8727|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 7'b1110001;
  assign _2404_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8723|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 7'b1110000;
  assign _2405_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8719|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 7'b1101111;
  assign _2406_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8715|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 7'b1101110;
  assign _2407_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8711|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 7'b1101101;
  assign _2408_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8707|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 7'b1101100;
  assign _2409_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8703|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 7'b1101011;
  assign _2410_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8699|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 7'b1101010;
  assign _2411_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8695|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 7'b1101001;
  assign _2412_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8691|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 7'b1101000;
  assign _2413_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8687|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 7'b1100111;
  assign _2414_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8683|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 7'b1100110;
  assign _2415_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8679|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 7'b1100101;
  assign _2416_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8675|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 7'b1100100;
  assign _2417_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8671|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 7'b1100011;
  assign _2418_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8667|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 7'b1100010;
  assign _2419_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8663|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 7'b1100001;
  assign _2420_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8659|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 7'b1100000;
  assign _2421_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8655|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 7'b1011111;
  assign _2422_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8651|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 7'b1011110;
  assign _2423_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8647|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 7'b1011101;
  assign _2424_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8643|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 7'b1011100;
  assign _2425_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8639|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 7'b1011011;
  assign _2426_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8635|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 7'b1011010;
  assign _2427_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8631|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 7'b1011001;
  assign _2428_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8627|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 7'b1011000;
  assign _2429_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8623|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 7'b1010111;
  assign _2430_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8619|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 7'b1010110;
  assign _2431_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8615|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 7'b1010101;
  assign _2432_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8611|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 7'b1010100;
  assign _2433_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8607|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 7'b1010011;
  assign _2434_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8603|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 7'b1010010;
  assign _2435_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8599|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 7'b1010001;
  assign _2436_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8595|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 7'b1010000;
  assign _2437_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8591|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 7'b1001111;
  assign _2438_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8587|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 7'b1001110;
  assign _2439_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8583|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 7'b1001101;
  assign _2440_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8579|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 7'b1001100;
  assign _2441_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8575|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 7'b1001011;
  assign _2442_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8571|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 7'b1001010;
  assign _2443_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8567|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 7'b1001001;
  assign _2444_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8563|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 7'b1001000;
  assign _2445_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8559|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 7'b1000111;
  assign _2446_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8555|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 7'b1000110;
  assign _2447_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8551|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 7'b1000101;
  assign _2448_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8547|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 7'b1000100;
  assign _2449_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8543|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 7'b1000011;
  assign _2450_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8539|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 7'b1000010;
  assign _2451_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8535|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 7'b1000001;
  assign _2452_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8531|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 7'b1000000;
  assign _2453_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8527|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 6'b111111;
  assign _2454_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8523|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 6'b111110;
  assign _2455_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8519|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 6'b111101;
  assign _2456_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8515|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 6'b111100;
  assign _2457_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8511|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 6'b111011;
  assign _2458_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8507|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 6'b111010;
  assign _2459_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8503|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 6'b111001;
  assign _2460_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8499|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 6'b111000;
  assign _2461_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8495|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 6'b110111;
  assign _2462_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8491|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 6'b110110;
  assign _2463_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8487|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 6'b110101;
  assign _2464_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8483|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 6'b110100;
  assign _2465_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8479|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 6'b110011;
  assign _2466_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8475|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 6'b110010;
  assign _2467_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8471|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 6'b110001;
  assign _2468_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8467|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 6'b110000;
  assign _2469_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8463|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 6'b101111;
  assign _2470_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8459|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 6'b101110;
  assign _2471_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8455|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 6'b101101;
  assign _2472_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8451|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 6'b101100;
  assign _2473_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8447|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 6'b101011;
  assign _2474_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8443|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 6'b101010;
  assign _2475_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8439|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 6'b101001;
  assign _2476_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8435|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 6'b101000;
  assign _2477_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8431|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 6'b100111;
  assign _2478_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8427|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 6'b100110;
  assign _2479_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8423|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 6'b100101;
  assign _2480_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8419|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 6'b100100;
  assign _2481_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8415|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 6'b100011;
  assign _2482_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8411|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 6'b100010;
  assign _2483_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8407|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 6'b100001;
  assign _2484_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8403|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 6'b100000;
  assign _2485_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8399|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 5'b11111;
  assign _2486_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8395|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 5'b11110;
  assign _2487_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8391|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 5'b11101;
  assign _2488_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8387|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 5'b11100;
  assign _2489_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8383|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 5'b11011;
  assign _2490_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8379|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 5'b11010;
  assign _2491_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8375|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 5'b11001;
  assign _2492_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8371|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 5'b11000;
  assign _2493_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8367|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 5'b10111;
  assign _2494_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8363|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 5'b10110;
  assign _2495_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8359|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 5'b10101;
  assign _2496_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8355|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 5'b10100;
  assign _2497_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8351|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 5'b10011;
  assign _2498_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8347|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 5'b10010;
  assign _2499_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8343|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 5'b10001;
  assign _2500_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8339|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 5'b10000;
  assign _2501_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8335|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 4'b1111;
  assign _2502_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8331|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 4'b1110;
  assign _2503_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8327|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 4'b1101;
  assign _2504_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8323|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 4'b1100;
  assign _2505_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8319|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 4'b1011;
  assign _2506_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8315|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 4'b1010;
  assign _2507_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8311|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 4'b1001;
  assign _2508_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8307|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 4'b1000;
  assign _2509_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8303|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 3'b111;
  assign _2510_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8299|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 3'b110;
  assign _2511_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8295|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 3'b101;
  assign _2512_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8291|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 3'b100;
  assign _2513_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8287|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 2'b11;
  assign _2514_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8283|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 2'b10;
  assign _2515_ = dp2lut_Y_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8279|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) 1'b1;
  assign _2516_ = ! (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8275|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *) dp2lut_Y_entry_1;
  assign _2517_ = dp2lut_Yinfo_1[17] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8270" *) density_reg256 : _2259_;
  assign _2518_ = dp2lut_Yinfo_1[16] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8267" *) density_reg0 : _2517_;
  assign _0288_ = _0401_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8266" *) _2518_ : lut_Y_data_11;
  function [15:0] _6375_;
    input [15:0] a;
    input [4095:0] b;
    input [255:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:9299|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8274" *)
    (* parallel_case *)
    casez (s)
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1:
        _6375_ = b[15:0];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?:
        _6375_ = b[31:16];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??:
        _6375_ = b[47:32];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???:
        _6375_ = b[63:48];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????:
        _6375_ = b[79:64];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????:
        _6375_ = b[95:80];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????:
        _6375_ = b[111:96];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????:
        _6375_ = b[127:112];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????:
        _6375_ = b[143:128];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????:
        _6375_ = b[159:144];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????:
        _6375_ = b[175:160];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????:
        _6375_ = b[191:176];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????:
        _6375_ = b[207:192];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????:
        _6375_ = b[223:208];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????:
        _6375_ = b[239:224];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????:
        _6375_ = b[255:240];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????:
        _6375_ = b[271:256];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????:
        _6375_ = b[287:272];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????:
        _6375_ = b[303:288];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????:
        _6375_ = b[319:304];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????:
        _6375_ = b[335:320];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????:
        _6375_ = b[351:336];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????:
        _6375_ = b[367:352];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????:
        _6375_ = b[383:368];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????:
        _6375_ = b[399:384];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????:
        _6375_ = b[415:400];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????:
        _6375_ = b[431:416];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????:
        _6375_ = b[447:432];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????:
        _6375_ = b[463:448];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????:
        _6375_ = b[479:464];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????:
        _6375_ = b[495:480];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????:
        _6375_ = b[511:496];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????:
        _6375_ = b[527:512];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????:
        _6375_ = b[543:528];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????:
        _6375_ = b[559:544];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????:
        _6375_ = b[575:560];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????:
        _6375_ = b[591:576];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????:
        _6375_ = b[607:592];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????:
        _6375_ = b[623:608];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????:
        _6375_ = b[639:624];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????:
        _6375_ = b[655:640];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????:
        _6375_ = b[671:656];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????:
        _6375_ = b[687:672];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????:
        _6375_ = b[703:688];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????:
        _6375_ = b[719:704];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????:
        _6375_ = b[735:720];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????:
        _6375_ = b[751:736];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????:
        _6375_ = b[767:752];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????:
        _6375_ = b[783:768];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????:
        _6375_ = b[799:784];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????:
        _6375_ = b[815:800];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????:
        _6375_ = b[831:816];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????:
        _6375_ = b[847:832];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????:
        _6375_ = b[863:848];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????:
        _6375_ = b[879:864];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????:
        _6375_ = b[895:880];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????:
        _6375_ = b[911:896];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????:
        _6375_ = b[927:912];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????:
        _6375_ = b[943:928];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????:
        _6375_ = b[959:944];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????:
        _6375_ = b[975:960];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????:
        _6375_ = b[991:976];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????:
        _6375_ = b[1007:992];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????:
        _6375_ = b[1023:1008];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????:
        _6375_ = b[1039:1024];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????:
        _6375_ = b[1055:1040];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????:
        _6375_ = b[1071:1056];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????:
        _6375_ = b[1087:1072];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????:
        _6375_ = b[1103:1088];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????:
        _6375_ = b[1119:1104];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????:
        _6375_ = b[1135:1120];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????:
        _6375_ = b[1151:1136];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????:
        _6375_ = b[1167:1152];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????:
        _6375_ = b[1183:1168];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????:
        _6375_ = b[1199:1184];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????:
        _6375_ = b[1215:1200];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????:
        _6375_ = b[1231:1216];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????:
        _6375_ = b[1247:1232];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????:
        _6375_ = b[1263:1248];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????:
        _6375_ = b[1279:1264];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????:
        _6375_ = b[1295:1280];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????:
        _6375_ = b[1311:1296];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????:
        _6375_ = b[1327:1312];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????:
        _6375_ = b[1343:1328];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????:
        _6375_ = b[1359:1344];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????:
        _6375_ = b[1375:1360];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????:
        _6375_ = b[1391:1376];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????:
        _6375_ = b[1407:1392];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????:
        _6375_ = b[1423:1408];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????:
        _6375_ = b[1439:1424];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????:
        _6375_ = b[1455:1440];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????:
        _6375_ = b[1471:1456];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????:
        _6375_ = b[1487:1472];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????:
        _6375_ = b[1503:1488];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????:
        _6375_ = b[1519:1504];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????:
        _6375_ = b[1535:1520];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????:
        _6375_ = b[1551:1536];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????:
        _6375_ = b[1567:1552];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????:
        _6375_ = b[1583:1568];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????:
        _6375_ = b[1599:1584];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6375_ = b[1615:1600];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6375_ = b[1631:1616];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6375_ = b[1647:1632];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6375_ = b[1663:1648];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6375_ = b[1679:1664];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6375_ = b[1695:1680];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6375_ = b[1711:1696];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6375_ = b[1727:1712];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6375_ = b[1743:1728];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6375_ = b[1759:1744];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6375_ = b[1775:1760];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6375_ = b[1791:1776];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6375_ = b[1807:1792];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6375_ = b[1823:1808];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6375_ = b[1839:1824];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6375_ = b[1855:1840];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6375_ = b[1871:1856];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6375_ = b[1887:1872];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6375_ = b[1903:1888];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6375_ = b[1919:1904];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6375_ = b[1935:1920];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6375_ = b[1951:1936];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6375_ = b[1967:1952];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6375_ = b[1983:1968];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6375_ = b[1999:1984];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6375_ = b[2015:2000];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6375_ = b[2031:2016];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6375_ = b[2047:2032];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6375_ = b[2063:2048];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6375_ = b[2079:2064];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6375_ = b[2095:2080];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6375_ = b[2111:2096];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6375_ = b[2127:2112];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6375_ = b[2143:2128];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6375_ = b[2159:2144];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6375_ = b[2175:2160];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6375_ = b[2191:2176];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6375_ = b[2207:2192];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6375_ = b[2223:2208];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6375_ = b[2239:2224];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6375_ = b[2255:2240];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6375_ = b[2271:2256];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6375_ = b[2287:2272];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6375_ = b[2303:2288];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6375_ = b[2319:2304];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6375_ = b[2335:2320];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6375_ = b[2351:2336];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6375_ = b[2367:2352];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6375_ = b[2383:2368];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6375_ = b[2399:2384];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6375_ = b[2415:2400];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6375_ = b[2431:2416];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6375_ = b[2447:2432];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6375_ = b[2463:2448];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6375_ = b[2479:2464];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6375_ = b[2495:2480];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6375_ = b[2511:2496];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6375_ = b[2527:2512];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6375_ = b[2543:2528];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6375_ = b[2559:2544];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6375_ = b[2575:2560];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6375_ = b[2591:2576];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6375_ = b[2607:2592];
      256'b????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6375_ = b[2623:2608];
      256'b???????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6375_ = b[2639:2624];
      256'b??????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6375_ = b[2655:2640];
      256'b?????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6375_ = b[2671:2656];
      256'b????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6375_ = b[2687:2672];
      256'b???????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6375_ = b[2703:2688];
      256'b??????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6375_ = b[2719:2704];
      256'b?????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6375_ = b[2735:2720];
      256'b????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6375_ = b[2751:2736];
      256'b???????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6375_ = b[2767:2752];
      256'b??????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6375_ = b[2783:2768];
      256'b?????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6375_ = b[2799:2784];
      256'b????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6375_ = b[2815:2800];
      256'b???????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6375_ = b[2831:2816];
      256'b??????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6375_ = b[2847:2832];
      256'b?????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6375_ = b[2863:2848];
      256'b????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6375_ = b[2879:2864];
      256'b???????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6375_ = b[2895:2880];
      256'b??????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6375_ = b[2911:2896];
      256'b?????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6375_ = b[2927:2912];
      256'b????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6375_ = b[2943:2928];
      256'b???????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6375_ = b[2959:2944];
      256'b??????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6375_ = b[2975:2960];
      256'b?????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6375_ = b[2991:2976];
      256'b????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6375_ = b[3007:2992];
      256'b???????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6375_ = b[3023:3008];
      256'b??????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6375_ = b[3039:3024];
      256'b?????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6375_ = b[3055:3040];
      256'b????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6375_ = b[3071:3056];
      256'b???????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6375_ = b[3087:3072];
      256'b??????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6375_ = b[3103:3088];
      256'b?????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6375_ = b[3119:3104];
      256'b????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6375_ = b[3135:3120];
      256'b???????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6375_ = b[3151:3136];
      256'b??????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6375_ = b[3167:3152];
      256'b?????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6375_ = b[3183:3168];
      256'b????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6375_ = b[3199:3184];
      256'b???????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6375_ = b[3215:3200];
      256'b??????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6375_ = b[3231:3216];
      256'b?????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6375_ = b[3247:3232];
      256'b????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6375_ = b[3263:3248];
      256'b???????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6375_ = b[3279:3264];
      256'b??????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6375_ = b[3295:3280];
      256'b?????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6375_ = b[3311:3296];
      256'b????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6375_ = b[3327:3312];
      256'b???????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6375_ = b[3343:3328];
      256'b??????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6375_ = b[3359:3344];
      256'b?????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6375_ = b[3375:3360];
      256'b????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6375_ = b[3391:3376];
      256'b???????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6375_ = b[3407:3392];
      256'b??????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6375_ = b[3423:3408];
      256'b?????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6375_ = b[3439:3424];
      256'b????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6375_ = b[3455:3440];
      256'b???????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6375_ = b[3471:3456];
      256'b??????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6375_ = b[3487:3472];
      256'b?????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6375_ = b[3503:3488];
      256'b????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6375_ = b[3519:3504];
      256'b???????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6375_ = b[3535:3520];
      256'b??????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6375_ = b[3551:3536];
      256'b?????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6375_ = b[3567:3552];
      256'b????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6375_ = b[3583:3568];
      256'b???????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6375_ = b[3599:3584];
      256'b??????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6375_ = b[3615:3600];
      256'b?????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6375_ = b[3631:3616];
      256'b????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6375_ = b[3647:3632];
      256'b???????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6375_ = b[3663:3648];
      256'b??????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6375_ = b[3679:3664];
      256'b?????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6375_ = b[3695:3680];
      256'b????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6375_ = b[3711:3696];
      256'b???????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6375_ = b[3727:3712];
      256'b??????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6375_ = b[3743:3728];
      256'b?????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6375_ = b[3759:3744];
      256'b????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6375_ = b[3775:3760];
      256'b???????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6375_ = b[3791:3776];
      256'b??????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6375_ = b[3807:3792];
      256'b?????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6375_ = b[3823:3808];
      256'b????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6375_ = b[3839:3824];
      256'b???????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6375_ = b[3855:3840];
      256'b??????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6375_ = b[3871:3856];
      256'b?????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6375_ = b[3887:3872];
      256'b????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6375_ = b[3903:3888];
      256'b???????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6375_ = b[3919:3904];
      256'b??????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6375_ = b[3935:3920];
      256'b?????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6375_ = b[3951:3936];
      256'b????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6375_ = b[3967:3952];
      256'b???????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6375_ = b[3983:3968];
      256'b??????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6375_ = b[3999:3984];
      256'b?????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6375_ = b[4015:4000];
      256'b????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6375_ = b[4031:4016];
      256'b???1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6375_ = b[4047:4032];
      256'b??1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6375_ = b[4063:4048];
      256'b?1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6375_ = b[4079:4064];
      256'b1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6375_ = b[4095:4080];
      default:
        _6375_ = a;
    endcase
  endfunction
  assign _2519_ = _6375_(density_reg0, { density_reg1, density_reg2, density_reg3, density_reg4, density_reg5, density_reg6, density_reg7, density_reg8, density_reg9, density_reg10, density_reg11, density_reg12, density_reg13, density_reg14, density_reg15, density_reg16, density_reg17, density_reg18, density_reg19, density_reg20, density_reg21, density_reg22, density_reg23, density_reg24, density_reg25, density_reg26, density_reg27, density_reg28, density_reg29, density_reg30, density_reg31, density_reg32, density_reg33, density_reg34, density_reg35, density_reg36, density_reg37, density_reg38, density_reg39, density_reg40, density_reg41, density_reg42, density_reg43, density_reg44, density_reg45, density_reg46, density_reg47, density_reg48, density_reg49, density_reg50, density_reg51, density_reg52, density_reg53, density_reg54, density_reg55, density_reg56, density_reg57, density_reg58, density_reg59, density_reg60, density_reg61, density_reg62, density_reg63, density_reg64, density_reg65, density_reg66, density_reg67, density_reg68, density_reg69, density_reg70, density_reg71, density_reg72, density_reg73, density_reg74, density_reg75, density_reg76, density_reg77, density_reg78, density_reg79, density_reg80, density_reg81, density_reg82, density_reg83, density_reg84, density_reg85, density_reg86, density_reg87, density_reg88, density_reg89, density_reg90, density_reg91, density_reg92, density_reg93, density_reg94, density_reg95, density_reg96, density_reg97, density_reg98, density_reg99, density_reg100, density_reg101, density_reg102, density_reg103, density_reg104, density_reg105, density_reg106, density_reg107, density_reg108, density_reg109, density_reg110, density_reg111, density_reg112, density_reg113, density_reg114, density_reg115, density_reg116, density_reg117, density_reg118, density_reg119, density_reg120, density_reg121, density_reg122, density_reg123, density_reg124, density_reg125, density_reg126, density_reg127, density_reg128, density_reg129, density_reg130, density_reg131, density_reg132, density_reg133, density_reg134, density_reg135, density_reg136, density_reg137, density_reg138, density_reg139, density_reg140, density_reg141, density_reg142, density_reg143, density_reg144, density_reg145, density_reg146, density_reg147, density_reg148, density_reg149, density_reg150, density_reg151, density_reg152, density_reg153, density_reg154, density_reg155, density_reg156, density_reg157, density_reg158, density_reg159, density_reg160, density_reg161, density_reg162, density_reg163, density_reg164, density_reg165, density_reg166, density_reg167, density_reg168, density_reg169, density_reg170, density_reg171, density_reg172, density_reg173, density_reg174, density_reg175, density_reg176, density_reg177, density_reg178, density_reg179, density_reg180, density_reg181, density_reg182, density_reg183, density_reg184, density_reg185, density_reg186, density_reg187, density_reg188, density_reg189, density_reg190, density_reg191, density_reg192, density_reg193, density_reg194, density_reg195, density_reg196, density_reg197, density_reg198, density_reg199, density_reg200, density_reg201, density_reg202, density_reg203, density_reg204, density_reg205, density_reg206, density_reg207, density_reg208, density_reg209, density_reg210, density_reg211, density_reg212, density_reg213, density_reg214, density_reg215, density_reg216, density_reg217, density_reg218, density_reg219, density_reg220, density_reg221, density_reg222, density_reg223, density_reg224, density_reg225, density_reg226, density_reg227, density_reg228, density_reg229, density_reg230, density_reg231, density_reg232, density_reg233, density_reg234, density_reg235, density_reg236, density_reg237, density_reg238, density_reg239, density_reg240, density_reg241, density_reg242, density_reg243, density_reg244, density_reg245, density_reg246, density_reg247, density_reg248, density_reg249, density_reg250, density_reg251, density_reg252, density_reg253, density_reg254, density_reg255, density_reg256 }, { _2515_, _2514_, _2513_, _2512_, _2511_, _2510_, _2509_, _2508_, _2507_, _2506_, _2505_, _2504_, _2503_, _2502_, _2501_, _2500_, _2499_, _2498_, _2497_, _2496_, _2495_, _2494_, _2493_, _2492_, _2491_, _2490_, _2489_, _2488_, _2487_, _2486_, _2485_, _2484_, _2483_, _2482_, _2481_, _2480_, _2479_, _2478_, _2477_, _2476_, _2475_, _2474_, _2473_, _2472_, _2471_, _2470_, _2469_, _2468_, _2467_, _2466_, _2465_, _2464_, _2463_, _2462_, _2461_, _2460_, _2459_, _2458_, _2457_, _2456_, _2455_, _2454_, _2453_, _2452_, _2451_, _2450_, _2449_, _2448_, _2447_, _2446_, _2445_, _2444_, _2443_, _2442_, _2441_, _2440_, _2439_, _2438_, _2437_, _2436_, _2435_, _2434_, _2433_, _2432_, _2431_, _2430_, _2429_, _2428_, _2427_, _2426_, _2425_, _2424_, _2423_, _2422_, _2421_, _2420_, _2419_, _2418_, _2417_, _2416_, _2415_, _2414_, _2413_, _2412_, _2411_, _2410_, _2409_, _2408_, _2407_, _2406_, _2405_, _2404_, _2403_, _2402_, _2401_, _2400_, _2399_, _2398_, _2397_, _2396_, _2395_, _2394_, _2393_, _2392_, _2391_, _2390_, _2389_, _2388_, _2387_, _2386_, _2385_, _2384_, _2383_, _2382_, _2381_, _2380_, _2379_, _2378_, _2377_, _2376_, _2375_, _2374_, _2373_, _2372_, _2371_, _2370_, _2369_, _2368_, _2367_, _2366_, _2365_, _2364_, _2363_, _2362_, _2361_, _2360_, _2359_, _2358_, _2357_, _2356_, _2355_, _2354_, _2353_, _2352_, _2351_, _2350_, _2349_, _2348_, _2347_, _2346_, _2345_, _2344_, _2343_, _2342_, _2341_, _2340_, _2339_, _2338_, _2337_, _2336_, _2335_, _2334_, _2333_, _2332_, _2331_, _2330_, _2329_, _2328_, _2327_, _2326_, _2325_, _2324_, _2323_, _2322_, _2321_, _2320_, _2319_, _2318_, _2317_, _2316_, _2315_, _2314_, _2313_, _2312_, _2311_, _2310_, _2309_, _2308_, _2307_, _2306_, _2305_, _2304_, _2303_, _2302_, _2301_, _2300_, _2299_, _2298_, _2297_, _2296_, _2295_, _2294_, _2293_, _2292_, _2291_, _2290_, _2289_, _2288_, _2287_, _2286_, _2285_, _2284_, _2283_, _2282_, _2281_, _2280_, _2279_, _2278_, _2277_, _2276_, _2275_, _2274_, _2273_, _2272_, _2271_, _2270_, _2269_, _2268_, _2267_, _2266_, _2265_, _2264_, _2263_, _2262_, _2261_, _2260_ });
  assign _2520_ = dp2lut_Yinfo_1[17] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8270" *) density_reg256 : _2519_;
  assign _2521_ = dp2lut_Yinfo_1[16] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8267" *) density_reg0 : _2520_;
  assign _0287_ = _0401_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8266" *) _2521_ : lut_Y_data_10;
  function [15:0] _6379_;
    input [15:0] a;
    input [4095:0] b;
    input [255:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8248|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *)
    (* parallel_case *)
    casez (s)
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1:
        _6379_ = b[15:0];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?:
        _6379_ = b[31:16];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??:
        _6379_ = b[47:32];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???:
        _6379_ = b[63:48];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????:
        _6379_ = b[79:64];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????:
        _6379_ = b[95:80];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????:
        _6379_ = b[111:96];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????:
        _6379_ = b[127:112];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????:
        _6379_ = b[143:128];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????:
        _6379_ = b[159:144];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????:
        _6379_ = b[175:160];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????:
        _6379_ = b[191:176];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????:
        _6379_ = b[207:192];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????:
        _6379_ = b[223:208];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????:
        _6379_ = b[239:224];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????:
        _6379_ = b[255:240];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????:
        _6379_ = b[271:256];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????:
        _6379_ = b[287:272];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????:
        _6379_ = b[303:288];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????:
        _6379_ = b[319:304];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????:
        _6379_ = b[335:320];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????:
        _6379_ = b[351:336];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????:
        _6379_ = b[367:352];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????:
        _6379_ = b[383:368];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????:
        _6379_ = b[399:384];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????:
        _6379_ = b[415:400];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????:
        _6379_ = b[431:416];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????:
        _6379_ = b[447:432];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????:
        _6379_ = b[463:448];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????:
        _6379_ = b[479:464];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????:
        _6379_ = b[495:480];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????:
        _6379_ = b[511:496];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????:
        _6379_ = b[527:512];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????:
        _6379_ = b[543:528];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????:
        _6379_ = b[559:544];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????:
        _6379_ = b[575:560];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????:
        _6379_ = b[591:576];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????:
        _6379_ = b[607:592];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????:
        _6379_ = b[623:608];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????:
        _6379_ = b[639:624];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????:
        _6379_ = b[655:640];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????:
        _6379_ = b[671:656];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????:
        _6379_ = b[687:672];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????:
        _6379_ = b[703:688];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????:
        _6379_ = b[719:704];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????:
        _6379_ = b[735:720];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????:
        _6379_ = b[751:736];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????:
        _6379_ = b[767:752];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????:
        _6379_ = b[783:768];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????:
        _6379_ = b[799:784];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????:
        _6379_ = b[815:800];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????:
        _6379_ = b[831:816];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????:
        _6379_ = b[847:832];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????:
        _6379_ = b[863:848];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????:
        _6379_ = b[879:864];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????:
        _6379_ = b[895:880];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????:
        _6379_ = b[911:896];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????:
        _6379_ = b[927:912];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????:
        _6379_ = b[943:928];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????:
        _6379_ = b[959:944];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????:
        _6379_ = b[975:960];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????:
        _6379_ = b[991:976];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????:
        _6379_ = b[1007:992];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????:
        _6379_ = b[1023:1008];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????:
        _6379_ = b[1039:1024];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????:
        _6379_ = b[1055:1040];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????:
        _6379_ = b[1071:1056];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????:
        _6379_ = b[1087:1072];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????:
        _6379_ = b[1103:1088];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????:
        _6379_ = b[1119:1104];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????:
        _6379_ = b[1135:1120];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????:
        _6379_ = b[1151:1136];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????:
        _6379_ = b[1167:1152];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????:
        _6379_ = b[1183:1168];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????:
        _6379_ = b[1199:1184];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????:
        _6379_ = b[1215:1200];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????:
        _6379_ = b[1231:1216];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????:
        _6379_ = b[1247:1232];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????:
        _6379_ = b[1263:1248];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????:
        _6379_ = b[1279:1264];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????:
        _6379_ = b[1295:1280];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????:
        _6379_ = b[1311:1296];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????:
        _6379_ = b[1327:1312];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????:
        _6379_ = b[1343:1328];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????:
        _6379_ = b[1359:1344];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????:
        _6379_ = b[1375:1360];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????:
        _6379_ = b[1391:1376];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????:
        _6379_ = b[1407:1392];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????:
        _6379_ = b[1423:1408];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????:
        _6379_ = b[1439:1424];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????:
        _6379_ = b[1455:1440];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????:
        _6379_ = b[1471:1456];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????:
        _6379_ = b[1487:1472];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????:
        _6379_ = b[1503:1488];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????:
        _6379_ = b[1519:1504];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????:
        _6379_ = b[1535:1520];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????:
        _6379_ = b[1551:1536];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????:
        _6379_ = b[1567:1552];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????:
        _6379_ = b[1583:1568];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????:
        _6379_ = b[1599:1584];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6379_ = b[1615:1600];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6379_ = b[1631:1616];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6379_ = b[1647:1632];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6379_ = b[1663:1648];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6379_ = b[1679:1664];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6379_ = b[1695:1680];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6379_ = b[1711:1696];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6379_ = b[1727:1712];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6379_ = b[1743:1728];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6379_ = b[1759:1744];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6379_ = b[1775:1760];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6379_ = b[1791:1776];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6379_ = b[1807:1792];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6379_ = b[1823:1808];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6379_ = b[1839:1824];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6379_ = b[1855:1840];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6379_ = b[1871:1856];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6379_ = b[1887:1872];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6379_ = b[1903:1888];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6379_ = b[1919:1904];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6379_ = b[1935:1920];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6379_ = b[1951:1936];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6379_ = b[1967:1952];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6379_ = b[1983:1968];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6379_ = b[1999:1984];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6379_ = b[2015:2000];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6379_ = b[2031:2016];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6379_ = b[2047:2032];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6379_ = b[2063:2048];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6379_ = b[2079:2064];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6379_ = b[2095:2080];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6379_ = b[2111:2096];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6379_ = b[2127:2112];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6379_ = b[2143:2128];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6379_ = b[2159:2144];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6379_ = b[2175:2160];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6379_ = b[2191:2176];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6379_ = b[2207:2192];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6379_ = b[2223:2208];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6379_ = b[2239:2224];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6379_ = b[2255:2240];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6379_ = b[2271:2256];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6379_ = b[2287:2272];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6379_ = b[2303:2288];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6379_ = b[2319:2304];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6379_ = b[2335:2320];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6379_ = b[2351:2336];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6379_ = b[2367:2352];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6379_ = b[2383:2368];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6379_ = b[2399:2384];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6379_ = b[2415:2400];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6379_ = b[2431:2416];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6379_ = b[2447:2432];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6379_ = b[2463:2448];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6379_ = b[2479:2464];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6379_ = b[2495:2480];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6379_ = b[2511:2496];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6379_ = b[2527:2512];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6379_ = b[2543:2528];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6379_ = b[2559:2544];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6379_ = b[2575:2560];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6379_ = b[2591:2576];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6379_ = b[2607:2592];
      256'b????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6379_ = b[2623:2608];
      256'b???????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6379_ = b[2639:2624];
      256'b??????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6379_ = b[2655:2640];
      256'b?????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6379_ = b[2671:2656];
      256'b????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6379_ = b[2687:2672];
      256'b???????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6379_ = b[2703:2688];
      256'b??????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6379_ = b[2719:2704];
      256'b?????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6379_ = b[2735:2720];
      256'b????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6379_ = b[2751:2736];
      256'b???????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6379_ = b[2767:2752];
      256'b??????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6379_ = b[2783:2768];
      256'b?????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6379_ = b[2799:2784];
      256'b????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6379_ = b[2815:2800];
      256'b???????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6379_ = b[2831:2816];
      256'b??????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6379_ = b[2847:2832];
      256'b?????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6379_ = b[2863:2848];
      256'b????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6379_ = b[2879:2864];
      256'b???????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6379_ = b[2895:2880];
      256'b??????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6379_ = b[2911:2896];
      256'b?????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6379_ = b[2927:2912];
      256'b????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6379_ = b[2943:2928];
      256'b???????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6379_ = b[2959:2944];
      256'b??????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6379_ = b[2975:2960];
      256'b?????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6379_ = b[2991:2976];
      256'b????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6379_ = b[3007:2992];
      256'b???????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6379_ = b[3023:3008];
      256'b??????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6379_ = b[3039:3024];
      256'b?????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6379_ = b[3055:3040];
      256'b????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6379_ = b[3071:3056];
      256'b???????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6379_ = b[3087:3072];
      256'b??????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6379_ = b[3103:3088];
      256'b?????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6379_ = b[3119:3104];
      256'b????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6379_ = b[3135:3120];
      256'b???????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6379_ = b[3151:3136];
      256'b??????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6379_ = b[3167:3152];
      256'b?????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6379_ = b[3183:3168];
      256'b????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6379_ = b[3199:3184];
      256'b???????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6379_ = b[3215:3200];
      256'b??????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6379_ = b[3231:3216];
      256'b?????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6379_ = b[3247:3232];
      256'b????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6379_ = b[3263:3248];
      256'b???????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6379_ = b[3279:3264];
      256'b??????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6379_ = b[3295:3280];
      256'b?????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6379_ = b[3311:3296];
      256'b????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6379_ = b[3327:3312];
      256'b???????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6379_ = b[3343:3328];
      256'b??????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6379_ = b[3359:3344];
      256'b?????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6379_ = b[3375:3360];
      256'b????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6379_ = b[3391:3376];
      256'b???????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6379_ = b[3407:3392];
      256'b??????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6379_ = b[3423:3408];
      256'b?????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6379_ = b[3439:3424];
      256'b????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6379_ = b[3455:3440];
      256'b???????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6379_ = b[3471:3456];
      256'b??????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6379_ = b[3487:3472];
      256'b?????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6379_ = b[3503:3488];
      256'b????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6379_ = b[3519:3504];
      256'b???????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6379_ = b[3535:3520];
      256'b??????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6379_ = b[3551:3536];
      256'b?????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6379_ = b[3567:3552];
      256'b????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6379_ = b[3583:3568];
      256'b???????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6379_ = b[3599:3584];
      256'b??????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6379_ = b[3615:3600];
      256'b?????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6379_ = b[3631:3616];
      256'b????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6379_ = b[3647:3632];
      256'b???????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6379_ = b[3663:3648];
      256'b??????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6379_ = b[3679:3664];
      256'b?????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6379_ = b[3695:3680];
      256'b????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6379_ = b[3711:3696];
      256'b???????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6379_ = b[3727:3712];
      256'b??????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6379_ = b[3743:3728];
      256'b?????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6379_ = b[3759:3744];
      256'b????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6379_ = b[3775:3760];
      256'b???????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6379_ = b[3791:3776];
      256'b??????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6379_ = b[3807:3792];
      256'b?????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6379_ = b[3823:3808];
      256'b????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6379_ = b[3839:3824];
      256'b???????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6379_ = b[3855:3840];
      256'b??????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6379_ = b[3871:3856];
      256'b?????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6379_ = b[3887:3872];
      256'b????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6379_ = b[3903:3888];
      256'b???????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6379_ = b[3919:3904];
      256'b??????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6379_ = b[3935:3920];
      256'b?????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6379_ = b[3951:3936];
      256'b????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6379_ = b[3967:3952];
      256'b???????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6379_ = b[3983:3968];
      256'b??????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6379_ = b[3999:3984];
      256'b?????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6379_ = b[4015:4000];
      256'b????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6379_ = b[4031:4016];
      256'b???1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6379_ = b[4047:4032];
      256'b??1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6379_ = b[4063:4048];
      256'b?1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6379_ = b[4079:4064];
      256'b1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6379_ = b[4095:4080];
      default:
        _6379_ = a;
    endcase
  endfunction
  assign _2522_ = _6379_(density_reg0, { density_reg1, density_reg2, density_reg3, density_reg4, density_reg5, density_reg6, density_reg7, density_reg8, density_reg9, density_reg10, density_reg11, density_reg12, density_reg13, density_reg14, density_reg15, density_reg16, density_reg17, density_reg18, density_reg19, density_reg20, density_reg21, density_reg22, density_reg23, density_reg24, density_reg25, density_reg26, density_reg27, density_reg28, density_reg29, density_reg30, density_reg31, density_reg32, density_reg33, density_reg34, density_reg35, density_reg36, density_reg37, density_reg38, density_reg39, density_reg40, density_reg41, density_reg42, density_reg43, density_reg44, density_reg45, density_reg46, density_reg47, density_reg48, density_reg49, density_reg50, density_reg51, density_reg52, density_reg53, density_reg54, density_reg55, density_reg56, density_reg57, density_reg58, density_reg59, density_reg60, density_reg61, density_reg62, density_reg63, density_reg64, density_reg65, density_reg66, density_reg67, density_reg68, density_reg69, density_reg70, density_reg71, density_reg72, density_reg73, density_reg74, density_reg75, density_reg76, density_reg77, density_reg78, density_reg79, density_reg80, density_reg81, density_reg82, density_reg83, density_reg84, density_reg85, density_reg86, density_reg87, density_reg88, density_reg89, density_reg90, density_reg91, density_reg92, density_reg93, density_reg94, density_reg95, density_reg96, density_reg97, density_reg98, density_reg99, density_reg100, density_reg101, density_reg102, density_reg103, density_reg104, density_reg105, density_reg106, density_reg107, density_reg108, density_reg109, density_reg110, density_reg111, density_reg112, density_reg113, density_reg114, density_reg115, density_reg116, density_reg117, density_reg118, density_reg119, density_reg120, density_reg121, density_reg122, density_reg123, density_reg124, density_reg125, density_reg126, density_reg127, density_reg128, density_reg129, density_reg130, density_reg131, density_reg132, density_reg133, density_reg134, density_reg135, density_reg136, density_reg137, density_reg138, density_reg139, density_reg140, density_reg141, density_reg142, density_reg143, density_reg144, density_reg145, density_reg146, density_reg147, density_reg148, density_reg149, density_reg150, density_reg151, density_reg152, density_reg153, density_reg154, density_reg155, density_reg156, density_reg157, density_reg158, density_reg159, density_reg160, density_reg161, density_reg162, density_reg163, density_reg164, density_reg165, density_reg166, density_reg167, density_reg168, density_reg169, density_reg170, density_reg171, density_reg172, density_reg173, density_reg174, density_reg175, density_reg176, density_reg177, density_reg178, density_reg179, density_reg180, density_reg181, density_reg182, density_reg183, density_reg184, density_reg185, density_reg186, density_reg187, density_reg188, density_reg189, density_reg190, density_reg191, density_reg192, density_reg193, density_reg194, density_reg195, density_reg196, density_reg197, density_reg198, density_reg199, density_reg200, density_reg201, density_reg202, density_reg203, density_reg204, density_reg205, density_reg206, density_reg207, density_reg208, density_reg209, density_reg210, density_reg211, density_reg212, density_reg213, density_reg214, density_reg215, density_reg216, density_reg217, density_reg218, density_reg219, density_reg220, density_reg221, density_reg222, density_reg223, density_reg224, density_reg225, density_reg226, density_reg227, density_reg228, density_reg229, density_reg230, density_reg231, density_reg232, density_reg233, density_reg234, density_reg235, density_reg236, density_reg237, density_reg238, density_reg239, density_reg240, density_reg241, density_reg242, density_reg243, density_reg244, density_reg245, density_reg246, density_reg247, density_reg248, density_reg249, density_reg250, density_reg251, density_reg252, density_reg253, density_reg254, density_reg255, density_reg256 }, { _2779_, _2778_, _2777_, _2776_, _2775_, _2774_, _2773_, _2772_, _2771_, _2770_, _2769_, _2768_, _2767_, _2766_, _2765_, _2764_, _2763_, _2762_, _2761_, _2760_, _2759_, _2758_, _2757_, _2756_, _2755_, _2754_, _2753_, _2752_, _2751_, _2750_, _2749_, _2748_, _2747_, _2746_, _2745_, _2744_, _2743_, _2742_, _2741_, _2740_, _2739_, _2738_, _2737_, _2736_, _2735_, _2734_, _2733_, _2732_, _2731_, _2730_, _2729_, _2728_, _2727_, _2726_, _2725_, _2724_, _2723_, _2722_, _2721_, _2720_, _2719_, _2718_, _2717_, _2716_, _2715_, _2714_, _2713_, _2712_, _2711_, _2710_, _2709_, _2708_, _2707_, _2706_, _2705_, _2704_, _2703_, _2702_, _2701_, _2700_, _2699_, _2698_, _2697_, _2696_, _2695_, _2694_, _2693_, _2692_, _2691_, _2690_, _2689_, _2688_, _2687_, _2686_, _2685_, _2684_, _2683_, _2682_, _2681_, _2680_, _2679_, _2678_, _2677_, _2676_, _2675_, _2674_, _2673_, _2672_, _2671_, _2670_, _2669_, _2668_, _2667_, _2666_, _2665_, _2664_, _2663_, _2662_, _2661_, _2660_, _2659_, _2658_, _2657_, _2656_, _2655_, _2654_, _2653_, _2652_, _2651_, _2650_, _2649_, _2648_, _2647_, _2646_, _2645_, _2644_, _2643_, _2642_, _2641_, _2640_, _2639_, _2638_, _2637_, _2636_, _2635_, _2634_, _2633_, _2632_, _2631_, _2630_, _2629_, _2628_, _2627_, _2626_, _2625_, _2624_, _2623_, _2622_, _2621_, _2620_, _2619_, _2618_, _2617_, _2616_, _2615_, _2614_, _2613_, _2612_, _2611_, _2610_, _2609_, _2608_, _2607_, _2606_, _2605_, _2604_, _2603_, _2602_, _2601_, _2600_, _2599_, _2598_, _2597_, _2596_, _2595_, _2594_, _2593_, _2592_, _2591_, _2590_, _2589_, _2588_, _2587_, _2586_, _2585_, _2584_, _2583_, _2582_, _2581_, _2580_, _2579_, _2578_, _2577_, _2576_, _2575_, _2574_, _2573_, _2572_, _2571_, _2570_, _2569_, _2568_, _2567_, _2566_, _2565_, _2564_, _2563_, _2562_, _2561_, _2560_, _2559_, _2558_, _2557_, _2556_, _2555_, _2554_, _2553_, _2552_, _2551_, _2550_, _2549_, _2548_, _2547_, _2546_, _2545_, _2544_, _2543_, _2542_, _2541_, _2540_, _2539_, _2538_, _2537_, _2536_, _2535_, _2534_, _2533_, _2532_, _2531_, _2530_, _2529_, _2528_, _2527_, _2526_, _2525_, _0406_ });
  assign _2523_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8248|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 9'b100000000;
  assign _2524_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8244|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 8'b11111111;
  assign _2525_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8240|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 8'b11111110;
  assign _2526_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8236|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 8'b11111101;
  assign _2527_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8232|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 8'b11111100;
  assign _2528_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8228|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 8'b11111011;
  assign _2529_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8224|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 8'b11111010;
  assign _2530_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8220|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 8'b11111001;
  assign _2531_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8216|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 8'b11111000;
  assign _2532_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8212|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 8'b11110111;
  assign _2533_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8208|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 8'b11110110;
  assign _2534_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8204|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 8'b11110101;
  assign _2535_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8200|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 8'b11110100;
  assign _2536_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8196|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 8'b11110011;
  assign _2537_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8192|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 8'b11110010;
  assign _2538_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8188|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 8'b11110001;
  assign _2539_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8184|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 8'b11110000;
  assign _2540_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8180|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 8'b11101111;
  assign _2541_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8176|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 8'b11101110;
  assign _2542_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8172|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 8'b11101101;
  assign _2543_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8168|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 8'b11101100;
  assign _2544_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8164|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 8'b11101011;
  assign _2545_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8160|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 8'b11101010;
  assign _2546_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8156|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 8'b11101001;
  assign _2547_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8152|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 8'b11101000;
  assign _2548_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8148|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 8'b11100111;
  assign _2549_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8144|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 8'b11100110;
  assign _2550_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8140|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 8'b11100101;
  assign _2551_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8136|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 8'b11100100;
  assign _2552_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8132|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 8'b11100011;
  assign _2553_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8128|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 8'b11100010;
  assign _2554_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8124|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 8'b11100001;
  assign _2555_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8120|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 8'b11100000;
  assign _2556_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8116|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 8'b11011111;
  assign _2557_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8112|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 8'b11011110;
  assign _2558_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8108|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 8'b11011101;
  assign _2559_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8104|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 8'b11011100;
  assign _2560_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8100|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 8'b11011011;
  assign _2561_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8096|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 8'b11011010;
  assign _2562_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8092|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 8'b11011001;
  assign _2563_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8088|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 8'b11011000;
  assign _2564_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8084|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 8'b11010111;
  assign _2565_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8080|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 8'b11010110;
  assign _2566_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8076|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 8'b11010101;
  assign _2567_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8072|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 8'b11010100;
  assign _2568_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8068|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 8'b11010011;
  assign _2569_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8064|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 8'b11010010;
  assign _2570_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8060|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 8'b11010001;
  assign _2571_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8056|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 8'b11010000;
  assign _2572_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8052|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 8'b11001111;
  assign _2573_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8048|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 8'b11001110;
  assign _2574_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8044|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 8'b11001101;
  assign _2575_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8040|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 8'b11001100;
  assign _2576_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8036|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 8'b11001011;
  assign _2577_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8032|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 8'b11001010;
  assign _2578_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8028|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 8'b11001001;
  assign _2579_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8024|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 8'b11001000;
  assign _2580_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8020|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 8'b11000111;
  assign _2581_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8016|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 8'b11000110;
  assign _2582_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8012|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 8'b11000101;
  assign _2583_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8008|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 8'b11000100;
  assign _2584_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8004|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 8'b11000011;
  assign _2585_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8000|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 8'b11000010;
  assign _2586_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7996|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 8'b11000001;
  assign _2587_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7992|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 8'b11000000;
  assign _2588_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7988|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 8'b10111111;
  assign _2589_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7984|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 8'b10111110;
  assign _2590_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7980|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 8'b10111101;
  assign _2591_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7976|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 8'b10111100;
  assign _2592_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7972|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 8'b10111011;
  assign _2593_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7968|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 8'b10111010;
  assign _2594_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7964|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 8'b10111001;
  assign _2595_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7960|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 8'b10111000;
  assign _2596_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7956|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 8'b10110111;
  assign _2597_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7952|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 8'b10110110;
  assign _2598_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7948|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 8'b10110101;
  assign _2599_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7944|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 8'b10110100;
  assign _2600_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7940|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 8'b10110011;
  assign _2601_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7936|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 8'b10110010;
  assign _2602_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7932|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 8'b10110001;
  assign _2603_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7928|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 8'b10110000;
  assign _2604_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7924|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 8'b10101111;
  assign _2605_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7920|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 8'b10101110;
  assign _2606_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7916|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 8'b10101101;
  assign _2607_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7912|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 8'b10101100;
  assign _2608_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7908|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 8'b10101011;
  assign _2609_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7904|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 8'b10101010;
  assign _2610_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7900|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 8'b10101001;
  assign _2611_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7896|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 8'b10101000;
  assign _2612_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7892|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 8'b10100111;
  assign _2613_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7888|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 8'b10100110;
  assign _2614_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7884|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 8'b10100101;
  assign _2615_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7880|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 8'b10100100;
  assign _2616_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7876|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 8'b10100011;
  assign _2617_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7872|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 8'b10100010;
  assign _2618_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7868|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 8'b10100001;
  assign _2619_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7864|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 8'b10100000;
  assign _2620_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7860|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 8'b10011111;
  assign _2621_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7856|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 8'b10011110;
  assign _2622_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7852|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 8'b10011101;
  assign _2623_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7848|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 8'b10011100;
  assign _2624_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7844|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 8'b10011011;
  assign _2625_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7840|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 8'b10011010;
  assign _2626_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7836|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 8'b10011001;
  assign _2627_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7832|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 8'b10011000;
  assign _2628_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7828|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 8'b10010111;
  assign _2629_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7824|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 8'b10010110;
  assign _2630_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7820|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 8'b10010101;
  assign _2631_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7816|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 8'b10010100;
  assign _2632_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7812|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 8'b10010011;
  assign _2633_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7808|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 8'b10010010;
  assign _2634_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7804|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 8'b10010001;
  assign _2635_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7800|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 8'b10010000;
  assign _2636_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7796|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 8'b10001111;
  assign _2637_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7792|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 8'b10001110;
  assign _2638_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7788|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 8'b10001101;
  assign _2639_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7784|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 8'b10001100;
  assign _2640_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7780|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 8'b10001011;
  assign _2641_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7776|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 8'b10001010;
  assign _2642_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7772|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 8'b10001001;
  assign _2643_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7768|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 8'b10001000;
  assign _2644_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7764|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 8'b10000111;
  assign _2645_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7760|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 8'b10000110;
  assign _2646_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7756|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 8'b10000101;
  assign _2647_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7752|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 8'b10000100;
  assign _2648_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7748|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 8'b10000011;
  assign _2649_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7744|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 8'b10000010;
  assign _2650_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7740|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 8'b10000001;
  assign _2651_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7736|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 8'b10000000;
  assign _2652_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7732|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 7'b1111111;
  assign _2653_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7728|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 7'b1111110;
  assign _2654_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7724|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 7'b1111101;
  assign _2655_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7720|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 7'b1111100;
  assign _2656_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7716|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 7'b1111011;
  assign _2657_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7712|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 7'b1111010;
  assign _2658_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7708|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 7'b1111001;
  assign _2659_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7704|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 7'b1111000;
  assign _2660_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7700|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 7'b1110111;
  assign _2661_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7696|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 7'b1110110;
  assign _2662_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7692|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 7'b1110101;
  assign _2663_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7688|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 7'b1110100;
  assign _2664_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7684|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 7'b1110011;
  assign _2665_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7680|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 7'b1110010;
  assign _2666_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7676|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 7'b1110001;
  assign _2667_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7672|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 7'b1110000;
  assign _2668_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7668|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 7'b1101111;
  assign _2669_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7664|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 7'b1101110;
  assign _2670_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7660|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 7'b1101101;
  assign _2671_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7656|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 7'b1101100;
  assign _2672_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7652|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 7'b1101011;
  assign _2673_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7648|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 7'b1101010;
  assign _2674_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7644|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 7'b1101001;
  assign _2675_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7640|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 7'b1101000;
  assign _2676_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7636|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 7'b1100111;
  assign _2677_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7632|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 7'b1100110;
  assign _2678_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7628|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 7'b1100101;
  assign _2679_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7624|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 7'b1100100;
  assign _2680_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7620|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 7'b1100011;
  assign _2681_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7616|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 7'b1100010;
  assign _2682_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7612|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 7'b1100001;
  assign _2683_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7608|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 7'b1100000;
  assign _2684_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7604|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 7'b1011111;
  assign _2685_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7600|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 7'b1011110;
  assign _2686_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7596|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 7'b1011101;
  assign _2687_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7592|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 7'b1011100;
  assign _2688_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7588|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 7'b1011011;
  assign _2689_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7584|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 7'b1011010;
  assign _2690_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7580|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 7'b1011001;
  assign _2691_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7576|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 7'b1011000;
  assign _2692_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7572|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 7'b1010111;
  assign _2693_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7568|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 7'b1010110;
  assign _2694_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7564|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 7'b1010101;
  assign _2695_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7560|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 7'b1010100;
  assign _2696_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7556|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 7'b1010011;
  assign _2697_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7552|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 7'b1010010;
  assign _2698_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7548|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 7'b1010001;
  assign _2699_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7544|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 7'b1010000;
  assign _2700_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7540|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 7'b1001111;
  assign _2701_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7536|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 7'b1001110;
  assign _2702_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7532|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 7'b1001101;
  assign _2703_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7528|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 7'b1001100;
  assign _2704_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7524|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 7'b1001011;
  assign _2705_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7520|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 7'b1001010;
  assign _2706_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7516|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 7'b1001001;
  assign _2707_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7512|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 7'b1001000;
  assign _2708_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7508|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 7'b1000111;
  assign _2709_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7504|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 7'b1000110;
  assign _2710_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7500|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 7'b1000101;
  assign _2711_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7496|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 7'b1000100;
  assign _2712_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7492|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 7'b1000011;
  assign _2713_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7488|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 7'b1000010;
  assign _2714_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7484|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 7'b1000001;
  assign _2715_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7480|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 7'b1000000;
  assign _2716_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7476|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 6'b111111;
  assign _2717_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7472|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 6'b111110;
  assign _2718_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7468|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 6'b111101;
  assign _2719_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7464|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 6'b111100;
  assign _2720_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7460|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 6'b111011;
  assign _2721_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7456|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 6'b111010;
  assign _2722_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7452|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 6'b111001;
  assign _2723_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7448|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 6'b111000;
  assign _2724_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7444|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 6'b110111;
  assign _2725_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7440|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 6'b110110;
  assign _2726_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7436|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 6'b110101;
  assign _2727_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7432|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 6'b110100;
  assign _2728_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7428|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 6'b110011;
  assign _2729_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7424|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 6'b110010;
  assign _2730_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7420|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 6'b110001;
  assign _2731_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7416|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 6'b110000;
  assign _2732_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7412|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 6'b101111;
  assign _2733_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7408|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 6'b101110;
  assign _2734_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7404|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 6'b101101;
  assign _2735_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7400|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 6'b101100;
  assign _2736_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7396|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 6'b101011;
  assign _2737_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7392|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 6'b101010;
  assign _2738_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7388|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 6'b101001;
  assign _2739_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7384|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 6'b101000;
  assign _2740_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7380|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 6'b100111;
  assign _2741_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7376|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 6'b100110;
  assign _2742_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7372|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 6'b100101;
  assign _2743_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7368|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 6'b100100;
  assign _2744_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7364|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 6'b100011;
  assign _2745_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7360|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 6'b100010;
  assign _2746_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7356|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 6'b100001;
  assign _2747_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7352|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 6'b100000;
  assign _2748_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7348|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 5'b11111;
  assign _2749_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7344|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 5'b11110;
  assign _2750_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7340|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 5'b11101;
  assign _2751_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7336|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 5'b11100;
  assign _2752_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7332|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 5'b11011;
  assign _2753_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7328|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 5'b11010;
  assign _2754_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7324|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 5'b11001;
  assign _2755_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7320|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 5'b11000;
  assign _2756_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7316|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 5'b10111;
  assign _2757_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7312|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 5'b10110;
  assign _2758_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7308|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 5'b10101;
  assign _2759_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7304|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 5'b10100;
  assign _2760_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7300|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 5'b10011;
  assign _2761_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7296|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 5'b10010;
  assign _2762_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7292|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 5'b10001;
  assign _2763_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7288|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 5'b10000;
  assign _2764_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7284|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 4'b1111;
  assign _2765_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7280|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 4'b1110;
  assign _2766_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7276|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 4'b1101;
  assign _2767_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7272|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 4'b1100;
  assign _2768_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7268|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 4'b1011;
  assign _2769_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7264|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 4'b1010;
  assign _2770_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7260|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 4'b1001;
  assign _2771_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7256|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 4'b1000;
  assign _2772_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7252|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 3'b111;
  assign _2773_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7248|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 3'b110;
  assign _2774_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7244|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 3'b101;
  assign _2775_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7240|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 3'b100;
  assign _2776_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7236|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 2'b11;
  assign _2777_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7232|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 2'b10;
  assign _2778_ = dp2lut_Y_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7228|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) 1'b1;
  assign _2779_ = ! (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7224|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *) dp2lut_Y_entry_0;
  assign _2780_ = dp2lut_Yinfo_0[17] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7219" *) density_reg256 : _2522_;
  assign _2781_ = dp2lut_Yinfo_0[16] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7216" *) density_reg0 : _2780_;
  assign _0286_ = _0400_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7215" *) _2781_ : lut_Y_data_01;
  function [15:0] _6640_;
    input [15:0] a;
    input [4095:0] b;
    input [255:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:8248|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7223" *)
    (* parallel_case *)
    casez (s)
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1:
        _6640_ = b[15:0];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?:
        _6640_ = b[31:16];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??:
        _6640_ = b[47:32];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???:
        _6640_ = b[63:48];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????:
        _6640_ = b[79:64];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????:
        _6640_ = b[95:80];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????:
        _6640_ = b[111:96];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????:
        _6640_ = b[127:112];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????:
        _6640_ = b[143:128];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????:
        _6640_ = b[159:144];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????:
        _6640_ = b[175:160];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????:
        _6640_ = b[191:176];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????:
        _6640_ = b[207:192];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????:
        _6640_ = b[223:208];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????:
        _6640_ = b[239:224];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????:
        _6640_ = b[255:240];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????:
        _6640_ = b[271:256];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????:
        _6640_ = b[287:272];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????:
        _6640_ = b[303:288];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????:
        _6640_ = b[319:304];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????:
        _6640_ = b[335:320];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????:
        _6640_ = b[351:336];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????:
        _6640_ = b[367:352];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????:
        _6640_ = b[383:368];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????:
        _6640_ = b[399:384];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????:
        _6640_ = b[415:400];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????:
        _6640_ = b[431:416];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????:
        _6640_ = b[447:432];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????:
        _6640_ = b[463:448];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????:
        _6640_ = b[479:464];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????:
        _6640_ = b[495:480];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????:
        _6640_ = b[511:496];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????:
        _6640_ = b[527:512];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????:
        _6640_ = b[543:528];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????:
        _6640_ = b[559:544];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????:
        _6640_ = b[575:560];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????:
        _6640_ = b[591:576];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????:
        _6640_ = b[607:592];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????:
        _6640_ = b[623:608];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????:
        _6640_ = b[639:624];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????:
        _6640_ = b[655:640];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????:
        _6640_ = b[671:656];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????:
        _6640_ = b[687:672];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????:
        _6640_ = b[703:688];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????:
        _6640_ = b[719:704];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????:
        _6640_ = b[735:720];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????:
        _6640_ = b[751:736];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????:
        _6640_ = b[767:752];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????:
        _6640_ = b[783:768];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????:
        _6640_ = b[799:784];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????:
        _6640_ = b[815:800];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????:
        _6640_ = b[831:816];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????:
        _6640_ = b[847:832];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????:
        _6640_ = b[863:848];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????:
        _6640_ = b[879:864];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????:
        _6640_ = b[895:880];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????:
        _6640_ = b[911:896];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????:
        _6640_ = b[927:912];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????:
        _6640_ = b[943:928];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????:
        _6640_ = b[959:944];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????:
        _6640_ = b[975:960];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????:
        _6640_ = b[991:976];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????:
        _6640_ = b[1007:992];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????:
        _6640_ = b[1023:1008];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????:
        _6640_ = b[1039:1024];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????:
        _6640_ = b[1055:1040];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????:
        _6640_ = b[1071:1056];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????:
        _6640_ = b[1087:1072];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????:
        _6640_ = b[1103:1088];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????:
        _6640_ = b[1119:1104];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????:
        _6640_ = b[1135:1120];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????:
        _6640_ = b[1151:1136];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????:
        _6640_ = b[1167:1152];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????:
        _6640_ = b[1183:1168];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????:
        _6640_ = b[1199:1184];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????:
        _6640_ = b[1215:1200];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????:
        _6640_ = b[1231:1216];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????:
        _6640_ = b[1247:1232];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????:
        _6640_ = b[1263:1248];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????:
        _6640_ = b[1279:1264];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????:
        _6640_ = b[1295:1280];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????:
        _6640_ = b[1311:1296];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????:
        _6640_ = b[1327:1312];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????:
        _6640_ = b[1343:1328];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????:
        _6640_ = b[1359:1344];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????:
        _6640_ = b[1375:1360];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????:
        _6640_ = b[1391:1376];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????:
        _6640_ = b[1407:1392];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????:
        _6640_ = b[1423:1408];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????:
        _6640_ = b[1439:1424];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????:
        _6640_ = b[1455:1440];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????:
        _6640_ = b[1471:1456];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????:
        _6640_ = b[1487:1472];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????:
        _6640_ = b[1503:1488];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????:
        _6640_ = b[1519:1504];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????:
        _6640_ = b[1535:1520];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????:
        _6640_ = b[1551:1536];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????:
        _6640_ = b[1567:1552];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????:
        _6640_ = b[1583:1568];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????:
        _6640_ = b[1599:1584];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6640_ = b[1615:1600];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6640_ = b[1631:1616];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6640_ = b[1647:1632];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6640_ = b[1663:1648];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6640_ = b[1679:1664];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6640_ = b[1695:1680];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6640_ = b[1711:1696];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6640_ = b[1727:1712];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6640_ = b[1743:1728];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6640_ = b[1759:1744];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6640_ = b[1775:1760];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6640_ = b[1791:1776];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6640_ = b[1807:1792];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6640_ = b[1823:1808];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6640_ = b[1839:1824];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6640_ = b[1855:1840];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6640_ = b[1871:1856];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6640_ = b[1887:1872];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6640_ = b[1903:1888];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6640_ = b[1919:1904];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6640_ = b[1935:1920];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6640_ = b[1951:1936];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6640_ = b[1967:1952];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6640_ = b[1983:1968];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6640_ = b[1999:1984];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6640_ = b[2015:2000];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6640_ = b[2031:2016];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6640_ = b[2047:2032];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6640_ = b[2063:2048];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6640_ = b[2079:2064];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6640_ = b[2095:2080];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6640_ = b[2111:2096];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6640_ = b[2127:2112];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6640_ = b[2143:2128];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6640_ = b[2159:2144];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6640_ = b[2175:2160];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6640_ = b[2191:2176];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6640_ = b[2207:2192];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6640_ = b[2223:2208];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6640_ = b[2239:2224];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6640_ = b[2255:2240];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6640_ = b[2271:2256];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6640_ = b[2287:2272];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6640_ = b[2303:2288];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6640_ = b[2319:2304];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6640_ = b[2335:2320];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6640_ = b[2351:2336];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6640_ = b[2367:2352];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6640_ = b[2383:2368];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6640_ = b[2399:2384];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6640_ = b[2415:2400];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6640_ = b[2431:2416];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6640_ = b[2447:2432];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6640_ = b[2463:2448];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6640_ = b[2479:2464];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6640_ = b[2495:2480];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6640_ = b[2511:2496];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6640_ = b[2527:2512];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6640_ = b[2543:2528];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6640_ = b[2559:2544];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6640_ = b[2575:2560];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6640_ = b[2591:2576];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6640_ = b[2607:2592];
      256'b????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6640_ = b[2623:2608];
      256'b???????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6640_ = b[2639:2624];
      256'b??????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6640_ = b[2655:2640];
      256'b?????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6640_ = b[2671:2656];
      256'b????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6640_ = b[2687:2672];
      256'b???????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6640_ = b[2703:2688];
      256'b??????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6640_ = b[2719:2704];
      256'b?????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6640_ = b[2735:2720];
      256'b????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6640_ = b[2751:2736];
      256'b???????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6640_ = b[2767:2752];
      256'b??????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6640_ = b[2783:2768];
      256'b?????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6640_ = b[2799:2784];
      256'b????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6640_ = b[2815:2800];
      256'b???????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6640_ = b[2831:2816];
      256'b??????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6640_ = b[2847:2832];
      256'b?????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6640_ = b[2863:2848];
      256'b????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6640_ = b[2879:2864];
      256'b???????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6640_ = b[2895:2880];
      256'b??????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6640_ = b[2911:2896];
      256'b?????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6640_ = b[2927:2912];
      256'b????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6640_ = b[2943:2928];
      256'b???????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6640_ = b[2959:2944];
      256'b??????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6640_ = b[2975:2960];
      256'b?????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6640_ = b[2991:2976];
      256'b????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6640_ = b[3007:2992];
      256'b???????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6640_ = b[3023:3008];
      256'b??????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6640_ = b[3039:3024];
      256'b?????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6640_ = b[3055:3040];
      256'b????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6640_ = b[3071:3056];
      256'b???????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6640_ = b[3087:3072];
      256'b??????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6640_ = b[3103:3088];
      256'b?????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6640_ = b[3119:3104];
      256'b????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6640_ = b[3135:3120];
      256'b???????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6640_ = b[3151:3136];
      256'b??????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6640_ = b[3167:3152];
      256'b?????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6640_ = b[3183:3168];
      256'b????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6640_ = b[3199:3184];
      256'b???????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6640_ = b[3215:3200];
      256'b??????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6640_ = b[3231:3216];
      256'b?????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6640_ = b[3247:3232];
      256'b????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6640_ = b[3263:3248];
      256'b???????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6640_ = b[3279:3264];
      256'b??????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6640_ = b[3295:3280];
      256'b?????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6640_ = b[3311:3296];
      256'b????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6640_ = b[3327:3312];
      256'b???????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6640_ = b[3343:3328];
      256'b??????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6640_ = b[3359:3344];
      256'b?????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6640_ = b[3375:3360];
      256'b????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6640_ = b[3391:3376];
      256'b???????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6640_ = b[3407:3392];
      256'b??????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6640_ = b[3423:3408];
      256'b?????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6640_ = b[3439:3424];
      256'b????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6640_ = b[3455:3440];
      256'b???????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6640_ = b[3471:3456];
      256'b??????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6640_ = b[3487:3472];
      256'b?????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6640_ = b[3503:3488];
      256'b????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6640_ = b[3519:3504];
      256'b???????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6640_ = b[3535:3520];
      256'b??????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6640_ = b[3551:3536];
      256'b?????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6640_ = b[3567:3552];
      256'b????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6640_ = b[3583:3568];
      256'b???????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6640_ = b[3599:3584];
      256'b??????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6640_ = b[3615:3600];
      256'b?????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6640_ = b[3631:3616];
      256'b????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6640_ = b[3647:3632];
      256'b???????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6640_ = b[3663:3648];
      256'b??????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6640_ = b[3679:3664];
      256'b?????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6640_ = b[3695:3680];
      256'b????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6640_ = b[3711:3696];
      256'b???????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6640_ = b[3727:3712];
      256'b??????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6640_ = b[3743:3728];
      256'b?????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6640_ = b[3759:3744];
      256'b????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6640_ = b[3775:3760];
      256'b???????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6640_ = b[3791:3776];
      256'b??????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6640_ = b[3807:3792];
      256'b?????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6640_ = b[3823:3808];
      256'b????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6640_ = b[3839:3824];
      256'b???????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6640_ = b[3855:3840];
      256'b??????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6640_ = b[3871:3856];
      256'b?????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6640_ = b[3887:3872];
      256'b????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6640_ = b[3903:3888];
      256'b???????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6640_ = b[3919:3904];
      256'b??????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6640_ = b[3935:3920];
      256'b?????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6640_ = b[3951:3936];
      256'b????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6640_ = b[3967:3952];
      256'b???????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6640_ = b[3983:3968];
      256'b??????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6640_ = b[3999:3984];
      256'b?????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6640_ = b[4015:4000];
      256'b????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6640_ = b[4031:4016];
      256'b???1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6640_ = b[4047:4032];
      256'b??1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6640_ = b[4063:4048];
      256'b?1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6640_ = b[4079:4064];
      256'b1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _6640_ = b[4095:4080];
      default:
        _6640_ = a;
    endcase
  endfunction
  assign _2782_ = _6640_(density_reg0, { density_reg1, density_reg2, density_reg3, density_reg4, density_reg5, density_reg6, density_reg7, density_reg8, density_reg9, density_reg10, density_reg11, density_reg12, density_reg13, density_reg14, density_reg15, density_reg16, density_reg17, density_reg18, density_reg19, density_reg20, density_reg21, density_reg22, density_reg23, density_reg24, density_reg25, density_reg26, density_reg27, density_reg28, density_reg29, density_reg30, density_reg31, density_reg32, density_reg33, density_reg34, density_reg35, density_reg36, density_reg37, density_reg38, density_reg39, density_reg40, density_reg41, density_reg42, density_reg43, density_reg44, density_reg45, density_reg46, density_reg47, density_reg48, density_reg49, density_reg50, density_reg51, density_reg52, density_reg53, density_reg54, density_reg55, density_reg56, density_reg57, density_reg58, density_reg59, density_reg60, density_reg61, density_reg62, density_reg63, density_reg64, density_reg65, density_reg66, density_reg67, density_reg68, density_reg69, density_reg70, density_reg71, density_reg72, density_reg73, density_reg74, density_reg75, density_reg76, density_reg77, density_reg78, density_reg79, density_reg80, density_reg81, density_reg82, density_reg83, density_reg84, density_reg85, density_reg86, density_reg87, density_reg88, density_reg89, density_reg90, density_reg91, density_reg92, density_reg93, density_reg94, density_reg95, density_reg96, density_reg97, density_reg98, density_reg99, density_reg100, density_reg101, density_reg102, density_reg103, density_reg104, density_reg105, density_reg106, density_reg107, density_reg108, density_reg109, density_reg110, density_reg111, density_reg112, density_reg113, density_reg114, density_reg115, density_reg116, density_reg117, density_reg118, density_reg119, density_reg120, density_reg121, density_reg122, density_reg123, density_reg124, density_reg125, density_reg126, density_reg127, density_reg128, density_reg129, density_reg130, density_reg131, density_reg132, density_reg133, density_reg134, density_reg135, density_reg136, density_reg137, density_reg138, density_reg139, density_reg140, density_reg141, density_reg142, density_reg143, density_reg144, density_reg145, density_reg146, density_reg147, density_reg148, density_reg149, density_reg150, density_reg151, density_reg152, density_reg153, density_reg154, density_reg155, density_reg156, density_reg157, density_reg158, density_reg159, density_reg160, density_reg161, density_reg162, density_reg163, density_reg164, density_reg165, density_reg166, density_reg167, density_reg168, density_reg169, density_reg170, density_reg171, density_reg172, density_reg173, density_reg174, density_reg175, density_reg176, density_reg177, density_reg178, density_reg179, density_reg180, density_reg181, density_reg182, density_reg183, density_reg184, density_reg185, density_reg186, density_reg187, density_reg188, density_reg189, density_reg190, density_reg191, density_reg192, density_reg193, density_reg194, density_reg195, density_reg196, density_reg197, density_reg198, density_reg199, density_reg200, density_reg201, density_reg202, density_reg203, density_reg204, density_reg205, density_reg206, density_reg207, density_reg208, density_reg209, density_reg210, density_reg211, density_reg212, density_reg213, density_reg214, density_reg215, density_reg216, density_reg217, density_reg218, density_reg219, density_reg220, density_reg221, density_reg222, density_reg223, density_reg224, density_reg225, density_reg226, density_reg227, density_reg228, density_reg229, density_reg230, density_reg231, density_reg232, density_reg233, density_reg234, density_reg235, density_reg236, density_reg237, density_reg238, density_reg239, density_reg240, density_reg241, density_reg242, density_reg243, density_reg244, density_reg245, density_reg246, density_reg247, density_reg248, density_reg249, density_reg250, density_reg251, density_reg252, density_reg253, density_reg254, density_reg255, density_reg256 }, { _2778_, _2777_, _2776_, _2775_, _2774_, _2773_, _2772_, _2771_, _2770_, _2769_, _2768_, _2767_, _2766_, _2765_, _2764_, _2763_, _2762_, _2761_, _2760_, _2759_, _2758_, _2757_, _2756_, _2755_, _2754_, _2753_, _2752_, _2751_, _2750_, _2749_, _2748_, _2747_, _2746_, _2745_, _2744_, _2743_, _2742_, _2741_, _2740_, _2739_, _2738_, _2737_, _2736_, _2735_, _2734_, _2733_, _2732_, _2731_, _2730_, _2729_, _2728_, _2727_, _2726_, _2725_, _2724_, _2723_, _2722_, _2721_, _2720_, _2719_, _2718_, _2717_, _2716_, _2715_, _2714_, _2713_, _2712_, _2711_, _2710_, _2709_, _2708_, _2707_, _2706_, _2705_, _2704_, _2703_, _2702_, _2701_, _2700_, _2699_, _2698_, _2697_, _2696_, _2695_, _2694_, _2693_, _2692_, _2691_, _2690_, _2689_, _2688_, _2687_, _2686_, _2685_, _2684_, _2683_, _2682_, _2681_, _2680_, _2679_, _2678_, _2677_, _2676_, _2675_, _2674_, _2673_, _2672_, _2671_, _2670_, _2669_, _2668_, _2667_, _2666_, _2665_, _2664_, _2663_, _2662_, _2661_, _2660_, _2659_, _2658_, _2657_, _2656_, _2655_, _2654_, _2653_, _2652_, _2651_, _2650_, _2649_, _2648_, _2647_, _2646_, _2645_, _2644_, _2643_, _2642_, _2641_, _2640_, _2639_, _2638_, _2637_, _2636_, _2635_, _2634_, _2633_, _2632_, _2631_, _2630_, _2629_, _2628_, _2627_, _2626_, _2625_, _2624_, _2623_, _2622_, _2621_, _2620_, _2619_, _2618_, _2617_, _2616_, _2615_, _2614_, _2613_, _2612_, _2611_, _2610_, _2609_, _2608_, _2607_, _2606_, _2605_, _2604_, _2603_, _2602_, _2601_, _2600_, _2599_, _2598_, _2597_, _2596_, _2595_, _2594_, _2593_, _2592_, _2591_, _2590_, _2589_, _2588_, _2587_, _2586_, _2585_, _2584_, _2583_, _2582_, _2581_, _2580_, _2579_, _2578_, _2577_, _2576_, _2575_, _2574_, _2573_, _2572_, _2571_, _2570_, _2569_, _2568_, _2567_, _2566_, _2565_, _2564_, _2563_, _2562_, _2561_, _2560_, _2559_, _2558_, _2557_, _2556_, _2555_, _2554_, _2553_, _2552_, _2551_, _2550_, _2549_, _2548_, _2547_, _2546_, _2545_, _2544_, _2543_, _2542_, _2541_, _2540_, _2539_, _2538_, _2537_, _2536_, _2535_, _2534_, _2533_, _2532_, _2531_, _2530_, _2529_, _2528_, _2527_, _2526_, _2525_, _2524_, _2523_ });
  assign _2783_ = dp2lut_Yinfo_0[17] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7219" *) density_reg256 : _2782_;
  assign _2784_ = dp2lut_Yinfo_0[16] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7216" *) density_reg0 : _2783_;
  assign _0285_ = _0400_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7215" *) _2784_ : lut_Y_data_00;
  function [15:0] _6644_;
    input [15:0] a;
    input [1023:0] b;
    input [63:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7196|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6939" *)
    (* parallel_case *)
    casez (s)
      64'b???????????????????????????????????????????????????????????????1:
        _6644_ = b[15:0];
      64'b??????????????????????????????????????????????????????????????1?:
        _6644_ = b[31:16];
      64'b?????????????????????????????????????????????????????????????1??:
        _6644_ = b[47:32];
      64'b????????????????????????????????????????????????????????????1???:
        _6644_ = b[63:48];
      64'b???????????????????????????????????????????????????????????1????:
        _6644_ = b[79:64];
      64'b??????????????????????????????????????????????????????????1?????:
        _6644_ = b[95:80];
      64'b?????????????????????????????????????????????????????????1??????:
        _6644_ = b[111:96];
      64'b????????????????????????????????????????????????????????1???????:
        _6644_ = b[127:112];
      64'b???????????????????????????????????????????????????????1????????:
        _6644_ = b[143:128];
      64'b??????????????????????????????????????????????????????1?????????:
        _6644_ = b[159:144];
      64'b?????????????????????????????????????????????????????1??????????:
        _6644_ = b[175:160];
      64'b????????????????????????????????????????????????????1???????????:
        _6644_ = b[191:176];
      64'b???????????????????????????????????????????????????1????????????:
        _6644_ = b[207:192];
      64'b??????????????????????????????????????????????????1?????????????:
        _6644_ = b[223:208];
      64'b?????????????????????????????????????????????????1??????????????:
        _6644_ = b[239:224];
      64'b????????????????????????????????????????????????1???????????????:
        _6644_ = b[255:240];
      64'b???????????????????????????????????????????????1????????????????:
        _6644_ = b[271:256];
      64'b??????????????????????????????????????????????1?????????????????:
        _6644_ = b[287:272];
      64'b?????????????????????????????????????????????1??????????????????:
        _6644_ = b[303:288];
      64'b????????????????????????????????????????????1???????????????????:
        _6644_ = b[319:304];
      64'b???????????????????????????????????????????1????????????????????:
        _6644_ = b[335:320];
      64'b??????????????????????????????????????????1?????????????????????:
        _6644_ = b[351:336];
      64'b?????????????????????????????????????????1??????????????????????:
        _6644_ = b[367:352];
      64'b????????????????????????????????????????1???????????????????????:
        _6644_ = b[383:368];
      64'b???????????????????????????????????????1????????????????????????:
        _6644_ = b[399:384];
      64'b??????????????????????????????????????1?????????????????????????:
        _6644_ = b[415:400];
      64'b?????????????????????????????????????1??????????????????????????:
        _6644_ = b[431:416];
      64'b????????????????????????????????????1???????????????????????????:
        _6644_ = b[447:432];
      64'b???????????????????????????????????1????????????????????????????:
        _6644_ = b[463:448];
      64'b??????????????????????????????????1?????????????????????????????:
        _6644_ = b[479:464];
      64'b?????????????????????????????????1??????????????????????????????:
        _6644_ = b[495:480];
      64'b????????????????????????????????1???????????????????????????????:
        _6644_ = b[511:496];
      64'b???????????????????????????????1????????????????????????????????:
        _6644_ = b[527:512];
      64'b??????????????????????????????1?????????????????????????????????:
        _6644_ = b[543:528];
      64'b?????????????????????????????1??????????????????????????????????:
        _6644_ = b[559:544];
      64'b????????????????????????????1???????????????????????????????????:
        _6644_ = b[575:560];
      64'b???????????????????????????1????????????????????????????????????:
        _6644_ = b[591:576];
      64'b??????????????????????????1?????????????????????????????????????:
        _6644_ = b[607:592];
      64'b?????????????????????????1??????????????????????????????????????:
        _6644_ = b[623:608];
      64'b????????????????????????1???????????????????????????????????????:
        _6644_ = b[639:624];
      64'b???????????????????????1????????????????????????????????????????:
        _6644_ = b[655:640];
      64'b??????????????????????1?????????????????????????????????????????:
        _6644_ = b[671:656];
      64'b?????????????????????1??????????????????????????????????????????:
        _6644_ = b[687:672];
      64'b????????????????????1???????????????????????????????????????????:
        _6644_ = b[703:688];
      64'b???????????????????1????????????????????????????????????????????:
        _6644_ = b[719:704];
      64'b??????????????????1?????????????????????????????????????????????:
        _6644_ = b[735:720];
      64'b?????????????????1??????????????????????????????????????????????:
        _6644_ = b[751:736];
      64'b????????????????1???????????????????????????????????????????????:
        _6644_ = b[767:752];
      64'b???????????????1????????????????????????????????????????????????:
        _6644_ = b[783:768];
      64'b??????????????1?????????????????????????????????????????????????:
        _6644_ = b[799:784];
      64'b?????????????1??????????????????????????????????????????????????:
        _6644_ = b[815:800];
      64'b????????????1???????????????????????????????????????????????????:
        _6644_ = b[831:816];
      64'b???????????1????????????????????????????????????????????????????:
        _6644_ = b[847:832];
      64'b??????????1?????????????????????????????????????????????????????:
        _6644_ = b[863:848];
      64'b?????????1??????????????????????????????????????????????????????:
        _6644_ = b[879:864];
      64'b????????1???????????????????????????????????????????????????????:
        _6644_ = b[895:880];
      64'b???????1????????????????????????????????????????????????????????:
        _6644_ = b[911:896];
      64'b??????1?????????????????????????????????????????????????????????:
        _6644_ = b[927:912];
      64'b?????1??????????????????????????????????????????????????????????:
        _6644_ = b[943:928];
      64'b????1???????????????????????????????????????????????????????????:
        _6644_ = b[959:944];
      64'b???1????????????????????????????????????????????????????????????:
        _6644_ = b[975:960];
      64'b??1?????????????????????????????????????????????????????????????:
        _6644_ = b[991:976];
      64'b?1??????????????????????????????????????????????????????????????:
        _6644_ = b[1007:992];
      64'b1???????????????????????????????????????????????????????????????:
        _6644_ = b[1023:1008];
      default:
        _6644_ = a;
    endcase
  endfunction
  assign _2785_ = _6644_(raw_reg0, { raw_reg1, raw_reg2, raw_reg3, raw_reg4, raw_reg5, raw_reg6, raw_reg7, raw_reg8, raw_reg9, raw_reg10, raw_reg11, raw_reg12, raw_reg13, raw_reg14, raw_reg15, raw_reg16, raw_reg17, raw_reg18, raw_reg19, raw_reg20, raw_reg21, raw_reg22, raw_reg23, raw_reg24, raw_reg25, raw_reg26, raw_reg27, raw_reg28, raw_reg29, raw_reg30, raw_reg31, raw_reg32, raw_reg33, raw_reg34, raw_reg35, raw_reg36, raw_reg37, raw_reg38, raw_reg39, raw_reg40, raw_reg41, raw_reg42, raw_reg43, raw_reg44, raw_reg45, raw_reg46, raw_reg47, raw_reg48, raw_reg49, raw_reg50, raw_reg51, raw_reg52, raw_reg53, raw_reg54, raw_reg55, raw_reg56, raw_reg57, raw_reg58, raw_reg59, raw_reg60, raw_reg61, raw_reg62, raw_reg63, raw_reg64 }, { _2850_, _2849_, _2848_, _2847_, _2846_, _2845_, _2844_, _2843_, _2842_, _2841_, _2840_, _2839_, _2838_, _2837_, _2836_, _2835_, _2834_, _2833_, _2832_, _2831_, _2830_, _2829_, _2828_, _2827_, _2826_, _2825_, _2824_, _2823_, _2822_, _2821_, _2820_, _2819_, _2818_, _2817_, _2816_, _2815_, _2814_, _2813_, _2812_, _2811_, _2810_, _2809_, _2808_, _2807_, _2806_, _2805_, _2804_, _2803_, _2802_, _2801_, _2800_, _2799_, _2798_, _2797_, _2796_, _2795_, _2794_, _2793_, _2792_, _2791_, _2790_, _2789_, _2788_, _0408_ });
  assign _2786_ = dp2lut_X_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7196|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6939" *) 7'b1000000;
  assign _2787_ = dp2lut_X_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7192|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6939" *) 6'b111111;
  assign _2788_ = dp2lut_X_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7188|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6939" *) 6'b111110;
  assign _2789_ = dp2lut_X_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7184|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6939" *) 6'b111101;
  assign _2790_ = dp2lut_X_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7180|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6939" *) 6'b111100;
  assign _2791_ = dp2lut_X_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7176|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6939" *) 6'b111011;
  assign _2792_ = dp2lut_X_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7172|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6939" *) 6'b111010;
  assign _2793_ = dp2lut_X_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7168|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6939" *) 6'b111001;
  assign _2794_ = dp2lut_X_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7164|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6939" *) 6'b111000;
  assign _2795_ = dp2lut_X_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7160|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6939" *) 6'b110111;
  assign _2796_ = dp2lut_X_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7156|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6939" *) 6'b110110;
  assign _2797_ = dp2lut_X_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7152|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6939" *) 6'b110101;
  assign _2798_ = dp2lut_X_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7148|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6939" *) 6'b110100;
  assign _2799_ = dp2lut_X_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7144|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6939" *) 6'b110011;
  assign _2800_ = dp2lut_X_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7140|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6939" *) 6'b110010;
  assign _2801_ = dp2lut_X_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7136|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6939" *) 6'b110001;
  assign _2802_ = dp2lut_X_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7132|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6939" *) 6'b110000;
  assign _2803_ = dp2lut_X_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7128|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6939" *) 6'b101111;
  assign _2804_ = dp2lut_X_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7124|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6939" *) 6'b101110;
  assign _2805_ = dp2lut_X_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7120|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6939" *) 6'b101101;
  assign _2806_ = dp2lut_X_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7116|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6939" *) 6'b101100;
  assign _2807_ = dp2lut_X_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7112|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6939" *) 6'b101011;
  assign _2808_ = dp2lut_X_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7108|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6939" *) 6'b101010;
  assign _2809_ = dp2lut_X_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7104|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6939" *) 6'b101001;
  assign _2810_ = dp2lut_X_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7100|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6939" *) 6'b101000;
  assign _2811_ = dp2lut_X_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7096|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6939" *) 6'b100111;
  assign _2812_ = dp2lut_X_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7092|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6939" *) 6'b100110;
  assign _2813_ = dp2lut_X_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7088|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6939" *) 6'b100101;
  assign _2814_ = dp2lut_X_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7084|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6939" *) 6'b100100;
  assign _2815_ = dp2lut_X_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7080|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6939" *) 6'b100011;
  assign _2816_ = dp2lut_X_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7076|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6939" *) 6'b100010;
  assign _2817_ = dp2lut_X_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7072|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6939" *) 6'b100001;
  assign _2818_ = dp2lut_X_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7068|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6939" *) 6'b100000;
  assign _2819_ = dp2lut_X_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7064|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6939" *) 5'b11111;
  assign _2820_ = dp2lut_X_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7060|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6939" *) 5'b11110;
  assign _2821_ = dp2lut_X_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7056|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6939" *) 5'b11101;
  assign _2822_ = dp2lut_X_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7052|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6939" *) 5'b11100;
  assign _2823_ = dp2lut_X_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7048|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6939" *) 5'b11011;
  assign _2824_ = dp2lut_X_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7044|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6939" *) 5'b11010;
  assign _2825_ = dp2lut_X_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7040|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6939" *) 5'b11001;
  assign _2826_ = dp2lut_X_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7036|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6939" *) 5'b11000;
  assign _2827_ = dp2lut_X_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7032|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6939" *) 5'b10111;
  assign _2828_ = dp2lut_X_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7028|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6939" *) 5'b10110;
  assign _2829_ = dp2lut_X_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7024|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6939" *) 5'b10101;
  assign _2830_ = dp2lut_X_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7020|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6939" *) 5'b10100;
  assign _2831_ = dp2lut_X_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7016|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6939" *) 5'b10011;
  assign _2832_ = dp2lut_X_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7012|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6939" *) 5'b10010;
  assign _2833_ = dp2lut_X_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7008|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6939" *) 5'b10001;
  assign _2834_ = dp2lut_X_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7004|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6939" *) 5'b10000;
  assign _2835_ = dp2lut_X_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7000|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6939" *) 4'b1111;
  assign _2836_ = dp2lut_X_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6996|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6939" *) 4'b1110;
  assign _2837_ = dp2lut_X_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6992|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6939" *) 4'b1101;
  assign _2838_ = dp2lut_X_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6988|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6939" *) 4'b1100;
  assign _2839_ = dp2lut_X_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6984|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6939" *) 4'b1011;
  assign _2840_ = dp2lut_X_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6980|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6939" *) 4'b1010;
  assign _2841_ = dp2lut_X_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6976|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6939" *) 4'b1001;
  assign _2842_ = dp2lut_X_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6972|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6939" *) 4'b1000;
  assign _2843_ = dp2lut_X_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6968|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6939" *) 3'b111;
  assign _2844_ = dp2lut_X_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6964|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6939" *) 3'b110;
  assign _2845_ = dp2lut_X_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6960|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6939" *) 3'b101;
  assign _2846_ = dp2lut_X_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6956|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6939" *) 3'b100;
  assign _2847_ = dp2lut_X_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6952|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6939" *) 2'b11;
  assign _2848_ = dp2lut_X_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6948|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6939" *) 2'b10;
  assign _2849_ = dp2lut_X_entry_7 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6944|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6939" *) 1'b1;
  assign _2850_ = ! (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6940|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6939" *) dp2lut_X_entry_7;
  assign _2851_ = dp2lut_Xinfo_7[17] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6935" *) raw_reg64 : _2785_;
  assign _2852_ = dp2lut_Xinfo_7[16] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6932" *) raw_reg0 : _2851_;
  assign _0276_ = _0399_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6931" *) _2852_ : lut_X_data_71;
  function [15:0] _6713_;
    input [15:0] a;
    input [1023:0] b;
    input [63:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:7196|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6939" *)
    (* parallel_case *)
    casez (s)
      64'b???????????????????????????????????????????????????????????????1:
        _6713_ = b[15:0];
      64'b??????????????????????????????????????????????????????????????1?:
        _6713_ = b[31:16];
      64'b?????????????????????????????????????????????????????????????1??:
        _6713_ = b[47:32];
      64'b????????????????????????????????????????????????????????????1???:
        _6713_ = b[63:48];
      64'b???????????????????????????????????????????????????????????1????:
        _6713_ = b[79:64];
      64'b??????????????????????????????????????????????????????????1?????:
        _6713_ = b[95:80];
      64'b?????????????????????????????????????????????????????????1??????:
        _6713_ = b[111:96];
      64'b????????????????????????????????????????????????????????1???????:
        _6713_ = b[127:112];
      64'b???????????????????????????????????????????????????????1????????:
        _6713_ = b[143:128];
      64'b??????????????????????????????????????????????????????1?????????:
        _6713_ = b[159:144];
      64'b?????????????????????????????????????????????????????1??????????:
        _6713_ = b[175:160];
      64'b????????????????????????????????????????????????????1???????????:
        _6713_ = b[191:176];
      64'b???????????????????????????????????????????????????1????????????:
        _6713_ = b[207:192];
      64'b??????????????????????????????????????????????????1?????????????:
        _6713_ = b[223:208];
      64'b?????????????????????????????????????????????????1??????????????:
        _6713_ = b[239:224];
      64'b????????????????????????????????????????????????1???????????????:
        _6713_ = b[255:240];
      64'b???????????????????????????????????????????????1????????????????:
        _6713_ = b[271:256];
      64'b??????????????????????????????????????????????1?????????????????:
        _6713_ = b[287:272];
      64'b?????????????????????????????????????????????1??????????????????:
        _6713_ = b[303:288];
      64'b????????????????????????????????????????????1???????????????????:
        _6713_ = b[319:304];
      64'b???????????????????????????????????????????1????????????????????:
        _6713_ = b[335:320];
      64'b??????????????????????????????????????????1?????????????????????:
        _6713_ = b[351:336];
      64'b?????????????????????????????????????????1??????????????????????:
        _6713_ = b[367:352];
      64'b????????????????????????????????????????1???????????????????????:
        _6713_ = b[383:368];
      64'b???????????????????????????????????????1????????????????????????:
        _6713_ = b[399:384];
      64'b??????????????????????????????????????1?????????????????????????:
        _6713_ = b[415:400];
      64'b?????????????????????????????????????1??????????????????????????:
        _6713_ = b[431:416];
      64'b????????????????????????????????????1???????????????????????????:
        _6713_ = b[447:432];
      64'b???????????????????????????????????1????????????????????????????:
        _6713_ = b[463:448];
      64'b??????????????????????????????????1?????????????????????????????:
        _6713_ = b[479:464];
      64'b?????????????????????????????????1??????????????????????????????:
        _6713_ = b[495:480];
      64'b????????????????????????????????1???????????????????????????????:
        _6713_ = b[511:496];
      64'b???????????????????????????????1????????????????????????????????:
        _6713_ = b[527:512];
      64'b??????????????????????????????1?????????????????????????????????:
        _6713_ = b[543:528];
      64'b?????????????????????????????1??????????????????????????????????:
        _6713_ = b[559:544];
      64'b????????????????????????????1???????????????????????????????????:
        _6713_ = b[575:560];
      64'b???????????????????????????1????????????????????????????????????:
        _6713_ = b[591:576];
      64'b??????????????????????????1?????????????????????????????????????:
        _6713_ = b[607:592];
      64'b?????????????????????????1??????????????????????????????????????:
        _6713_ = b[623:608];
      64'b????????????????????????1???????????????????????????????????????:
        _6713_ = b[639:624];
      64'b???????????????????????1????????????????????????????????????????:
        _6713_ = b[655:640];
      64'b??????????????????????1?????????????????????????????????????????:
        _6713_ = b[671:656];
      64'b?????????????????????1??????????????????????????????????????????:
        _6713_ = b[687:672];
      64'b????????????????????1???????????????????????????????????????????:
        _6713_ = b[703:688];
      64'b???????????????????1????????????????????????????????????????????:
        _6713_ = b[719:704];
      64'b??????????????????1?????????????????????????????????????????????:
        _6713_ = b[735:720];
      64'b?????????????????1??????????????????????????????????????????????:
        _6713_ = b[751:736];
      64'b????????????????1???????????????????????????????????????????????:
        _6713_ = b[767:752];
      64'b???????????????1????????????????????????????????????????????????:
        _6713_ = b[783:768];
      64'b??????????????1?????????????????????????????????????????????????:
        _6713_ = b[799:784];
      64'b?????????????1??????????????????????????????????????????????????:
        _6713_ = b[815:800];
      64'b????????????1???????????????????????????????????????????????????:
        _6713_ = b[831:816];
      64'b???????????1????????????????????????????????????????????????????:
        _6713_ = b[847:832];
      64'b??????????1?????????????????????????????????????????????????????:
        _6713_ = b[863:848];
      64'b?????????1??????????????????????????????????????????????????????:
        _6713_ = b[879:864];
      64'b????????1???????????????????????????????????????????????????????:
        _6713_ = b[895:880];
      64'b???????1????????????????????????????????????????????????????????:
        _6713_ = b[911:896];
      64'b??????1?????????????????????????????????????????????????????????:
        _6713_ = b[927:912];
      64'b?????1??????????????????????????????????????????????????????????:
        _6713_ = b[943:928];
      64'b????1???????????????????????????????????????????????????????????:
        _6713_ = b[959:944];
      64'b???1????????????????????????????????????????????????????????????:
        _6713_ = b[975:960];
      64'b??1?????????????????????????????????????????????????????????????:
        _6713_ = b[991:976];
      64'b?1??????????????????????????????????????????????????????????????:
        _6713_ = b[1007:992];
      64'b1???????????????????????????????????????????????????????????????:
        _6713_ = b[1023:1008];
      default:
        _6713_ = a;
    endcase
  endfunction
  assign _2853_ = _6713_(raw_reg0, { raw_reg1, raw_reg2, raw_reg3, raw_reg4, raw_reg5, raw_reg6, raw_reg7, raw_reg8, raw_reg9, raw_reg10, raw_reg11, raw_reg12, raw_reg13, raw_reg14, raw_reg15, raw_reg16, raw_reg17, raw_reg18, raw_reg19, raw_reg20, raw_reg21, raw_reg22, raw_reg23, raw_reg24, raw_reg25, raw_reg26, raw_reg27, raw_reg28, raw_reg29, raw_reg30, raw_reg31, raw_reg32, raw_reg33, raw_reg34, raw_reg35, raw_reg36, raw_reg37, raw_reg38, raw_reg39, raw_reg40, raw_reg41, raw_reg42, raw_reg43, raw_reg44, raw_reg45, raw_reg46, raw_reg47, raw_reg48, raw_reg49, raw_reg50, raw_reg51, raw_reg52, raw_reg53, raw_reg54, raw_reg55, raw_reg56, raw_reg57, raw_reg58, raw_reg59, raw_reg60, raw_reg61, raw_reg62, raw_reg63, raw_reg64 }, { _2849_, _2848_, _2847_, _2846_, _2845_, _2844_, _2843_, _2842_, _2841_, _2840_, _2839_, _2838_, _2837_, _2836_, _2835_, _2834_, _2833_, _2832_, _2831_, _2830_, _2829_, _2828_, _2827_, _2826_, _2825_, _2824_, _2823_, _2822_, _2821_, _2820_, _2819_, _2818_, _2817_, _2816_, _2815_, _2814_, _2813_, _2812_, _2811_, _2810_, _2809_, _2808_, _2807_, _2806_, _2805_, _2804_, _2803_, _2802_, _2801_, _2800_, _2799_, _2798_, _2797_, _2796_, _2795_, _2794_, _2793_, _2792_, _2791_, _2790_, _2789_, _2788_, _2787_, _2786_ });
  assign _2854_ = dp2lut_Xinfo_7[17] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6935" *) raw_reg64 : _2853_;
  assign _2855_ = dp2lut_Xinfo_7[16] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6932" *) raw_reg0 : _2854_;
  assign _0275_ = _0399_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6931" *) _2855_ : lut_X_data_70;
  function [15:0] _6717_;
    input [15:0] a;
    input [1023:0] b;
    input [63:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6913|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6656" *)
    (* parallel_case *)
    casez (s)
      64'b???????????????????????????????????????????????????????????????1:
        _6717_ = b[15:0];
      64'b??????????????????????????????????????????????????????????????1?:
        _6717_ = b[31:16];
      64'b?????????????????????????????????????????????????????????????1??:
        _6717_ = b[47:32];
      64'b????????????????????????????????????????????????????????????1???:
        _6717_ = b[63:48];
      64'b???????????????????????????????????????????????????????????1????:
        _6717_ = b[79:64];
      64'b??????????????????????????????????????????????????????????1?????:
        _6717_ = b[95:80];
      64'b?????????????????????????????????????????????????????????1??????:
        _6717_ = b[111:96];
      64'b????????????????????????????????????????????????????????1???????:
        _6717_ = b[127:112];
      64'b???????????????????????????????????????????????????????1????????:
        _6717_ = b[143:128];
      64'b??????????????????????????????????????????????????????1?????????:
        _6717_ = b[159:144];
      64'b?????????????????????????????????????????????????????1??????????:
        _6717_ = b[175:160];
      64'b????????????????????????????????????????????????????1???????????:
        _6717_ = b[191:176];
      64'b???????????????????????????????????????????????????1????????????:
        _6717_ = b[207:192];
      64'b??????????????????????????????????????????????????1?????????????:
        _6717_ = b[223:208];
      64'b?????????????????????????????????????????????????1??????????????:
        _6717_ = b[239:224];
      64'b????????????????????????????????????????????????1???????????????:
        _6717_ = b[255:240];
      64'b???????????????????????????????????????????????1????????????????:
        _6717_ = b[271:256];
      64'b??????????????????????????????????????????????1?????????????????:
        _6717_ = b[287:272];
      64'b?????????????????????????????????????????????1??????????????????:
        _6717_ = b[303:288];
      64'b????????????????????????????????????????????1???????????????????:
        _6717_ = b[319:304];
      64'b???????????????????????????????????????????1????????????????????:
        _6717_ = b[335:320];
      64'b??????????????????????????????????????????1?????????????????????:
        _6717_ = b[351:336];
      64'b?????????????????????????????????????????1??????????????????????:
        _6717_ = b[367:352];
      64'b????????????????????????????????????????1???????????????????????:
        _6717_ = b[383:368];
      64'b???????????????????????????????????????1????????????????????????:
        _6717_ = b[399:384];
      64'b??????????????????????????????????????1?????????????????????????:
        _6717_ = b[415:400];
      64'b?????????????????????????????????????1??????????????????????????:
        _6717_ = b[431:416];
      64'b????????????????????????????????????1???????????????????????????:
        _6717_ = b[447:432];
      64'b???????????????????????????????????1????????????????????????????:
        _6717_ = b[463:448];
      64'b??????????????????????????????????1?????????????????????????????:
        _6717_ = b[479:464];
      64'b?????????????????????????????????1??????????????????????????????:
        _6717_ = b[495:480];
      64'b????????????????????????????????1???????????????????????????????:
        _6717_ = b[511:496];
      64'b???????????????????????????????1????????????????????????????????:
        _6717_ = b[527:512];
      64'b??????????????????????????????1?????????????????????????????????:
        _6717_ = b[543:528];
      64'b?????????????????????????????1??????????????????????????????????:
        _6717_ = b[559:544];
      64'b????????????????????????????1???????????????????????????????????:
        _6717_ = b[575:560];
      64'b???????????????????????????1????????????????????????????????????:
        _6717_ = b[591:576];
      64'b??????????????????????????1?????????????????????????????????????:
        _6717_ = b[607:592];
      64'b?????????????????????????1??????????????????????????????????????:
        _6717_ = b[623:608];
      64'b????????????????????????1???????????????????????????????????????:
        _6717_ = b[639:624];
      64'b???????????????????????1????????????????????????????????????????:
        _6717_ = b[655:640];
      64'b??????????????????????1?????????????????????????????????????????:
        _6717_ = b[671:656];
      64'b?????????????????????1??????????????????????????????????????????:
        _6717_ = b[687:672];
      64'b????????????????????1???????????????????????????????????????????:
        _6717_ = b[703:688];
      64'b???????????????????1????????????????????????????????????????????:
        _6717_ = b[719:704];
      64'b??????????????????1?????????????????????????????????????????????:
        _6717_ = b[735:720];
      64'b?????????????????1??????????????????????????????????????????????:
        _6717_ = b[751:736];
      64'b????????????????1???????????????????????????????????????????????:
        _6717_ = b[767:752];
      64'b???????????????1????????????????????????????????????????????????:
        _6717_ = b[783:768];
      64'b??????????????1?????????????????????????????????????????????????:
        _6717_ = b[799:784];
      64'b?????????????1??????????????????????????????????????????????????:
        _6717_ = b[815:800];
      64'b????????????1???????????????????????????????????????????????????:
        _6717_ = b[831:816];
      64'b???????????1????????????????????????????????????????????????????:
        _6717_ = b[847:832];
      64'b??????????1?????????????????????????????????????????????????????:
        _6717_ = b[863:848];
      64'b?????????1??????????????????????????????????????????????????????:
        _6717_ = b[879:864];
      64'b????????1???????????????????????????????????????????????????????:
        _6717_ = b[895:880];
      64'b???????1????????????????????????????????????????????????????????:
        _6717_ = b[911:896];
      64'b??????1?????????????????????????????????????????????????????????:
        _6717_ = b[927:912];
      64'b?????1??????????????????????????????????????????????????????????:
        _6717_ = b[943:928];
      64'b????1???????????????????????????????????????????????????????????:
        _6717_ = b[959:944];
      64'b???1????????????????????????????????????????????????????????????:
        _6717_ = b[975:960];
      64'b??1?????????????????????????????????????????????????????????????:
        _6717_ = b[991:976];
      64'b?1??????????????????????????????????????????????????????????????:
        _6717_ = b[1007:992];
      64'b1???????????????????????????????????????????????????????????????:
        _6717_ = b[1023:1008];
      default:
        _6717_ = a;
    endcase
  endfunction
  assign _2856_ = _6717_(raw_reg0, { raw_reg1, raw_reg2, raw_reg3, raw_reg4, raw_reg5, raw_reg6, raw_reg7, raw_reg8, raw_reg9, raw_reg10, raw_reg11, raw_reg12, raw_reg13, raw_reg14, raw_reg15, raw_reg16, raw_reg17, raw_reg18, raw_reg19, raw_reg20, raw_reg21, raw_reg22, raw_reg23, raw_reg24, raw_reg25, raw_reg26, raw_reg27, raw_reg28, raw_reg29, raw_reg30, raw_reg31, raw_reg32, raw_reg33, raw_reg34, raw_reg35, raw_reg36, raw_reg37, raw_reg38, raw_reg39, raw_reg40, raw_reg41, raw_reg42, raw_reg43, raw_reg44, raw_reg45, raw_reg46, raw_reg47, raw_reg48, raw_reg49, raw_reg50, raw_reg51, raw_reg52, raw_reg53, raw_reg54, raw_reg55, raw_reg56, raw_reg57, raw_reg58, raw_reg59, raw_reg60, raw_reg61, raw_reg62, raw_reg63, raw_reg64 }, { _2921_, _2920_, _2919_, _2918_, _2917_, _2916_, _2915_, _2914_, _2913_, _2912_, _2911_, _2910_, _2909_, _2908_, _2907_, _2906_, _2905_, _2904_, _2903_, _2902_, _2901_, _2900_, _2899_, _2898_, _2897_, _2896_, _2895_, _2894_, _2893_, _2892_, _2891_, _2890_, _2889_, _2888_, _2887_, _2886_, _2885_, _2884_, _2883_, _2882_, _2881_, _2880_, _2879_, _2878_, _2877_, _2876_, _2875_, _2874_, _2873_, _2872_, _2871_, _2870_, _2869_, _2868_, _2867_, _2866_, _2865_, _2864_, _2863_, _2862_, _2861_, _2860_, _2859_, _0409_ });
  assign _2857_ = dp2lut_X_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6913|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6656" *) 7'b1000000;
  assign _2858_ = dp2lut_X_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6909|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6656" *) 6'b111111;
  assign _2859_ = dp2lut_X_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6905|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6656" *) 6'b111110;
  assign _2860_ = dp2lut_X_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6901|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6656" *) 6'b111101;
  assign _2861_ = dp2lut_X_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6897|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6656" *) 6'b111100;
  assign _2862_ = dp2lut_X_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6893|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6656" *) 6'b111011;
  assign _2863_ = dp2lut_X_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6889|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6656" *) 6'b111010;
  assign _2864_ = dp2lut_X_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6885|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6656" *) 6'b111001;
  assign _2865_ = dp2lut_X_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6881|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6656" *) 6'b111000;
  assign _2866_ = dp2lut_X_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6877|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6656" *) 6'b110111;
  assign _2867_ = dp2lut_X_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6873|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6656" *) 6'b110110;
  assign _2868_ = dp2lut_X_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6869|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6656" *) 6'b110101;
  assign _2869_ = dp2lut_X_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6865|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6656" *) 6'b110100;
  assign _2870_ = dp2lut_X_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6861|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6656" *) 6'b110011;
  assign _2871_ = dp2lut_X_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6857|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6656" *) 6'b110010;
  assign _2872_ = dp2lut_X_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6853|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6656" *) 6'b110001;
  assign _2873_ = dp2lut_X_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6849|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6656" *) 6'b110000;
  assign _2874_ = dp2lut_X_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6845|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6656" *) 6'b101111;
  assign _2875_ = dp2lut_X_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6841|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6656" *) 6'b101110;
  assign _2876_ = dp2lut_X_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6837|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6656" *) 6'b101101;
  assign _2877_ = dp2lut_X_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6833|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6656" *) 6'b101100;
  assign _2878_ = dp2lut_X_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6829|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6656" *) 6'b101011;
  assign _2879_ = dp2lut_X_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6825|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6656" *) 6'b101010;
  assign _2880_ = dp2lut_X_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6821|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6656" *) 6'b101001;
  assign _2881_ = dp2lut_X_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6817|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6656" *) 6'b101000;
  assign _2882_ = dp2lut_X_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6813|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6656" *) 6'b100111;
  assign _2883_ = dp2lut_X_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6809|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6656" *) 6'b100110;
  assign _2884_ = dp2lut_X_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6805|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6656" *) 6'b100101;
  assign _2885_ = dp2lut_X_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6801|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6656" *) 6'b100100;
  assign _2886_ = dp2lut_X_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6797|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6656" *) 6'b100011;
  assign _2887_ = dp2lut_X_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6793|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6656" *) 6'b100010;
  assign _2888_ = dp2lut_X_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6789|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6656" *) 6'b100001;
  assign _2889_ = dp2lut_X_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6785|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6656" *) 6'b100000;
  assign _2890_ = dp2lut_X_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6781|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6656" *) 5'b11111;
  assign _2891_ = dp2lut_X_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6777|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6656" *) 5'b11110;
  assign _2892_ = dp2lut_X_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6773|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6656" *) 5'b11101;
  assign _2893_ = dp2lut_X_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6769|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6656" *) 5'b11100;
  assign _2894_ = dp2lut_X_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6765|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6656" *) 5'b11011;
  assign _2895_ = dp2lut_X_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6761|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6656" *) 5'b11010;
  assign _2896_ = dp2lut_X_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6757|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6656" *) 5'b11001;
  assign _2897_ = dp2lut_X_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6753|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6656" *) 5'b11000;
  assign _2898_ = dp2lut_X_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6749|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6656" *) 5'b10111;
  assign _2899_ = dp2lut_X_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6745|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6656" *) 5'b10110;
  assign _2900_ = dp2lut_X_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6741|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6656" *) 5'b10101;
  assign _2901_ = dp2lut_X_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6737|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6656" *) 5'b10100;
  assign _2902_ = dp2lut_X_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6733|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6656" *) 5'b10011;
  assign _2903_ = dp2lut_X_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6729|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6656" *) 5'b10010;
  assign _2904_ = dp2lut_X_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6725|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6656" *) 5'b10001;
  assign _2905_ = dp2lut_X_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6721|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6656" *) 5'b10000;
  assign _2906_ = dp2lut_X_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6717|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6656" *) 4'b1111;
  assign _2907_ = dp2lut_X_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6713|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6656" *) 4'b1110;
  assign _2908_ = dp2lut_X_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6709|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6656" *) 4'b1101;
  assign _2909_ = dp2lut_X_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6705|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6656" *) 4'b1100;
  assign _2910_ = dp2lut_X_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6701|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6656" *) 4'b1011;
  assign _2911_ = dp2lut_X_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6697|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6656" *) 4'b1010;
  assign _2912_ = dp2lut_X_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6693|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6656" *) 4'b1001;
  assign _2913_ = dp2lut_X_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6689|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6656" *) 4'b1000;
  assign _2914_ = dp2lut_X_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6685|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6656" *) 3'b111;
  assign _2915_ = dp2lut_X_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6681|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6656" *) 3'b110;
  assign _2916_ = dp2lut_X_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6677|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6656" *) 3'b101;
  assign _2917_ = dp2lut_X_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6673|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6656" *) 3'b100;
  assign _2918_ = dp2lut_X_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6669|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6656" *) 2'b11;
  assign _2919_ = dp2lut_X_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6665|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6656" *) 2'b10;
  assign _2920_ = dp2lut_X_entry_6 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6661|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6656" *) 1'b1;
  assign _2921_ = ! (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6657|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6656" *) dp2lut_X_entry_6;
  assign _2922_ = dp2lut_Xinfo_6[17] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6652" *) raw_reg64 : _2856_;
  assign _2923_ = dp2lut_Xinfo_6[16] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6649" *) raw_reg0 : _2922_;
  assign _0274_ = _0398_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6648" *) _2923_ : lut_X_data_61;
  function [15:0] _6786_;
    input [15:0] a;
    input [1023:0] b;
    input [63:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6913|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6656" *)
    (* parallel_case *)
    casez (s)
      64'b???????????????????????????????????????????????????????????????1:
        _6786_ = b[15:0];
      64'b??????????????????????????????????????????????????????????????1?:
        _6786_ = b[31:16];
      64'b?????????????????????????????????????????????????????????????1??:
        _6786_ = b[47:32];
      64'b????????????????????????????????????????????????????????????1???:
        _6786_ = b[63:48];
      64'b???????????????????????????????????????????????????????????1????:
        _6786_ = b[79:64];
      64'b??????????????????????????????????????????????????????????1?????:
        _6786_ = b[95:80];
      64'b?????????????????????????????????????????????????????????1??????:
        _6786_ = b[111:96];
      64'b????????????????????????????????????????????????????????1???????:
        _6786_ = b[127:112];
      64'b???????????????????????????????????????????????????????1????????:
        _6786_ = b[143:128];
      64'b??????????????????????????????????????????????????????1?????????:
        _6786_ = b[159:144];
      64'b?????????????????????????????????????????????????????1??????????:
        _6786_ = b[175:160];
      64'b????????????????????????????????????????????????????1???????????:
        _6786_ = b[191:176];
      64'b???????????????????????????????????????????????????1????????????:
        _6786_ = b[207:192];
      64'b??????????????????????????????????????????????????1?????????????:
        _6786_ = b[223:208];
      64'b?????????????????????????????????????????????????1??????????????:
        _6786_ = b[239:224];
      64'b????????????????????????????????????????????????1???????????????:
        _6786_ = b[255:240];
      64'b???????????????????????????????????????????????1????????????????:
        _6786_ = b[271:256];
      64'b??????????????????????????????????????????????1?????????????????:
        _6786_ = b[287:272];
      64'b?????????????????????????????????????????????1??????????????????:
        _6786_ = b[303:288];
      64'b????????????????????????????????????????????1???????????????????:
        _6786_ = b[319:304];
      64'b???????????????????????????????????????????1????????????????????:
        _6786_ = b[335:320];
      64'b??????????????????????????????????????????1?????????????????????:
        _6786_ = b[351:336];
      64'b?????????????????????????????????????????1??????????????????????:
        _6786_ = b[367:352];
      64'b????????????????????????????????????????1???????????????????????:
        _6786_ = b[383:368];
      64'b???????????????????????????????????????1????????????????????????:
        _6786_ = b[399:384];
      64'b??????????????????????????????????????1?????????????????????????:
        _6786_ = b[415:400];
      64'b?????????????????????????????????????1??????????????????????????:
        _6786_ = b[431:416];
      64'b????????????????????????????????????1???????????????????????????:
        _6786_ = b[447:432];
      64'b???????????????????????????????????1????????????????????????????:
        _6786_ = b[463:448];
      64'b??????????????????????????????????1?????????????????????????????:
        _6786_ = b[479:464];
      64'b?????????????????????????????????1??????????????????????????????:
        _6786_ = b[495:480];
      64'b????????????????????????????????1???????????????????????????????:
        _6786_ = b[511:496];
      64'b???????????????????????????????1????????????????????????????????:
        _6786_ = b[527:512];
      64'b??????????????????????????????1?????????????????????????????????:
        _6786_ = b[543:528];
      64'b?????????????????????????????1??????????????????????????????????:
        _6786_ = b[559:544];
      64'b????????????????????????????1???????????????????????????????????:
        _6786_ = b[575:560];
      64'b???????????????????????????1????????????????????????????????????:
        _6786_ = b[591:576];
      64'b??????????????????????????1?????????????????????????????????????:
        _6786_ = b[607:592];
      64'b?????????????????????????1??????????????????????????????????????:
        _6786_ = b[623:608];
      64'b????????????????????????1???????????????????????????????????????:
        _6786_ = b[639:624];
      64'b???????????????????????1????????????????????????????????????????:
        _6786_ = b[655:640];
      64'b??????????????????????1?????????????????????????????????????????:
        _6786_ = b[671:656];
      64'b?????????????????????1??????????????????????????????????????????:
        _6786_ = b[687:672];
      64'b????????????????????1???????????????????????????????????????????:
        _6786_ = b[703:688];
      64'b???????????????????1????????????????????????????????????????????:
        _6786_ = b[719:704];
      64'b??????????????????1?????????????????????????????????????????????:
        _6786_ = b[735:720];
      64'b?????????????????1??????????????????????????????????????????????:
        _6786_ = b[751:736];
      64'b????????????????1???????????????????????????????????????????????:
        _6786_ = b[767:752];
      64'b???????????????1????????????????????????????????????????????????:
        _6786_ = b[783:768];
      64'b??????????????1?????????????????????????????????????????????????:
        _6786_ = b[799:784];
      64'b?????????????1??????????????????????????????????????????????????:
        _6786_ = b[815:800];
      64'b????????????1???????????????????????????????????????????????????:
        _6786_ = b[831:816];
      64'b???????????1????????????????????????????????????????????????????:
        _6786_ = b[847:832];
      64'b??????????1?????????????????????????????????????????????????????:
        _6786_ = b[863:848];
      64'b?????????1??????????????????????????????????????????????????????:
        _6786_ = b[879:864];
      64'b????????1???????????????????????????????????????????????????????:
        _6786_ = b[895:880];
      64'b???????1????????????????????????????????????????????????????????:
        _6786_ = b[911:896];
      64'b??????1?????????????????????????????????????????????????????????:
        _6786_ = b[927:912];
      64'b?????1??????????????????????????????????????????????????????????:
        _6786_ = b[943:928];
      64'b????1???????????????????????????????????????????????????????????:
        _6786_ = b[959:944];
      64'b???1????????????????????????????????????????????????????????????:
        _6786_ = b[975:960];
      64'b??1?????????????????????????????????????????????????????????????:
        _6786_ = b[991:976];
      64'b?1??????????????????????????????????????????????????????????????:
        _6786_ = b[1007:992];
      64'b1???????????????????????????????????????????????????????????????:
        _6786_ = b[1023:1008];
      default:
        _6786_ = a;
    endcase
  endfunction
  assign _2924_ = _6786_(raw_reg0, { raw_reg1, raw_reg2, raw_reg3, raw_reg4, raw_reg5, raw_reg6, raw_reg7, raw_reg8, raw_reg9, raw_reg10, raw_reg11, raw_reg12, raw_reg13, raw_reg14, raw_reg15, raw_reg16, raw_reg17, raw_reg18, raw_reg19, raw_reg20, raw_reg21, raw_reg22, raw_reg23, raw_reg24, raw_reg25, raw_reg26, raw_reg27, raw_reg28, raw_reg29, raw_reg30, raw_reg31, raw_reg32, raw_reg33, raw_reg34, raw_reg35, raw_reg36, raw_reg37, raw_reg38, raw_reg39, raw_reg40, raw_reg41, raw_reg42, raw_reg43, raw_reg44, raw_reg45, raw_reg46, raw_reg47, raw_reg48, raw_reg49, raw_reg50, raw_reg51, raw_reg52, raw_reg53, raw_reg54, raw_reg55, raw_reg56, raw_reg57, raw_reg58, raw_reg59, raw_reg60, raw_reg61, raw_reg62, raw_reg63, raw_reg64 }, { _2920_, _2919_, _2918_, _2917_, _2916_, _2915_, _2914_, _2913_, _2912_, _2911_, _2910_, _2909_, _2908_, _2907_, _2906_, _2905_, _2904_, _2903_, _2902_, _2901_, _2900_, _2899_, _2898_, _2897_, _2896_, _2895_, _2894_, _2893_, _2892_, _2891_, _2890_, _2889_, _2888_, _2887_, _2886_, _2885_, _2884_, _2883_, _2882_, _2881_, _2880_, _2879_, _2878_, _2877_, _2876_, _2875_, _2874_, _2873_, _2872_, _2871_, _2870_, _2869_, _2868_, _2867_, _2866_, _2865_, _2864_, _2863_, _2862_, _2861_, _2860_, _2859_, _2858_, _2857_ });
  assign _2925_ = dp2lut_Xinfo_6[17] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6652" *) raw_reg64 : _2924_;
  assign _2926_ = dp2lut_Xinfo_6[16] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6649" *) raw_reg0 : _2925_;
  assign _0273_ = _0398_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6648" *) _2926_ : lut_X_data_60;
  function [15:0] _6790_;
    input [15:0] a;
    input [1023:0] b;
    input [63:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6630|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6373" *)
    (* parallel_case *)
    casez (s)
      64'b???????????????????????????????????????????????????????????????1:
        _6790_ = b[15:0];
      64'b??????????????????????????????????????????????????????????????1?:
        _6790_ = b[31:16];
      64'b?????????????????????????????????????????????????????????????1??:
        _6790_ = b[47:32];
      64'b????????????????????????????????????????????????????????????1???:
        _6790_ = b[63:48];
      64'b???????????????????????????????????????????????????????????1????:
        _6790_ = b[79:64];
      64'b??????????????????????????????????????????????????????????1?????:
        _6790_ = b[95:80];
      64'b?????????????????????????????????????????????????????????1??????:
        _6790_ = b[111:96];
      64'b????????????????????????????????????????????????????????1???????:
        _6790_ = b[127:112];
      64'b???????????????????????????????????????????????????????1????????:
        _6790_ = b[143:128];
      64'b??????????????????????????????????????????????????????1?????????:
        _6790_ = b[159:144];
      64'b?????????????????????????????????????????????????????1??????????:
        _6790_ = b[175:160];
      64'b????????????????????????????????????????????????????1???????????:
        _6790_ = b[191:176];
      64'b???????????????????????????????????????????????????1????????????:
        _6790_ = b[207:192];
      64'b??????????????????????????????????????????????????1?????????????:
        _6790_ = b[223:208];
      64'b?????????????????????????????????????????????????1??????????????:
        _6790_ = b[239:224];
      64'b????????????????????????????????????????????????1???????????????:
        _6790_ = b[255:240];
      64'b???????????????????????????????????????????????1????????????????:
        _6790_ = b[271:256];
      64'b??????????????????????????????????????????????1?????????????????:
        _6790_ = b[287:272];
      64'b?????????????????????????????????????????????1??????????????????:
        _6790_ = b[303:288];
      64'b????????????????????????????????????????????1???????????????????:
        _6790_ = b[319:304];
      64'b???????????????????????????????????????????1????????????????????:
        _6790_ = b[335:320];
      64'b??????????????????????????????????????????1?????????????????????:
        _6790_ = b[351:336];
      64'b?????????????????????????????????????????1??????????????????????:
        _6790_ = b[367:352];
      64'b????????????????????????????????????????1???????????????????????:
        _6790_ = b[383:368];
      64'b???????????????????????????????????????1????????????????????????:
        _6790_ = b[399:384];
      64'b??????????????????????????????????????1?????????????????????????:
        _6790_ = b[415:400];
      64'b?????????????????????????????????????1??????????????????????????:
        _6790_ = b[431:416];
      64'b????????????????????????????????????1???????????????????????????:
        _6790_ = b[447:432];
      64'b???????????????????????????????????1????????????????????????????:
        _6790_ = b[463:448];
      64'b??????????????????????????????????1?????????????????????????????:
        _6790_ = b[479:464];
      64'b?????????????????????????????????1??????????????????????????????:
        _6790_ = b[495:480];
      64'b????????????????????????????????1???????????????????????????????:
        _6790_ = b[511:496];
      64'b???????????????????????????????1????????????????????????????????:
        _6790_ = b[527:512];
      64'b??????????????????????????????1?????????????????????????????????:
        _6790_ = b[543:528];
      64'b?????????????????????????????1??????????????????????????????????:
        _6790_ = b[559:544];
      64'b????????????????????????????1???????????????????????????????????:
        _6790_ = b[575:560];
      64'b???????????????????????????1????????????????????????????????????:
        _6790_ = b[591:576];
      64'b??????????????????????????1?????????????????????????????????????:
        _6790_ = b[607:592];
      64'b?????????????????????????1??????????????????????????????????????:
        _6790_ = b[623:608];
      64'b????????????????????????1???????????????????????????????????????:
        _6790_ = b[639:624];
      64'b???????????????????????1????????????????????????????????????????:
        _6790_ = b[655:640];
      64'b??????????????????????1?????????????????????????????????????????:
        _6790_ = b[671:656];
      64'b?????????????????????1??????????????????????????????????????????:
        _6790_ = b[687:672];
      64'b????????????????????1???????????????????????????????????????????:
        _6790_ = b[703:688];
      64'b???????????????????1????????????????????????????????????????????:
        _6790_ = b[719:704];
      64'b??????????????????1?????????????????????????????????????????????:
        _6790_ = b[735:720];
      64'b?????????????????1??????????????????????????????????????????????:
        _6790_ = b[751:736];
      64'b????????????????1???????????????????????????????????????????????:
        _6790_ = b[767:752];
      64'b???????????????1????????????????????????????????????????????????:
        _6790_ = b[783:768];
      64'b??????????????1?????????????????????????????????????????????????:
        _6790_ = b[799:784];
      64'b?????????????1??????????????????????????????????????????????????:
        _6790_ = b[815:800];
      64'b????????????1???????????????????????????????????????????????????:
        _6790_ = b[831:816];
      64'b???????????1????????????????????????????????????????????????????:
        _6790_ = b[847:832];
      64'b??????????1?????????????????????????????????????????????????????:
        _6790_ = b[863:848];
      64'b?????????1??????????????????????????????????????????????????????:
        _6790_ = b[879:864];
      64'b????????1???????????????????????????????????????????????????????:
        _6790_ = b[895:880];
      64'b???????1????????????????????????????????????????????????????????:
        _6790_ = b[911:896];
      64'b??????1?????????????????????????????????????????????????????????:
        _6790_ = b[927:912];
      64'b?????1??????????????????????????????????????????????????????????:
        _6790_ = b[943:928];
      64'b????1???????????????????????????????????????????????????????????:
        _6790_ = b[959:944];
      64'b???1????????????????????????????????????????????????????????????:
        _6790_ = b[975:960];
      64'b??1?????????????????????????????????????????????????????????????:
        _6790_ = b[991:976];
      64'b?1??????????????????????????????????????????????????????????????:
        _6790_ = b[1007:992];
      64'b1???????????????????????????????????????????????????????????????:
        _6790_ = b[1023:1008];
      default:
        _6790_ = a;
    endcase
  endfunction
  assign _2927_ = _6790_(raw_reg0, { raw_reg1, raw_reg2, raw_reg3, raw_reg4, raw_reg5, raw_reg6, raw_reg7, raw_reg8, raw_reg9, raw_reg10, raw_reg11, raw_reg12, raw_reg13, raw_reg14, raw_reg15, raw_reg16, raw_reg17, raw_reg18, raw_reg19, raw_reg20, raw_reg21, raw_reg22, raw_reg23, raw_reg24, raw_reg25, raw_reg26, raw_reg27, raw_reg28, raw_reg29, raw_reg30, raw_reg31, raw_reg32, raw_reg33, raw_reg34, raw_reg35, raw_reg36, raw_reg37, raw_reg38, raw_reg39, raw_reg40, raw_reg41, raw_reg42, raw_reg43, raw_reg44, raw_reg45, raw_reg46, raw_reg47, raw_reg48, raw_reg49, raw_reg50, raw_reg51, raw_reg52, raw_reg53, raw_reg54, raw_reg55, raw_reg56, raw_reg57, raw_reg58, raw_reg59, raw_reg60, raw_reg61, raw_reg62, raw_reg63, raw_reg64 }, { _2992_, _2991_, _2990_, _2989_, _2988_, _2987_, _2986_, _2985_, _2984_, _2983_, _2982_, _2981_, _2980_, _2979_, _2978_, _2977_, _2976_, _2975_, _2974_, _2973_, _2972_, _2971_, _2970_, _2969_, _2968_, _2967_, _2966_, _2965_, _2964_, _2963_, _2962_, _2961_, _2960_, _2959_, _2958_, _2957_, _2956_, _2955_, _2954_, _2953_, _2952_, _2951_, _2950_, _2949_, _2948_, _2947_, _2946_, _2945_, _2944_, _2943_, _2942_, _2941_, _2940_, _2939_, _2938_, _2937_, _2936_, _2935_, _2934_, _2933_, _2932_, _2931_, _2930_, _0410_ });
  assign _2928_ = dp2lut_X_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6630|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6373" *) 7'b1000000;
  assign _2929_ = dp2lut_X_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6626|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6373" *) 6'b111111;
  assign _2930_ = dp2lut_X_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6622|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6373" *) 6'b111110;
  assign _2931_ = dp2lut_X_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6618|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6373" *) 6'b111101;
  assign _2932_ = dp2lut_X_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6614|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6373" *) 6'b111100;
  assign _2933_ = dp2lut_X_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6610|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6373" *) 6'b111011;
  assign _2934_ = dp2lut_X_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6606|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6373" *) 6'b111010;
  assign _2935_ = dp2lut_X_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6602|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6373" *) 6'b111001;
  assign _2936_ = dp2lut_X_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6598|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6373" *) 6'b111000;
  assign _2937_ = dp2lut_X_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6594|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6373" *) 6'b110111;
  assign _2938_ = dp2lut_X_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6590|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6373" *) 6'b110110;
  assign _2939_ = dp2lut_X_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6586|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6373" *) 6'b110101;
  assign _2940_ = dp2lut_X_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6582|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6373" *) 6'b110100;
  assign _2941_ = dp2lut_X_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6578|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6373" *) 6'b110011;
  assign _2942_ = dp2lut_X_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6574|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6373" *) 6'b110010;
  assign _2943_ = dp2lut_X_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6570|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6373" *) 6'b110001;
  assign _2944_ = dp2lut_X_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6566|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6373" *) 6'b110000;
  assign _2945_ = dp2lut_X_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6562|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6373" *) 6'b101111;
  assign _2946_ = dp2lut_X_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6558|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6373" *) 6'b101110;
  assign _2947_ = dp2lut_X_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6554|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6373" *) 6'b101101;
  assign _2948_ = dp2lut_X_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6550|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6373" *) 6'b101100;
  assign _2949_ = dp2lut_X_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6546|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6373" *) 6'b101011;
  assign _2950_ = dp2lut_X_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6542|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6373" *) 6'b101010;
  assign _2951_ = dp2lut_X_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6538|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6373" *) 6'b101001;
  assign _2952_ = dp2lut_X_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6534|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6373" *) 6'b101000;
  assign _2953_ = dp2lut_X_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6530|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6373" *) 6'b100111;
  assign _2954_ = dp2lut_X_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6526|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6373" *) 6'b100110;
  assign _2955_ = dp2lut_X_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6522|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6373" *) 6'b100101;
  assign _2956_ = dp2lut_X_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6518|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6373" *) 6'b100100;
  assign _2957_ = dp2lut_X_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6514|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6373" *) 6'b100011;
  assign _2958_ = dp2lut_X_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6510|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6373" *) 6'b100010;
  assign _2959_ = dp2lut_X_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6506|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6373" *) 6'b100001;
  assign _2960_ = dp2lut_X_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6502|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6373" *) 6'b100000;
  assign _2961_ = dp2lut_X_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6498|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6373" *) 5'b11111;
  assign _2962_ = dp2lut_X_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6494|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6373" *) 5'b11110;
  assign _2963_ = dp2lut_X_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6490|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6373" *) 5'b11101;
  assign _2964_ = dp2lut_X_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6486|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6373" *) 5'b11100;
  assign _2965_ = dp2lut_X_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6482|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6373" *) 5'b11011;
  assign _2966_ = dp2lut_X_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6478|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6373" *) 5'b11010;
  assign _2967_ = dp2lut_X_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6474|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6373" *) 5'b11001;
  assign _2968_ = dp2lut_X_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6470|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6373" *) 5'b11000;
  assign _2969_ = dp2lut_X_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6466|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6373" *) 5'b10111;
  assign _2970_ = dp2lut_X_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6462|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6373" *) 5'b10110;
  assign _2971_ = dp2lut_X_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6458|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6373" *) 5'b10101;
  assign _2972_ = dp2lut_X_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6454|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6373" *) 5'b10100;
  assign _2973_ = dp2lut_X_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6450|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6373" *) 5'b10011;
  assign _2974_ = dp2lut_X_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6446|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6373" *) 5'b10010;
  assign _2975_ = dp2lut_X_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6442|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6373" *) 5'b10001;
  assign _2976_ = dp2lut_X_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6438|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6373" *) 5'b10000;
  assign _2977_ = dp2lut_X_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6434|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6373" *) 4'b1111;
  assign _2978_ = dp2lut_X_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6430|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6373" *) 4'b1110;
  assign _2979_ = dp2lut_X_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6426|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6373" *) 4'b1101;
  assign _2980_ = dp2lut_X_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6422|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6373" *) 4'b1100;
  assign _2981_ = dp2lut_X_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6418|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6373" *) 4'b1011;
  assign _2982_ = dp2lut_X_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6414|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6373" *) 4'b1010;
  assign _2983_ = dp2lut_X_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6410|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6373" *) 4'b1001;
  assign _2984_ = dp2lut_X_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6406|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6373" *) 4'b1000;
  assign _2985_ = dp2lut_X_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6402|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6373" *) 3'b111;
  assign _2986_ = dp2lut_X_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6398|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6373" *) 3'b110;
  assign _2987_ = dp2lut_X_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6394|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6373" *) 3'b101;
  assign _2988_ = dp2lut_X_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6390|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6373" *) 3'b100;
  assign _2989_ = dp2lut_X_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6386|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6373" *) 2'b11;
  assign _2990_ = dp2lut_X_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6382|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6373" *) 2'b10;
  assign _2991_ = dp2lut_X_entry_5 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6378|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6373" *) 1'b1;
  assign _2992_ = ! (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6374|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6373" *) dp2lut_X_entry_5;
  assign _2993_ = dp2lut_Xinfo_5[17] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6369" *) raw_reg64 : _2927_;
  assign _2994_ = dp2lut_Xinfo_5[16] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6366" *) raw_reg0 : _2993_;
  assign _0272_ = _0397_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6365" *) _2994_ : lut_X_data_51;
  function [15:0] _6859_;
    input [15:0] a;
    input [1023:0] b;
    input [63:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6630|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6373" *)
    (* parallel_case *)
    casez (s)
      64'b???????????????????????????????????????????????????????????????1:
        _6859_ = b[15:0];
      64'b??????????????????????????????????????????????????????????????1?:
        _6859_ = b[31:16];
      64'b?????????????????????????????????????????????????????????????1??:
        _6859_ = b[47:32];
      64'b????????????????????????????????????????????????????????????1???:
        _6859_ = b[63:48];
      64'b???????????????????????????????????????????????????????????1????:
        _6859_ = b[79:64];
      64'b??????????????????????????????????????????????????????????1?????:
        _6859_ = b[95:80];
      64'b?????????????????????????????????????????????????????????1??????:
        _6859_ = b[111:96];
      64'b????????????????????????????????????????????????????????1???????:
        _6859_ = b[127:112];
      64'b???????????????????????????????????????????????????????1????????:
        _6859_ = b[143:128];
      64'b??????????????????????????????????????????????????????1?????????:
        _6859_ = b[159:144];
      64'b?????????????????????????????????????????????????????1??????????:
        _6859_ = b[175:160];
      64'b????????????????????????????????????????????????????1???????????:
        _6859_ = b[191:176];
      64'b???????????????????????????????????????????????????1????????????:
        _6859_ = b[207:192];
      64'b??????????????????????????????????????????????????1?????????????:
        _6859_ = b[223:208];
      64'b?????????????????????????????????????????????????1??????????????:
        _6859_ = b[239:224];
      64'b????????????????????????????????????????????????1???????????????:
        _6859_ = b[255:240];
      64'b???????????????????????????????????????????????1????????????????:
        _6859_ = b[271:256];
      64'b??????????????????????????????????????????????1?????????????????:
        _6859_ = b[287:272];
      64'b?????????????????????????????????????????????1??????????????????:
        _6859_ = b[303:288];
      64'b????????????????????????????????????????????1???????????????????:
        _6859_ = b[319:304];
      64'b???????????????????????????????????????????1????????????????????:
        _6859_ = b[335:320];
      64'b??????????????????????????????????????????1?????????????????????:
        _6859_ = b[351:336];
      64'b?????????????????????????????????????????1??????????????????????:
        _6859_ = b[367:352];
      64'b????????????????????????????????????????1???????????????????????:
        _6859_ = b[383:368];
      64'b???????????????????????????????????????1????????????????????????:
        _6859_ = b[399:384];
      64'b??????????????????????????????????????1?????????????????????????:
        _6859_ = b[415:400];
      64'b?????????????????????????????????????1??????????????????????????:
        _6859_ = b[431:416];
      64'b????????????????????????????????????1???????????????????????????:
        _6859_ = b[447:432];
      64'b???????????????????????????????????1????????????????????????????:
        _6859_ = b[463:448];
      64'b??????????????????????????????????1?????????????????????????????:
        _6859_ = b[479:464];
      64'b?????????????????????????????????1??????????????????????????????:
        _6859_ = b[495:480];
      64'b????????????????????????????????1???????????????????????????????:
        _6859_ = b[511:496];
      64'b???????????????????????????????1????????????????????????????????:
        _6859_ = b[527:512];
      64'b??????????????????????????????1?????????????????????????????????:
        _6859_ = b[543:528];
      64'b?????????????????????????????1??????????????????????????????????:
        _6859_ = b[559:544];
      64'b????????????????????????????1???????????????????????????????????:
        _6859_ = b[575:560];
      64'b???????????????????????????1????????????????????????????????????:
        _6859_ = b[591:576];
      64'b??????????????????????????1?????????????????????????????????????:
        _6859_ = b[607:592];
      64'b?????????????????????????1??????????????????????????????????????:
        _6859_ = b[623:608];
      64'b????????????????????????1???????????????????????????????????????:
        _6859_ = b[639:624];
      64'b???????????????????????1????????????????????????????????????????:
        _6859_ = b[655:640];
      64'b??????????????????????1?????????????????????????????????????????:
        _6859_ = b[671:656];
      64'b?????????????????????1??????????????????????????????????????????:
        _6859_ = b[687:672];
      64'b????????????????????1???????????????????????????????????????????:
        _6859_ = b[703:688];
      64'b???????????????????1????????????????????????????????????????????:
        _6859_ = b[719:704];
      64'b??????????????????1?????????????????????????????????????????????:
        _6859_ = b[735:720];
      64'b?????????????????1??????????????????????????????????????????????:
        _6859_ = b[751:736];
      64'b????????????????1???????????????????????????????????????????????:
        _6859_ = b[767:752];
      64'b???????????????1????????????????????????????????????????????????:
        _6859_ = b[783:768];
      64'b??????????????1?????????????????????????????????????????????????:
        _6859_ = b[799:784];
      64'b?????????????1??????????????????????????????????????????????????:
        _6859_ = b[815:800];
      64'b????????????1???????????????????????????????????????????????????:
        _6859_ = b[831:816];
      64'b???????????1????????????????????????????????????????????????????:
        _6859_ = b[847:832];
      64'b??????????1?????????????????????????????????????????????????????:
        _6859_ = b[863:848];
      64'b?????????1??????????????????????????????????????????????????????:
        _6859_ = b[879:864];
      64'b????????1???????????????????????????????????????????????????????:
        _6859_ = b[895:880];
      64'b???????1????????????????????????????????????????????????????????:
        _6859_ = b[911:896];
      64'b??????1?????????????????????????????????????????????????????????:
        _6859_ = b[927:912];
      64'b?????1??????????????????????????????????????????????????????????:
        _6859_ = b[943:928];
      64'b????1???????????????????????????????????????????????????????????:
        _6859_ = b[959:944];
      64'b???1????????????????????????????????????????????????????????????:
        _6859_ = b[975:960];
      64'b??1?????????????????????????????????????????????????????????????:
        _6859_ = b[991:976];
      64'b?1??????????????????????????????????????????????????????????????:
        _6859_ = b[1007:992];
      64'b1???????????????????????????????????????????????????????????????:
        _6859_ = b[1023:1008];
      default:
        _6859_ = a;
    endcase
  endfunction
  assign _2995_ = _6859_(raw_reg0, { raw_reg1, raw_reg2, raw_reg3, raw_reg4, raw_reg5, raw_reg6, raw_reg7, raw_reg8, raw_reg9, raw_reg10, raw_reg11, raw_reg12, raw_reg13, raw_reg14, raw_reg15, raw_reg16, raw_reg17, raw_reg18, raw_reg19, raw_reg20, raw_reg21, raw_reg22, raw_reg23, raw_reg24, raw_reg25, raw_reg26, raw_reg27, raw_reg28, raw_reg29, raw_reg30, raw_reg31, raw_reg32, raw_reg33, raw_reg34, raw_reg35, raw_reg36, raw_reg37, raw_reg38, raw_reg39, raw_reg40, raw_reg41, raw_reg42, raw_reg43, raw_reg44, raw_reg45, raw_reg46, raw_reg47, raw_reg48, raw_reg49, raw_reg50, raw_reg51, raw_reg52, raw_reg53, raw_reg54, raw_reg55, raw_reg56, raw_reg57, raw_reg58, raw_reg59, raw_reg60, raw_reg61, raw_reg62, raw_reg63, raw_reg64 }, { _2991_, _2990_, _2989_, _2988_, _2987_, _2986_, _2985_, _2984_, _2983_, _2982_, _2981_, _2980_, _2979_, _2978_, _2977_, _2976_, _2975_, _2974_, _2973_, _2972_, _2971_, _2970_, _2969_, _2968_, _2967_, _2966_, _2965_, _2964_, _2963_, _2962_, _2961_, _2960_, _2959_, _2958_, _2957_, _2956_, _2955_, _2954_, _2953_, _2952_, _2951_, _2950_, _2949_, _2948_, _2947_, _2946_, _2945_, _2944_, _2943_, _2942_, _2941_, _2940_, _2939_, _2938_, _2937_, _2936_, _2935_, _2934_, _2933_, _2932_, _2931_, _2930_, _2929_, _2928_ });
  assign _2996_ = dp2lut_Xinfo_5[17] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6369" *) raw_reg64 : _2995_;
  assign _2997_ = dp2lut_Xinfo_5[16] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6366" *) raw_reg0 : _2996_;
  assign _0271_ = _0397_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6365" *) _2997_ : lut_X_data_50;
  function [15:0] _6863_;
    input [15:0] a;
    input [1023:0] b;
    input [63:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6347|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6090" *)
    (* parallel_case *)
    casez (s)
      64'b???????????????????????????????????????????????????????????????1:
        _6863_ = b[15:0];
      64'b??????????????????????????????????????????????????????????????1?:
        _6863_ = b[31:16];
      64'b?????????????????????????????????????????????????????????????1??:
        _6863_ = b[47:32];
      64'b????????????????????????????????????????????????????????????1???:
        _6863_ = b[63:48];
      64'b???????????????????????????????????????????????????????????1????:
        _6863_ = b[79:64];
      64'b??????????????????????????????????????????????????????????1?????:
        _6863_ = b[95:80];
      64'b?????????????????????????????????????????????????????????1??????:
        _6863_ = b[111:96];
      64'b????????????????????????????????????????????????????????1???????:
        _6863_ = b[127:112];
      64'b???????????????????????????????????????????????????????1????????:
        _6863_ = b[143:128];
      64'b??????????????????????????????????????????????????????1?????????:
        _6863_ = b[159:144];
      64'b?????????????????????????????????????????????????????1??????????:
        _6863_ = b[175:160];
      64'b????????????????????????????????????????????????????1???????????:
        _6863_ = b[191:176];
      64'b???????????????????????????????????????????????????1????????????:
        _6863_ = b[207:192];
      64'b??????????????????????????????????????????????????1?????????????:
        _6863_ = b[223:208];
      64'b?????????????????????????????????????????????????1??????????????:
        _6863_ = b[239:224];
      64'b????????????????????????????????????????????????1???????????????:
        _6863_ = b[255:240];
      64'b???????????????????????????????????????????????1????????????????:
        _6863_ = b[271:256];
      64'b??????????????????????????????????????????????1?????????????????:
        _6863_ = b[287:272];
      64'b?????????????????????????????????????????????1??????????????????:
        _6863_ = b[303:288];
      64'b????????????????????????????????????????????1???????????????????:
        _6863_ = b[319:304];
      64'b???????????????????????????????????????????1????????????????????:
        _6863_ = b[335:320];
      64'b??????????????????????????????????????????1?????????????????????:
        _6863_ = b[351:336];
      64'b?????????????????????????????????????????1??????????????????????:
        _6863_ = b[367:352];
      64'b????????????????????????????????????????1???????????????????????:
        _6863_ = b[383:368];
      64'b???????????????????????????????????????1????????????????????????:
        _6863_ = b[399:384];
      64'b??????????????????????????????????????1?????????????????????????:
        _6863_ = b[415:400];
      64'b?????????????????????????????????????1??????????????????????????:
        _6863_ = b[431:416];
      64'b????????????????????????????????????1???????????????????????????:
        _6863_ = b[447:432];
      64'b???????????????????????????????????1????????????????????????????:
        _6863_ = b[463:448];
      64'b??????????????????????????????????1?????????????????????????????:
        _6863_ = b[479:464];
      64'b?????????????????????????????????1??????????????????????????????:
        _6863_ = b[495:480];
      64'b????????????????????????????????1???????????????????????????????:
        _6863_ = b[511:496];
      64'b???????????????????????????????1????????????????????????????????:
        _6863_ = b[527:512];
      64'b??????????????????????????????1?????????????????????????????????:
        _6863_ = b[543:528];
      64'b?????????????????????????????1??????????????????????????????????:
        _6863_ = b[559:544];
      64'b????????????????????????????1???????????????????????????????????:
        _6863_ = b[575:560];
      64'b???????????????????????????1????????????????????????????????????:
        _6863_ = b[591:576];
      64'b??????????????????????????1?????????????????????????????????????:
        _6863_ = b[607:592];
      64'b?????????????????????????1??????????????????????????????????????:
        _6863_ = b[623:608];
      64'b????????????????????????1???????????????????????????????????????:
        _6863_ = b[639:624];
      64'b???????????????????????1????????????????????????????????????????:
        _6863_ = b[655:640];
      64'b??????????????????????1?????????????????????????????????????????:
        _6863_ = b[671:656];
      64'b?????????????????????1??????????????????????????????????????????:
        _6863_ = b[687:672];
      64'b????????????????????1???????????????????????????????????????????:
        _6863_ = b[703:688];
      64'b???????????????????1????????????????????????????????????????????:
        _6863_ = b[719:704];
      64'b??????????????????1?????????????????????????????????????????????:
        _6863_ = b[735:720];
      64'b?????????????????1??????????????????????????????????????????????:
        _6863_ = b[751:736];
      64'b????????????????1???????????????????????????????????????????????:
        _6863_ = b[767:752];
      64'b???????????????1????????????????????????????????????????????????:
        _6863_ = b[783:768];
      64'b??????????????1?????????????????????????????????????????????????:
        _6863_ = b[799:784];
      64'b?????????????1??????????????????????????????????????????????????:
        _6863_ = b[815:800];
      64'b????????????1???????????????????????????????????????????????????:
        _6863_ = b[831:816];
      64'b???????????1????????????????????????????????????????????????????:
        _6863_ = b[847:832];
      64'b??????????1?????????????????????????????????????????????????????:
        _6863_ = b[863:848];
      64'b?????????1??????????????????????????????????????????????????????:
        _6863_ = b[879:864];
      64'b????????1???????????????????????????????????????????????????????:
        _6863_ = b[895:880];
      64'b???????1????????????????????????????????????????????????????????:
        _6863_ = b[911:896];
      64'b??????1?????????????????????????????????????????????????????????:
        _6863_ = b[927:912];
      64'b?????1??????????????????????????????????????????????????????????:
        _6863_ = b[943:928];
      64'b????1???????????????????????????????????????????????????????????:
        _6863_ = b[959:944];
      64'b???1????????????????????????????????????????????????????????????:
        _6863_ = b[975:960];
      64'b??1?????????????????????????????????????????????????????????????:
        _6863_ = b[991:976];
      64'b?1??????????????????????????????????????????????????????????????:
        _6863_ = b[1007:992];
      64'b1???????????????????????????????????????????????????????????????:
        _6863_ = b[1023:1008];
      default:
        _6863_ = a;
    endcase
  endfunction
  assign _2998_ = _6863_(raw_reg0, { raw_reg1, raw_reg2, raw_reg3, raw_reg4, raw_reg5, raw_reg6, raw_reg7, raw_reg8, raw_reg9, raw_reg10, raw_reg11, raw_reg12, raw_reg13, raw_reg14, raw_reg15, raw_reg16, raw_reg17, raw_reg18, raw_reg19, raw_reg20, raw_reg21, raw_reg22, raw_reg23, raw_reg24, raw_reg25, raw_reg26, raw_reg27, raw_reg28, raw_reg29, raw_reg30, raw_reg31, raw_reg32, raw_reg33, raw_reg34, raw_reg35, raw_reg36, raw_reg37, raw_reg38, raw_reg39, raw_reg40, raw_reg41, raw_reg42, raw_reg43, raw_reg44, raw_reg45, raw_reg46, raw_reg47, raw_reg48, raw_reg49, raw_reg50, raw_reg51, raw_reg52, raw_reg53, raw_reg54, raw_reg55, raw_reg56, raw_reg57, raw_reg58, raw_reg59, raw_reg60, raw_reg61, raw_reg62, raw_reg63, raw_reg64 }, { _3063_, _3062_, _3061_, _3060_, _3059_, _3058_, _3057_, _3056_, _3055_, _3054_, _3053_, _3052_, _3051_, _3050_, _3049_, _3048_, _3047_, _3046_, _3045_, _3044_, _3043_, _3042_, _3041_, _3040_, _3039_, _3038_, _3037_, _3036_, _3035_, _3034_, _3033_, _3032_, _3031_, _3030_, _3029_, _3028_, _3027_, _3026_, _3025_, _3024_, _3023_, _3022_, _3021_, _3020_, _3019_, _3018_, _3017_, _3016_, _3015_, _3014_, _3013_, _3012_, _3011_, _3010_, _3009_, _3008_, _3007_, _3006_, _3005_, _3004_, _3003_, _3002_, _3001_, _0411_ });
  assign _2999_ = dp2lut_X_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6347|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6090" *) 7'b1000000;
  assign _3000_ = dp2lut_X_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6343|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6090" *) 6'b111111;
  assign _3001_ = dp2lut_X_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6339|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6090" *) 6'b111110;
  assign _3002_ = dp2lut_X_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6335|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6090" *) 6'b111101;
  assign _3003_ = dp2lut_X_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6331|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6090" *) 6'b111100;
  assign _3004_ = dp2lut_X_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6327|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6090" *) 6'b111011;
  assign _3005_ = dp2lut_X_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6323|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6090" *) 6'b111010;
  assign _3006_ = dp2lut_X_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6319|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6090" *) 6'b111001;
  assign _3007_ = dp2lut_X_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6315|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6090" *) 6'b111000;
  assign _3008_ = dp2lut_X_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6311|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6090" *) 6'b110111;
  assign _3009_ = dp2lut_X_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6307|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6090" *) 6'b110110;
  assign _3010_ = dp2lut_X_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6303|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6090" *) 6'b110101;
  assign _3011_ = dp2lut_X_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6299|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6090" *) 6'b110100;
  assign _3012_ = dp2lut_X_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6295|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6090" *) 6'b110011;
  assign _3013_ = dp2lut_X_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6291|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6090" *) 6'b110010;
  assign _3014_ = dp2lut_X_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6287|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6090" *) 6'b110001;
  assign _3015_ = dp2lut_X_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6283|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6090" *) 6'b110000;
  assign _3016_ = dp2lut_X_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6279|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6090" *) 6'b101111;
  assign _3017_ = dp2lut_X_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6275|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6090" *) 6'b101110;
  assign _3018_ = dp2lut_X_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6271|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6090" *) 6'b101101;
  assign _3019_ = dp2lut_X_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6267|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6090" *) 6'b101100;
  assign _3020_ = dp2lut_X_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6263|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6090" *) 6'b101011;
  assign _3021_ = dp2lut_X_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6259|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6090" *) 6'b101010;
  assign _3022_ = dp2lut_X_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6255|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6090" *) 6'b101001;
  assign _3023_ = dp2lut_X_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6251|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6090" *) 6'b101000;
  assign _3024_ = dp2lut_X_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6247|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6090" *) 6'b100111;
  assign _3025_ = dp2lut_X_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6243|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6090" *) 6'b100110;
  assign _3026_ = dp2lut_X_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6239|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6090" *) 6'b100101;
  assign _3027_ = dp2lut_X_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6235|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6090" *) 6'b100100;
  assign _3028_ = dp2lut_X_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6231|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6090" *) 6'b100011;
  assign _3029_ = dp2lut_X_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6227|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6090" *) 6'b100010;
  assign _3030_ = dp2lut_X_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6223|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6090" *) 6'b100001;
  assign _3031_ = dp2lut_X_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6219|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6090" *) 6'b100000;
  assign _3032_ = dp2lut_X_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6215|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6090" *) 5'b11111;
  assign _3033_ = dp2lut_X_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6211|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6090" *) 5'b11110;
  assign _3034_ = dp2lut_X_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6207|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6090" *) 5'b11101;
  assign _3035_ = dp2lut_X_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6203|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6090" *) 5'b11100;
  assign _3036_ = dp2lut_X_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6199|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6090" *) 5'b11011;
  assign _3037_ = dp2lut_X_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6195|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6090" *) 5'b11010;
  assign _3038_ = dp2lut_X_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6191|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6090" *) 5'b11001;
  assign _3039_ = dp2lut_X_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6187|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6090" *) 5'b11000;
  assign _3040_ = dp2lut_X_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6183|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6090" *) 5'b10111;
  assign _3041_ = dp2lut_X_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6179|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6090" *) 5'b10110;
  assign _3042_ = dp2lut_X_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6175|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6090" *) 5'b10101;
  assign _3043_ = dp2lut_X_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6171|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6090" *) 5'b10100;
  assign _3044_ = dp2lut_X_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6167|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6090" *) 5'b10011;
  assign _3045_ = dp2lut_X_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6163|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6090" *) 5'b10010;
  assign _3046_ = dp2lut_X_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6159|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6090" *) 5'b10001;
  assign _3047_ = dp2lut_X_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6155|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6090" *) 5'b10000;
  assign _3048_ = dp2lut_X_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6151|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6090" *) 4'b1111;
  assign _3049_ = dp2lut_X_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6147|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6090" *) 4'b1110;
  assign _3050_ = dp2lut_X_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6143|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6090" *) 4'b1101;
  assign _3051_ = dp2lut_X_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6139|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6090" *) 4'b1100;
  assign _3052_ = dp2lut_X_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6135|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6090" *) 4'b1011;
  assign _3053_ = dp2lut_X_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6131|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6090" *) 4'b1010;
  assign _3054_ = dp2lut_X_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6127|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6090" *) 4'b1001;
  assign _3055_ = dp2lut_X_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6123|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6090" *) 4'b1000;
  assign _3056_ = dp2lut_X_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6119|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6090" *) 3'b111;
  assign _3057_ = dp2lut_X_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6115|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6090" *) 3'b110;
  assign _3058_ = dp2lut_X_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6111|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6090" *) 3'b101;
  assign _3059_ = dp2lut_X_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6107|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6090" *) 3'b100;
  assign _3060_ = dp2lut_X_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6103|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6090" *) 2'b11;
  assign _3061_ = dp2lut_X_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6099|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6090" *) 2'b10;
  assign _3062_ = dp2lut_X_entry_4 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6095|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6090" *) 1'b1;
  assign _3063_ = ! (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6091|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6090" *) dp2lut_X_entry_4;
  assign _3064_ = dp2lut_Xinfo_4[17] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6086" *) raw_reg64 : _2998_;
  assign _3065_ = dp2lut_Xinfo_4[16] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6083" *) raw_reg0 : _3064_;
  assign _0270_ = _0396_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6082" *) _3065_ : lut_X_data_41;
  function [15:0] _6932_;
    input [15:0] a;
    input [1023:0] b;
    input [63:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6347|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6090" *)
    (* parallel_case *)
    casez (s)
      64'b???????????????????????????????????????????????????????????????1:
        _6932_ = b[15:0];
      64'b??????????????????????????????????????????????????????????????1?:
        _6932_ = b[31:16];
      64'b?????????????????????????????????????????????????????????????1??:
        _6932_ = b[47:32];
      64'b????????????????????????????????????????????????????????????1???:
        _6932_ = b[63:48];
      64'b???????????????????????????????????????????????????????????1????:
        _6932_ = b[79:64];
      64'b??????????????????????????????????????????????????????????1?????:
        _6932_ = b[95:80];
      64'b?????????????????????????????????????????????????????????1??????:
        _6932_ = b[111:96];
      64'b????????????????????????????????????????????????????????1???????:
        _6932_ = b[127:112];
      64'b???????????????????????????????????????????????????????1????????:
        _6932_ = b[143:128];
      64'b??????????????????????????????????????????????????????1?????????:
        _6932_ = b[159:144];
      64'b?????????????????????????????????????????????????????1??????????:
        _6932_ = b[175:160];
      64'b????????????????????????????????????????????????????1???????????:
        _6932_ = b[191:176];
      64'b???????????????????????????????????????????????????1????????????:
        _6932_ = b[207:192];
      64'b??????????????????????????????????????????????????1?????????????:
        _6932_ = b[223:208];
      64'b?????????????????????????????????????????????????1??????????????:
        _6932_ = b[239:224];
      64'b????????????????????????????????????????????????1???????????????:
        _6932_ = b[255:240];
      64'b???????????????????????????????????????????????1????????????????:
        _6932_ = b[271:256];
      64'b??????????????????????????????????????????????1?????????????????:
        _6932_ = b[287:272];
      64'b?????????????????????????????????????????????1??????????????????:
        _6932_ = b[303:288];
      64'b????????????????????????????????????????????1???????????????????:
        _6932_ = b[319:304];
      64'b???????????????????????????????????????????1????????????????????:
        _6932_ = b[335:320];
      64'b??????????????????????????????????????????1?????????????????????:
        _6932_ = b[351:336];
      64'b?????????????????????????????????????????1??????????????????????:
        _6932_ = b[367:352];
      64'b????????????????????????????????????????1???????????????????????:
        _6932_ = b[383:368];
      64'b???????????????????????????????????????1????????????????????????:
        _6932_ = b[399:384];
      64'b??????????????????????????????????????1?????????????????????????:
        _6932_ = b[415:400];
      64'b?????????????????????????????????????1??????????????????????????:
        _6932_ = b[431:416];
      64'b????????????????????????????????????1???????????????????????????:
        _6932_ = b[447:432];
      64'b???????????????????????????????????1????????????????????????????:
        _6932_ = b[463:448];
      64'b??????????????????????????????????1?????????????????????????????:
        _6932_ = b[479:464];
      64'b?????????????????????????????????1??????????????????????????????:
        _6932_ = b[495:480];
      64'b????????????????????????????????1???????????????????????????????:
        _6932_ = b[511:496];
      64'b???????????????????????????????1????????????????????????????????:
        _6932_ = b[527:512];
      64'b??????????????????????????????1?????????????????????????????????:
        _6932_ = b[543:528];
      64'b?????????????????????????????1??????????????????????????????????:
        _6932_ = b[559:544];
      64'b????????????????????????????1???????????????????????????????????:
        _6932_ = b[575:560];
      64'b???????????????????????????1????????????????????????????????????:
        _6932_ = b[591:576];
      64'b??????????????????????????1?????????????????????????????????????:
        _6932_ = b[607:592];
      64'b?????????????????????????1??????????????????????????????????????:
        _6932_ = b[623:608];
      64'b????????????????????????1???????????????????????????????????????:
        _6932_ = b[639:624];
      64'b???????????????????????1????????????????????????????????????????:
        _6932_ = b[655:640];
      64'b??????????????????????1?????????????????????????????????????????:
        _6932_ = b[671:656];
      64'b?????????????????????1??????????????????????????????????????????:
        _6932_ = b[687:672];
      64'b????????????????????1???????????????????????????????????????????:
        _6932_ = b[703:688];
      64'b???????????????????1????????????????????????????????????????????:
        _6932_ = b[719:704];
      64'b??????????????????1?????????????????????????????????????????????:
        _6932_ = b[735:720];
      64'b?????????????????1??????????????????????????????????????????????:
        _6932_ = b[751:736];
      64'b????????????????1???????????????????????????????????????????????:
        _6932_ = b[767:752];
      64'b???????????????1????????????????????????????????????????????????:
        _6932_ = b[783:768];
      64'b??????????????1?????????????????????????????????????????????????:
        _6932_ = b[799:784];
      64'b?????????????1??????????????????????????????????????????????????:
        _6932_ = b[815:800];
      64'b????????????1???????????????????????????????????????????????????:
        _6932_ = b[831:816];
      64'b???????????1????????????????????????????????????????????????????:
        _6932_ = b[847:832];
      64'b??????????1?????????????????????????????????????????????????????:
        _6932_ = b[863:848];
      64'b?????????1??????????????????????????????????????????????????????:
        _6932_ = b[879:864];
      64'b????????1???????????????????????????????????????????????????????:
        _6932_ = b[895:880];
      64'b???????1????????????????????????????????????????????????????????:
        _6932_ = b[911:896];
      64'b??????1?????????????????????????????????????????????????????????:
        _6932_ = b[927:912];
      64'b?????1??????????????????????????????????????????????????????????:
        _6932_ = b[943:928];
      64'b????1???????????????????????????????????????????????????????????:
        _6932_ = b[959:944];
      64'b???1????????????????????????????????????????????????????????????:
        _6932_ = b[975:960];
      64'b??1?????????????????????????????????????????????????????????????:
        _6932_ = b[991:976];
      64'b?1??????????????????????????????????????????????????????????????:
        _6932_ = b[1007:992];
      64'b1???????????????????????????????????????????????????????????????:
        _6932_ = b[1023:1008];
      default:
        _6932_ = a;
    endcase
  endfunction
  assign _3066_ = _6932_(raw_reg0, { raw_reg1, raw_reg2, raw_reg3, raw_reg4, raw_reg5, raw_reg6, raw_reg7, raw_reg8, raw_reg9, raw_reg10, raw_reg11, raw_reg12, raw_reg13, raw_reg14, raw_reg15, raw_reg16, raw_reg17, raw_reg18, raw_reg19, raw_reg20, raw_reg21, raw_reg22, raw_reg23, raw_reg24, raw_reg25, raw_reg26, raw_reg27, raw_reg28, raw_reg29, raw_reg30, raw_reg31, raw_reg32, raw_reg33, raw_reg34, raw_reg35, raw_reg36, raw_reg37, raw_reg38, raw_reg39, raw_reg40, raw_reg41, raw_reg42, raw_reg43, raw_reg44, raw_reg45, raw_reg46, raw_reg47, raw_reg48, raw_reg49, raw_reg50, raw_reg51, raw_reg52, raw_reg53, raw_reg54, raw_reg55, raw_reg56, raw_reg57, raw_reg58, raw_reg59, raw_reg60, raw_reg61, raw_reg62, raw_reg63, raw_reg64 }, { _3062_, _3061_, _3060_, _3059_, _3058_, _3057_, _3056_, _3055_, _3054_, _3053_, _3052_, _3051_, _3050_, _3049_, _3048_, _3047_, _3046_, _3045_, _3044_, _3043_, _3042_, _3041_, _3040_, _3039_, _3038_, _3037_, _3036_, _3035_, _3034_, _3033_, _3032_, _3031_, _3030_, _3029_, _3028_, _3027_, _3026_, _3025_, _3024_, _3023_, _3022_, _3021_, _3020_, _3019_, _3018_, _3017_, _3016_, _3015_, _3014_, _3013_, _3012_, _3011_, _3010_, _3009_, _3008_, _3007_, _3006_, _3005_, _3004_, _3003_, _3002_, _3001_, _3000_, _2999_ });
  assign _3067_ = dp2lut_Xinfo_4[17] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6086" *) raw_reg64 : _3066_;
  assign _3068_ = dp2lut_Xinfo_4[16] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6083" *) raw_reg0 : _3067_;
  assign _0269_ = _0396_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6082" *) _3068_ : lut_X_data_40;
  function [15:0] _6936_;
    input [15:0] a;
    input [1023:0] b;
    input [63:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6064|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5807" *)
    (* parallel_case *)
    casez (s)
      64'b???????????????????????????????????????????????????????????????1:
        _6936_ = b[15:0];
      64'b??????????????????????????????????????????????????????????????1?:
        _6936_ = b[31:16];
      64'b?????????????????????????????????????????????????????????????1??:
        _6936_ = b[47:32];
      64'b????????????????????????????????????????????????????????????1???:
        _6936_ = b[63:48];
      64'b???????????????????????????????????????????????????????????1????:
        _6936_ = b[79:64];
      64'b??????????????????????????????????????????????????????????1?????:
        _6936_ = b[95:80];
      64'b?????????????????????????????????????????????????????????1??????:
        _6936_ = b[111:96];
      64'b????????????????????????????????????????????????????????1???????:
        _6936_ = b[127:112];
      64'b???????????????????????????????????????????????????????1????????:
        _6936_ = b[143:128];
      64'b??????????????????????????????????????????????????????1?????????:
        _6936_ = b[159:144];
      64'b?????????????????????????????????????????????????????1??????????:
        _6936_ = b[175:160];
      64'b????????????????????????????????????????????????????1???????????:
        _6936_ = b[191:176];
      64'b???????????????????????????????????????????????????1????????????:
        _6936_ = b[207:192];
      64'b??????????????????????????????????????????????????1?????????????:
        _6936_ = b[223:208];
      64'b?????????????????????????????????????????????????1??????????????:
        _6936_ = b[239:224];
      64'b????????????????????????????????????????????????1???????????????:
        _6936_ = b[255:240];
      64'b???????????????????????????????????????????????1????????????????:
        _6936_ = b[271:256];
      64'b??????????????????????????????????????????????1?????????????????:
        _6936_ = b[287:272];
      64'b?????????????????????????????????????????????1??????????????????:
        _6936_ = b[303:288];
      64'b????????????????????????????????????????????1???????????????????:
        _6936_ = b[319:304];
      64'b???????????????????????????????????????????1????????????????????:
        _6936_ = b[335:320];
      64'b??????????????????????????????????????????1?????????????????????:
        _6936_ = b[351:336];
      64'b?????????????????????????????????????????1??????????????????????:
        _6936_ = b[367:352];
      64'b????????????????????????????????????????1???????????????????????:
        _6936_ = b[383:368];
      64'b???????????????????????????????????????1????????????????????????:
        _6936_ = b[399:384];
      64'b??????????????????????????????????????1?????????????????????????:
        _6936_ = b[415:400];
      64'b?????????????????????????????????????1??????????????????????????:
        _6936_ = b[431:416];
      64'b????????????????????????????????????1???????????????????????????:
        _6936_ = b[447:432];
      64'b???????????????????????????????????1????????????????????????????:
        _6936_ = b[463:448];
      64'b??????????????????????????????????1?????????????????????????????:
        _6936_ = b[479:464];
      64'b?????????????????????????????????1??????????????????????????????:
        _6936_ = b[495:480];
      64'b????????????????????????????????1???????????????????????????????:
        _6936_ = b[511:496];
      64'b???????????????????????????????1????????????????????????????????:
        _6936_ = b[527:512];
      64'b??????????????????????????????1?????????????????????????????????:
        _6936_ = b[543:528];
      64'b?????????????????????????????1??????????????????????????????????:
        _6936_ = b[559:544];
      64'b????????????????????????????1???????????????????????????????????:
        _6936_ = b[575:560];
      64'b???????????????????????????1????????????????????????????????????:
        _6936_ = b[591:576];
      64'b??????????????????????????1?????????????????????????????????????:
        _6936_ = b[607:592];
      64'b?????????????????????????1??????????????????????????????????????:
        _6936_ = b[623:608];
      64'b????????????????????????1???????????????????????????????????????:
        _6936_ = b[639:624];
      64'b???????????????????????1????????????????????????????????????????:
        _6936_ = b[655:640];
      64'b??????????????????????1?????????????????????????????????????????:
        _6936_ = b[671:656];
      64'b?????????????????????1??????????????????????????????????????????:
        _6936_ = b[687:672];
      64'b????????????????????1???????????????????????????????????????????:
        _6936_ = b[703:688];
      64'b???????????????????1????????????????????????????????????????????:
        _6936_ = b[719:704];
      64'b??????????????????1?????????????????????????????????????????????:
        _6936_ = b[735:720];
      64'b?????????????????1??????????????????????????????????????????????:
        _6936_ = b[751:736];
      64'b????????????????1???????????????????????????????????????????????:
        _6936_ = b[767:752];
      64'b???????????????1????????????????????????????????????????????????:
        _6936_ = b[783:768];
      64'b??????????????1?????????????????????????????????????????????????:
        _6936_ = b[799:784];
      64'b?????????????1??????????????????????????????????????????????????:
        _6936_ = b[815:800];
      64'b????????????1???????????????????????????????????????????????????:
        _6936_ = b[831:816];
      64'b???????????1????????????????????????????????????????????????????:
        _6936_ = b[847:832];
      64'b??????????1?????????????????????????????????????????????????????:
        _6936_ = b[863:848];
      64'b?????????1??????????????????????????????????????????????????????:
        _6936_ = b[879:864];
      64'b????????1???????????????????????????????????????????????????????:
        _6936_ = b[895:880];
      64'b???????1????????????????????????????????????????????????????????:
        _6936_ = b[911:896];
      64'b??????1?????????????????????????????????????????????????????????:
        _6936_ = b[927:912];
      64'b?????1??????????????????????????????????????????????????????????:
        _6936_ = b[943:928];
      64'b????1???????????????????????????????????????????????????????????:
        _6936_ = b[959:944];
      64'b???1????????????????????????????????????????????????????????????:
        _6936_ = b[975:960];
      64'b??1?????????????????????????????????????????????????????????????:
        _6936_ = b[991:976];
      64'b?1??????????????????????????????????????????????????????????????:
        _6936_ = b[1007:992];
      64'b1???????????????????????????????????????????????????????????????:
        _6936_ = b[1023:1008];
      default:
        _6936_ = a;
    endcase
  endfunction
  assign _3069_ = _6936_(raw_reg0, { raw_reg1, raw_reg2, raw_reg3, raw_reg4, raw_reg5, raw_reg6, raw_reg7, raw_reg8, raw_reg9, raw_reg10, raw_reg11, raw_reg12, raw_reg13, raw_reg14, raw_reg15, raw_reg16, raw_reg17, raw_reg18, raw_reg19, raw_reg20, raw_reg21, raw_reg22, raw_reg23, raw_reg24, raw_reg25, raw_reg26, raw_reg27, raw_reg28, raw_reg29, raw_reg30, raw_reg31, raw_reg32, raw_reg33, raw_reg34, raw_reg35, raw_reg36, raw_reg37, raw_reg38, raw_reg39, raw_reg40, raw_reg41, raw_reg42, raw_reg43, raw_reg44, raw_reg45, raw_reg46, raw_reg47, raw_reg48, raw_reg49, raw_reg50, raw_reg51, raw_reg52, raw_reg53, raw_reg54, raw_reg55, raw_reg56, raw_reg57, raw_reg58, raw_reg59, raw_reg60, raw_reg61, raw_reg62, raw_reg63, raw_reg64 }, { _3134_, _3133_, _3132_, _3131_, _3130_, _3129_, _3128_, _3127_, _3126_, _3125_, _3124_, _3123_, _3122_, _3121_, _3120_, _3119_, _3118_, _3117_, _3116_, _3115_, _3114_, _3113_, _3112_, _3111_, _3110_, _3109_, _3108_, _3107_, _3106_, _3105_, _3104_, _3103_, _3102_, _3101_, _3100_, _3099_, _3098_, _3097_, _3096_, _3095_, _3094_, _3093_, _3092_, _3091_, _3090_, _3089_, _3088_, _3087_, _3086_, _3085_, _3084_, _3083_, _3082_, _3081_, _3080_, _3079_, _3078_, _3077_, _3076_, _3075_, _3074_, _3073_, _3072_, _0413_ });
  assign _3070_ = dp2lut_X_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6064|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5807" *) 7'b1000000;
  assign _3071_ = dp2lut_X_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6060|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5807" *) 6'b111111;
  assign _3072_ = dp2lut_X_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6056|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5807" *) 6'b111110;
  assign _3073_ = dp2lut_X_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6052|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5807" *) 6'b111101;
  assign _3074_ = dp2lut_X_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6048|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5807" *) 6'b111100;
  assign _3075_ = dp2lut_X_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6044|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5807" *) 6'b111011;
  assign _3076_ = dp2lut_X_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6040|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5807" *) 6'b111010;
  assign _3077_ = dp2lut_X_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6036|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5807" *) 6'b111001;
  assign _3078_ = dp2lut_X_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6032|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5807" *) 6'b111000;
  assign _3079_ = dp2lut_X_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6028|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5807" *) 6'b110111;
  assign _3080_ = dp2lut_X_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6024|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5807" *) 6'b110110;
  assign _3081_ = dp2lut_X_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6020|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5807" *) 6'b110101;
  assign _3082_ = dp2lut_X_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6016|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5807" *) 6'b110100;
  assign _3083_ = dp2lut_X_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6012|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5807" *) 6'b110011;
  assign _3084_ = dp2lut_X_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6008|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5807" *) 6'b110010;
  assign _3085_ = dp2lut_X_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6004|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5807" *) 6'b110001;
  assign _3086_ = dp2lut_X_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6000|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5807" *) 6'b110000;
  assign _3087_ = dp2lut_X_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5996|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5807" *) 6'b101111;
  assign _3088_ = dp2lut_X_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5992|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5807" *) 6'b101110;
  assign _3089_ = dp2lut_X_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5988|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5807" *) 6'b101101;
  assign _3090_ = dp2lut_X_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5984|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5807" *) 6'b101100;
  assign _3091_ = dp2lut_X_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5980|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5807" *) 6'b101011;
  assign _3092_ = dp2lut_X_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5976|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5807" *) 6'b101010;
  assign _3093_ = dp2lut_X_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5972|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5807" *) 6'b101001;
  assign _3094_ = dp2lut_X_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5968|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5807" *) 6'b101000;
  assign _3095_ = dp2lut_X_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5964|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5807" *) 6'b100111;
  assign _3096_ = dp2lut_X_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5960|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5807" *) 6'b100110;
  assign _3097_ = dp2lut_X_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5956|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5807" *) 6'b100101;
  assign _3098_ = dp2lut_X_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5952|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5807" *) 6'b100100;
  assign _3099_ = dp2lut_X_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5948|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5807" *) 6'b100011;
  assign _3100_ = dp2lut_X_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5944|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5807" *) 6'b100010;
  assign _3101_ = dp2lut_X_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5940|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5807" *) 6'b100001;
  assign _3102_ = dp2lut_X_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5936|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5807" *) 6'b100000;
  assign _3103_ = dp2lut_X_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5932|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5807" *) 5'b11111;
  assign _3104_ = dp2lut_X_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5928|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5807" *) 5'b11110;
  assign _3105_ = dp2lut_X_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5924|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5807" *) 5'b11101;
  assign _3106_ = dp2lut_X_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5920|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5807" *) 5'b11100;
  assign _3107_ = dp2lut_X_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5916|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5807" *) 5'b11011;
  assign _3108_ = dp2lut_X_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5912|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5807" *) 5'b11010;
  assign _3109_ = dp2lut_X_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5908|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5807" *) 5'b11001;
  assign _3110_ = dp2lut_X_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5904|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5807" *) 5'b11000;
  assign _3111_ = dp2lut_X_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5900|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5807" *) 5'b10111;
  assign _3112_ = dp2lut_X_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5896|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5807" *) 5'b10110;
  assign _3113_ = dp2lut_X_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5892|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5807" *) 5'b10101;
  assign _3114_ = dp2lut_X_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5888|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5807" *) 5'b10100;
  assign _3115_ = dp2lut_X_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5884|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5807" *) 5'b10011;
  assign _3116_ = dp2lut_X_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5880|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5807" *) 5'b10010;
  assign _3117_ = dp2lut_X_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5876|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5807" *) 5'b10001;
  assign _3118_ = dp2lut_X_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5872|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5807" *) 5'b10000;
  assign _3119_ = dp2lut_X_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5868|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5807" *) 4'b1111;
  assign _3120_ = dp2lut_X_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5864|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5807" *) 4'b1110;
  assign _3121_ = dp2lut_X_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5860|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5807" *) 4'b1101;
  assign _3122_ = dp2lut_X_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5856|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5807" *) 4'b1100;
  assign _3123_ = dp2lut_X_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5852|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5807" *) 4'b1011;
  assign _3124_ = dp2lut_X_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5848|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5807" *) 4'b1010;
  assign _3125_ = dp2lut_X_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5844|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5807" *) 4'b1001;
  assign _3126_ = dp2lut_X_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5840|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5807" *) 4'b1000;
  assign _3127_ = dp2lut_X_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5836|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5807" *) 3'b111;
  assign _3128_ = dp2lut_X_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5832|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5807" *) 3'b110;
  assign _3129_ = dp2lut_X_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5828|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5807" *) 3'b101;
  assign _3130_ = dp2lut_X_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5824|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5807" *) 3'b100;
  assign _3131_ = dp2lut_X_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5820|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5807" *) 2'b11;
  assign _3132_ = dp2lut_X_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5816|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5807" *) 2'b10;
  assign _3133_ = dp2lut_X_entry_3 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5812|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5807" *) 1'b1;
  assign _3134_ = ! (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5808|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5807" *) dp2lut_X_entry_3;
  assign _3135_ = dp2lut_Xinfo_3[17] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5803" *) raw_reg64 : _3069_;
  assign _3136_ = dp2lut_Xinfo_3[16] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5800" *) raw_reg0 : _3135_;
  assign _0268_ = _0395_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5799" *) _3136_ : lut_X_data_31;
  function [15:0] _7005_;
    input [15:0] a;
    input [1023:0] b;
    input [63:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:6064|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5807" *)
    (* parallel_case *)
    casez (s)
      64'b???????????????????????????????????????????????????????????????1:
        _7005_ = b[15:0];
      64'b??????????????????????????????????????????????????????????????1?:
        _7005_ = b[31:16];
      64'b?????????????????????????????????????????????????????????????1??:
        _7005_ = b[47:32];
      64'b????????????????????????????????????????????????????????????1???:
        _7005_ = b[63:48];
      64'b???????????????????????????????????????????????????????????1????:
        _7005_ = b[79:64];
      64'b??????????????????????????????????????????????????????????1?????:
        _7005_ = b[95:80];
      64'b?????????????????????????????????????????????????????????1??????:
        _7005_ = b[111:96];
      64'b????????????????????????????????????????????????????????1???????:
        _7005_ = b[127:112];
      64'b???????????????????????????????????????????????????????1????????:
        _7005_ = b[143:128];
      64'b??????????????????????????????????????????????????????1?????????:
        _7005_ = b[159:144];
      64'b?????????????????????????????????????????????????????1??????????:
        _7005_ = b[175:160];
      64'b????????????????????????????????????????????????????1???????????:
        _7005_ = b[191:176];
      64'b???????????????????????????????????????????????????1????????????:
        _7005_ = b[207:192];
      64'b??????????????????????????????????????????????????1?????????????:
        _7005_ = b[223:208];
      64'b?????????????????????????????????????????????????1??????????????:
        _7005_ = b[239:224];
      64'b????????????????????????????????????????????????1???????????????:
        _7005_ = b[255:240];
      64'b???????????????????????????????????????????????1????????????????:
        _7005_ = b[271:256];
      64'b??????????????????????????????????????????????1?????????????????:
        _7005_ = b[287:272];
      64'b?????????????????????????????????????????????1??????????????????:
        _7005_ = b[303:288];
      64'b????????????????????????????????????????????1???????????????????:
        _7005_ = b[319:304];
      64'b???????????????????????????????????????????1????????????????????:
        _7005_ = b[335:320];
      64'b??????????????????????????????????????????1?????????????????????:
        _7005_ = b[351:336];
      64'b?????????????????????????????????????????1??????????????????????:
        _7005_ = b[367:352];
      64'b????????????????????????????????????????1???????????????????????:
        _7005_ = b[383:368];
      64'b???????????????????????????????????????1????????????????????????:
        _7005_ = b[399:384];
      64'b??????????????????????????????????????1?????????????????????????:
        _7005_ = b[415:400];
      64'b?????????????????????????????????????1??????????????????????????:
        _7005_ = b[431:416];
      64'b????????????????????????????????????1???????????????????????????:
        _7005_ = b[447:432];
      64'b???????????????????????????????????1????????????????????????????:
        _7005_ = b[463:448];
      64'b??????????????????????????????????1?????????????????????????????:
        _7005_ = b[479:464];
      64'b?????????????????????????????????1??????????????????????????????:
        _7005_ = b[495:480];
      64'b????????????????????????????????1???????????????????????????????:
        _7005_ = b[511:496];
      64'b???????????????????????????????1????????????????????????????????:
        _7005_ = b[527:512];
      64'b??????????????????????????????1?????????????????????????????????:
        _7005_ = b[543:528];
      64'b?????????????????????????????1??????????????????????????????????:
        _7005_ = b[559:544];
      64'b????????????????????????????1???????????????????????????????????:
        _7005_ = b[575:560];
      64'b???????????????????????????1????????????????????????????????????:
        _7005_ = b[591:576];
      64'b??????????????????????????1?????????????????????????????????????:
        _7005_ = b[607:592];
      64'b?????????????????????????1??????????????????????????????????????:
        _7005_ = b[623:608];
      64'b????????????????????????1???????????????????????????????????????:
        _7005_ = b[639:624];
      64'b???????????????????????1????????????????????????????????????????:
        _7005_ = b[655:640];
      64'b??????????????????????1?????????????????????????????????????????:
        _7005_ = b[671:656];
      64'b?????????????????????1??????????????????????????????????????????:
        _7005_ = b[687:672];
      64'b????????????????????1???????????????????????????????????????????:
        _7005_ = b[703:688];
      64'b???????????????????1????????????????????????????????????????????:
        _7005_ = b[719:704];
      64'b??????????????????1?????????????????????????????????????????????:
        _7005_ = b[735:720];
      64'b?????????????????1??????????????????????????????????????????????:
        _7005_ = b[751:736];
      64'b????????????????1???????????????????????????????????????????????:
        _7005_ = b[767:752];
      64'b???????????????1????????????????????????????????????????????????:
        _7005_ = b[783:768];
      64'b??????????????1?????????????????????????????????????????????????:
        _7005_ = b[799:784];
      64'b?????????????1??????????????????????????????????????????????????:
        _7005_ = b[815:800];
      64'b????????????1???????????????????????????????????????????????????:
        _7005_ = b[831:816];
      64'b???????????1????????????????????????????????????????????????????:
        _7005_ = b[847:832];
      64'b??????????1?????????????????????????????????????????????????????:
        _7005_ = b[863:848];
      64'b?????????1??????????????????????????????????????????????????????:
        _7005_ = b[879:864];
      64'b????????1???????????????????????????????????????????????????????:
        _7005_ = b[895:880];
      64'b???????1????????????????????????????????????????????????????????:
        _7005_ = b[911:896];
      64'b??????1?????????????????????????????????????????????????????????:
        _7005_ = b[927:912];
      64'b?????1??????????????????????????????????????????????????????????:
        _7005_ = b[943:928];
      64'b????1???????????????????????????????????????????????????????????:
        _7005_ = b[959:944];
      64'b???1????????????????????????????????????????????????????????????:
        _7005_ = b[975:960];
      64'b??1?????????????????????????????????????????????????????????????:
        _7005_ = b[991:976];
      64'b?1??????????????????????????????????????????????????????????????:
        _7005_ = b[1007:992];
      64'b1???????????????????????????????????????????????????????????????:
        _7005_ = b[1023:1008];
      default:
        _7005_ = a;
    endcase
  endfunction
  assign _3137_ = _7005_(raw_reg0, { raw_reg1, raw_reg2, raw_reg3, raw_reg4, raw_reg5, raw_reg6, raw_reg7, raw_reg8, raw_reg9, raw_reg10, raw_reg11, raw_reg12, raw_reg13, raw_reg14, raw_reg15, raw_reg16, raw_reg17, raw_reg18, raw_reg19, raw_reg20, raw_reg21, raw_reg22, raw_reg23, raw_reg24, raw_reg25, raw_reg26, raw_reg27, raw_reg28, raw_reg29, raw_reg30, raw_reg31, raw_reg32, raw_reg33, raw_reg34, raw_reg35, raw_reg36, raw_reg37, raw_reg38, raw_reg39, raw_reg40, raw_reg41, raw_reg42, raw_reg43, raw_reg44, raw_reg45, raw_reg46, raw_reg47, raw_reg48, raw_reg49, raw_reg50, raw_reg51, raw_reg52, raw_reg53, raw_reg54, raw_reg55, raw_reg56, raw_reg57, raw_reg58, raw_reg59, raw_reg60, raw_reg61, raw_reg62, raw_reg63, raw_reg64 }, { _3133_, _3132_, _3131_, _3130_, _3129_, _3128_, _3127_, _3126_, _3125_, _3124_, _3123_, _3122_, _3121_, _3120_, _3119_, _3118_, _3117_, _3116_, _3115_, _3114_, _3113_, _3112_, _3111_, _3110_, _3109_, _3108_, _3107_, _3106_, _3105_, _3104_, _3103_, _3102_, _3101_, _3100_, _3099_, _3098_, _3097_, _3096_, _3095_, _3094_, _3093_, _3092_, _3091_, _3090_, _3089_, _3088_, _3087_, _3086_, _3085_, _3084_, _3083_, _3082_, _3081_, _3080_, _3079_, _3078_, _3077_, _3076_, _3075_, _3074_, _3073_, _3072_, _3071_, _3070_ });
  assign _3138_ = dp2lut_Xinfo_3[17] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5803" *) raw_reg64 : _3137_;
  assign _3139_ = dp2lut_Xinfo_3[16] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5800" *) raw_reg0 : _3138_;
  assign _0267_ = _0395_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5799" *) _3139_ : lut_X_data_30;
  function [15:0] _7009_;
    input [15:0] a;
    input [1023:0] b;
    input [63:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5781|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5524" *)
    (* parallel_case *)
    casez (s)
      64'b???????????????????????????????????????????????????????????????1:
        _7009_ = b[15:0];
      64'b??????????????????????????????????????????????????????????????1?:
        _7009_ = b[31:16];
      64'b?????????????????????????????????????????????????????????????1??:
        _7009_ = b[47:32];
      64'b????????????????????????????????????????????????????????????1???:
        _7009_ = b[63:48];
      64'b???????????????????????????????????????????????????????????1????:
        _7009_ = b[79:64];
      64'b??????????????????????????????????????????????????????????1?????:
        _7009_ = b[95:80];
      64'b?????????????????????????????????????????????????????????1??????:
        _7009_ = b[111:96];
      64'b????????????????????????????????????????????????????????1???????:
        _7009_ = b[127:112];
      64'b???????????????????????????????????????????????????????1????????:
        _7009_ = b[143:128];
      64'b??????????????????????????????????????????????????????1?????????:
        _7009_ = b[159:144];
      64'b?????????????????????????????????????????????????????1??????????:
        _7009_ = b[175:160];
      64'b????????????????????????????????????????????????????1???????????:
        _7009_ = b[191:176];
      64'b???????????????????????????????????????????????????1????????????:
        _7009_ = b[207:192];
      64'b??????????????????????????????????????????????????1?????????????:
        _7009_ = b[223:208];
      64'b?????????????????????????????????????????????????1??????????????:
        _7009_ = b[239:224];
      64'b????????????????????????????????????????????????1???????????????:
        _7009_ = b[255:240];
      64'b???????????????????????????????????????????????1????????????????:
        _7009_ = b[271:256];
      64'b??????????????????????????????????????????????1?????????????????:
        _7009_ = b[287:272];
      64'b?????????????????????????????????????????????1??????????????????:
        _7009_ = b[303:288];
      64'b????????????????????????????????????????????1???????????????????:
        _7009_ = b[319:304];
      64'b???????????????????????????????????????????1????????????????????:
        _7009_ = b[335:320];
      64'b??????????????????????????????????????????1?????????????????????:
        _7009_ = b[351:336];
      64'b?????????????????????????????????????????1??????????????????????:
        _7009_ = b[367:352];
      64'b????????????????????????????????????????1???????????????????????:
        _7009_ = b[383:368];
      64'b???????????????????????????????????????1????????????????????????:
        _7009_ = b[399:384];
      64'b??????????????????????????????????????1?????????????????????????:
        _7009_ = b[415:400];
      64'b?????????????????????????????????????1??????????????????????????:
        _7009_ = b[431:416];
      64'b????????????????????????????????????1???????????????????????????:
        _7009_ = b[447:432];
      64'b???????????????????????????????????1????????????????????????????:
        _7009_ = b[463:448];
      64'b??????????????????????????????????1?????????????????????????????:
        _7009_ = b[479:464];
      64'b?????????????????????????????????1??????????????????????????????:
        _7009_ = b[495:480];
      64'b????????????????????????????????1???????????????????????????????:
        _7009_ = b[511:496];
      64'b???????????????????????????????1????????????????????????????????:
        _7009_ = b[527:512];
      64'b??????????????????????????????1?????????????????????????????????:
        _7009_ = b[543:528];
      64'b?????????????????????????????1??????????????????????????????????:
        _7009_ = b[559:544];
      64'b????????????????????????????1???????????????????????????????????:
        _7009_ = b[575:560];
      64'b???????????????????????????1????????????????????????????????????:
        _7009_ = b[591:576];
      64'b??????????????????????????1?????????????????????????????????????:
        _7009_ = b[607:592];
      64'b?????????????????????????1??????????????????????????????????????:
        _7009_ = b[623:608];
      64'b????????????????????????1???????????????????????????????????????:
        _7009_ = b[639:624];
      64'b???????????????????????1????????????????????????????????????????:
        _7009_ = b[655:640];
      64'b??????????????????????1?????????????????????????????????????????:
        _7009_ = b[671:656];
      64'b?????????????????????1??????????????????????????????????????????:
        _7009_ = b[687:672];
      64'b????????????????????1???????????????????????????????????????????:
        _7009_ = b[703:688];
      64'b???????????????????1????????????????????????????????????????????:
        _7009_ = b[719:704];
      64'b??????????????????1?????????????????????????????????????????????:
        _7009_ = b[735:720];
      64'b?????????????????1??????????????????????????????????????????????:
        _7009_ = b[751:736];
      64'b????????????????1???????????????????????????????????????????????:
        _7009_ = b[767:752];
      64'b???????????????1????????????????????????????????????????????????:
        _7009_ = b[783:768];
      64'b??????????????1?????????????????????????????????????????????????:
        _7009_ = b[799:784];
      64'b?????????????1??????????????????????????????????????????????????:
        _7009_ = b[815:800];
      64'b????????????1???????????????????????????????????????????????????:
        _7009_ = b[831:816];
      64'b???????????1????????????????????????????????????????????????????:
        _7009_ = b[847:832];
      64'b??????????1?????????????????????????????????????????????????????:
        _7009_ = b[863:848];
      64'b?????????1??????????????????????????????????????????????????????:
        _7009_ = b[879:864];
      64'b????????1???????????????????????????????????????????????????????:
        _7009_ = b[895:880];
      64'b???????1????????????????????????????????????????????????????????:
        _7009_ = b[911:896];
      64'b??????1?????????????????????????????????????????????????????????:
        _7009_ = b[927:912];
      64'b?????1??????????????????????????????????????????????????????????:
        _7009_ = b[943:928];
      64'b????1???????????????????????????????????????????????????????????:
        _7009_ = b[959:944];
      64'b???1????????????????????????????????????????????????????????????:
        _7009_ = b[975:960];
      64'b??1?????????????????????????????????????????????????????????????:
        _7009_ = b[991:976];
      64'b?1??????????????????????????????????????????????????????????????:
        _7009_ = b[1007:992];
      64'b1???????????????????????????????????????????????????????????????:
        _7009_ = b[1023:1008];
      default:
        _7009_ = a;
    endcase
  endfunction
  assign _3140_ = _7009_(raw_reg0, { raw_reg1, raw_reg2, raw_reg3, raw_reg4, raw_reg5, raw_reg6, raw_reg7, raw_reg8, raw_reg9, raw_reg10, raw_reg11, raw_reg12, raw_reg13, raw_reg14, raw_reg15, raw_reg16, raw_reg17, raw_reg18, raw_reg19, raw_reg20, raw_reg21, raw_reg22, raw_reg23, raw_reg24, raw_reg25, raw_reg26, raw_reg27, raw_reg28, raw_reg29, raw_reg30, raw_reg31, raw_reg32, raw_reg33, raw_reg34, raw_reg35, raw_reg36, raw_reg37, raw_reg38, raw_reg39, raw_reg40, raw_reg41, raw_reg42, raw_reg43, raw_reg44, raw_reg45, raw_reg46, raw_reg47, raw_reg48, raw_reg49, raw_reg50, raw_reg51, raw_reg52, raw_reg53, raw_reg54, raw_reg55, raw_reg56, raw_reg57, raw_reg58, raw_reg59, raw_reg60, raw_reg61, raw_reg62, raw_reg63, raw_reg64 }, { _3205_, _3204_, _3203_, _3202_, _3201_, _3200_, _3199_, _3198_, _3197_, _3196_, _3195_, _3194_, _3193_, _3192_, _3191_, _3190_, _3189_, _3188_, _3187_, _3186_, _3185_, _3184_, _3183_, _3182_, _3181_, _3180_, _3179_, _3178_, _3177_, _3176_, _3175_, _3174_, _3173_, _3172_, _3171_, _3170_, _3169_, _3168_, _3167_, _3166_, _3165_, _3164_, _3163_, _3162_, _3161_, _3160_, _3159_, _3158_, _3157_, _3156_, _3155_, _3154_, _3153_, _3152_, _3151_, _3150_, _3149_, _3148_, _3147_, _3146_, _3145_, _3144_, _3143_, _0415_ });
  assign _3141_ = dp2lut_X_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5781|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5524" *) 7'b1000000;
  assign _3142_ = dp2lut_X_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5777|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5524" *) 6'b111111;
  assign _3143_ = dp2lut_X_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5773|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5524" *) 6'b111110;
  assign _3144_ = dp2lut_X_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5769|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5524" *) 6'b111101;
  assign _3145_ = dp2lut_X_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5765|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5524" *) 6'b111100;
  assign _3146_ = dp2lut_X_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5761|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5524" *) 6'b111011;
  assign _3147_ = dp2lut_X_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5757|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5524" *) 6'b111010;
  assign _3148_ = dp2lut_X_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5753|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5524" *) 6'b111001;
  assign _3149_ = dp2lut_X_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5749|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5524" *) 6'b111000;
  assign _3150_ = dp2lut_X_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5745|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5524" *) 6'b110111;
  assign _3151_ = dp2lut_X_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5741|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5524" *) 6'b110110;
  assign _3152_ = dp2lut_X_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5737|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5524" *) 6'b110101;
  assign _3153_ = dp2lut_X_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5733|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5524" *) 6'b110100;
  assign _3154_ = dp2lut_X_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5729|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5524" *) 6'b110011;
  assign _3155_ = dp2lut_X_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5725|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5524" *) 6'b110010;
  assign _3156_ = dp2lut_X_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5721|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5524" *) 6'b110001;
  assign _3157_ = dp2lut_X_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5717|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5524" *) 6'b110000;
  assign _3158_ = dp2lut_X_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5713|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5524" *) 6'b101111;
  assign _3159_ = dp2lut_X_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5709|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5524" *) 6'b101110;
  assign _3160_ = dp2lut_X_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5705|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5524" *) 6'b101101;
  assign _3161_ = dp2lut_X_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5701|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5524" *) 6'b101100;
  assign _3162_ = dp2lut_X_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5697|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5524" *) 6'b101011;
  assign _3163_ = dp2lut_X_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5693|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5524" *) 6'b101010;
  assign _3164_ = dp2lut_X_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5689|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5524" *) 6'b101001;
  assign _3165_ = dp2lut_X_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5685|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5524" *) 6'b101000;
  assign _3166_ = dp2lut_X_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5681|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5524" *) 6'b100111;
  assign _3167_ = dp2lut_X_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5677|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5524" *) 6'b100110;
  assign _3168_ = dp2lut_X_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5673|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5524" *) 6'b100101;
  assign _3169_ = dp2lut_X_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5669|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5524" *) 6'b100100;
  assign _3170_ = dp2lut_X_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5665|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5524" *) 6'b100011;
  assign _3171_ = dp2lut_X_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5661|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5524" *) 6'b100010;
  assign _3172_ = dp2lut_X_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5657|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5524" *) 6'b100001;
  assign _3173_ = dp2lut_X_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5653|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5524" *) 6'b100000;
  assign _3174_ = dp2lut_X_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5649|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5524" *) 5'b11111;
  assign _3175_ = dp2lut_X_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5645|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5524" *) 5'b11110;
  assign _3176_ = dp2lut_X_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5641|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5524" *) 5'b11101;
  assign _3177_ = dp2lut_X_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5637|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5524" *) 5'b11100;
  assign _3178_ = dp2lut_X_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5633|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5524" *) 5'b11011;
  assign _3179_ = dp2lut_X_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5629|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5524" *) 5'b11010;
  assign _3180_ = dp2lut_X_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5625|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5524" *) 5'b11001;
  assign _3181_ = dp2lut_X_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5621|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5524" *) 5'b11000;
  assign _3182_ = dp2lut_X_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5617|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5524" *) 5'b10111;
  assign _3183_ = dp2lut_X_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5613|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5524" *) 5'b10110;
  assign _3184_ = dp2lut_X_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5609|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5524" *) 5'b10101;
  assign _3185_ = dp2lut_X_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5605|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5524" *) 5'b10100;
  assign _3186_ = dp2lut_X_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5601|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5524" *) 5'b10011;
  assign _3187_ = dp2lut_X_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5597|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5524" *) 5'b10010;
  assign _3188_ = dp2lut_X_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5593|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5524" *) 5'b10001;
  assign _3189_ = dp2lut_X_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5589|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5524" *) 5'b10000;
  assign _3190_ = dp2lut_X_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5585|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5524" *) 4'b1111;
  assign _3191_ = dp2lut_X_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5581|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5524" *) 4'b1110;
  assign _3192_ = dp2lut_X_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5577|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5524" *) 4'b1101;
  assign _3193_ = dp2lut_X_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5573|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5524" *) 4'b1100;
  assign _3194_ = dp2lut_X_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5569|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5524" *) 4'b1011;
  assign _3195_ = dp2lut_X_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5565|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5524" *) 4'b1010;
  assign _3196_ = dp2lut_X_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5561|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5524" *) 4'b1001;
  assign _3197_ = dp2lut_X_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5557|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5524" *) 4'b1000;
  assign _3198_ = dp2lut_X_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5553|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5524" *) 3'b111;
  assign _3199_ = dp2lut_X_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5549|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5524" *) 3'b110;
  assign _3200_ = dp2lut_X_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5545|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5524" *) 3'b101;
  assign _3201_ = dp2lut_X_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5541|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5524" *) 3'b100;
  assign _3202_ = dp2lut_X_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5537|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5524" *) 2'b11;
  assign _3203_ = dp2lut_X_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5533|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5524" *) 2'b10;
  assign _3204_ = dp2lut_X_entry_2 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5529|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5524" *) 1'b1;
  assign _3205_ = ! (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5525|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5524" *) dp2lut_X_entry_2;
  assign _3206_ = dp2lut_Xinfo_2[17] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5520" *) raw_reg64 : _3140_;
  assign _3207_ = dp2lut_Xinfo_2[16] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5517" *) raw_reg0 : _3206_;
  assign _0266_ = _0394_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5516" *) _3207_ : lut_X_data_21;
  function [15:0] _7078_;
    input [15:0] a;
    input [1023:0] b;
    input [63:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5781|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5524" *)
    (* parallel_case *)
    casez (s)
      64'b???????????????????????????????????????????????????????????????1:
        _7078_ = b[15:0];
      64'b??????????????????????????????????????????????????????????????1?:
        _7078_ = b[31:16];
      64'b?????????????????????????????????????????????????????????????1??:
        _7078_ = b[47:32];
      64'b????????????????????????????????????????????????????????????1???:
        _7078_ = b[63:48];
      64'b???????????????????????????????????????????????????????????1????:
        _7078_ = b[79:64];
      64'b??????????????????????????????????????????????????????????1?????:
        _7078_ = b[95:80];
      64'b?????????????????????????????????????????????????????????1??????:
        _7078_ = b[111:96];
      64'b????????????????????????????????????????????????????????1???????:
        _7078_ = b[127:112];
      64'b???????????????????????????????????????????????????????1????????:
        _7078_ = b[143:128];
      64'b??????????????????????????????????????????????????????1?????????:
        _7078_ = b[159:144];
      64'b?????????????????????????????????????????????????????1??????????:
        _7078_ = b[175:160];
      64'b????????????????????????????????????????????????????1???????????:
        _7078_ = b[191:176];
      64'b???????????????????????????????????????????????????1????????????:
        _7078_ = b[207:192];
      64'b??????????????????????????????????????????????????1?????????????:
        _7078_ = b[223:208];
      64'b?????????????????????????????????????????????????1??????????????:
        _7078_ = b[239:224];
      64'b????????????????????????????????????????????????1???????????????:
        _7078_ = b[255:240];
      64'b???????????????????????????????????????????????1????????????????:
        _7078_ = b[271:256];
      64'b??????????????????????????????????????????????1?????????????????:
        _7078_ = b[287:272];
      64'b?????????????????????????????????????????????1??????????????????:
        _7078_ = b[303:288];
      64'b????????????????????????????????????????????1???????????????????:
        _7078_ = b[319:304];
      64'b???????????????????????????????????????????1????????????????????:
        _7078_ = b[335:320];
      64'b??????????????????????????????????????????1?????????????????????:
        _7078_ = b[351:336];
      64'b?????????????????????????????????????????1??????????????????????:
        _7078_ = b[367:352];
      64'b????????????????????????????????????????1???????????????????????:
        _7078_ = b[383:368];
      64'b???????????????????????????????????????1????????????????????????:
        _7078_ = b[399:384];
      64'b??????????????????????????????????????1?????????????????????????:
        _7078_ = b[415:400];
      64'b?????????????????????????????????????1??????????????????????????:
        _7078_ = b[431:416];
      64'b????????????????????????????????????1???????????????????????????:
        _7078_ = b[447:432];
      64'b???????????????????????????????????1????????????????????????????:
        _7078_ = b[463:448];
      64'b??????????????????????????????????1?????????????????????????????:
        _7078_ = b[479:464];
      64'b?????????????????????????????????1??????????????????????????????:
        _7078_ = b[495:480];
      64'b????????????????????????????????1???????????????????????????????:
        _7078_ = b[511:496];
      64'b???????????????????????????????1????????????????????????????????:
        _7078_ = b[527:512];
      64'b??????????????????????????????1?????????????????????????????????:
        _7078_ = b[543:528];
      64'b?????????????????????????????1??????????????????????????????????:
        _7078_ = b[559:544];
      64'b????????????????????????????1???????????????????????????????????:
        _7078_ = b[575:560];
      64'b???????????????????????????1????????????????????????????????????:
        _7078_ = b[591:576];
      64'b??????????????????????????1?????????????????????????????????????:
        _7078_ = b[607:592];
      64'b?????????????????????????1??????????????????????????????????????:
        _7078_ = b[623:608];
      64'b????????????????????????1???????????????????????????????????????:
        _7078_ = b[639:624];
      64'b???????????????????????1????????????????????????????????????????:
        _7078_ = b[655:640];
      64'b??????????????????????1?????????????????????????????????????????:
        _7078_ = b[671:656];
      64'b?????????????????????1??????????????????????????????????????????:
        _7078_ = b[687:672];
      64'b????????????????????1???????????????????????????????????????????:
        _7078_ = b[703:688];
      64'b???????????????????1????????????????????????????????????????????:
        _7078_ = b[719:704];
      64'b??????????????????1?????????????????????????????????????????????:
        _7078_ = b[735:720];
      64'b?????????????????1??????????????????????????????????????????????:
        _7078_ = b[751:736];
      64'b????????????????1???????????????????????????????????????????????:
        _7078_ = b[767:752];
      64'b???????????????1????????????????????????????????????????????????:
        _7078_ = b[783:768];
      64'b??????????????1?????????????????????????????????????????????????:
        _7078_ = b[799:784];
      64'b?????????????1??????????????????????????????????????????????????:
        _7078_ = b[815:800];
      64'b????????????1???????????????????????????????????????????????????:
        _7078_ = b[831:816];
      64'b???????????1????????????????????????????????????????????????????:
        _7078_ = b[847:832];
      64'b??????????1?????????????????????????????????????????????????????:
        _7078_ = b[863:848];
      64'b?????????1??????????????????????????????????????????????????????:
        _7078_ = b[879:864];
      64'b????????1???????????????????????????????????????????????????????:
        _7078_ = b[895:880];
      64'b???????1????????????????????????????????????????????????????????:
        _7078_ = b[911:896];
      64'b??????1?????????????????????????????????????????????????????????:
        _7078_ = b[927:912];
      64'b?????1??????????????????????????????????????????????????????????:
        _7078_ = b[943:928];
      64'b????1???????????????????????????????????????????????????????????:
        _7078_ = b[959:944];
      64'b???1????????????????????????????????????????????????????????????:
        _7078_ = b[975:960];
      64'b??1?????????????????????????????????????????????????????????????:
        _7078_ = b[991:976];
      64'b?1??????????????????????????????????????????????????????????????:
        _7078_ = b[1007:992];
      64'b1???????????????????????????????????????????????????????????????:
        _7078_ = b[1023:1008];
      default:
        _7078_ = a;
    endcase
  endfunction
  assign _3208_ = _7078_(raw_reg0, { raw_reg1, raw_reg2, raw_reg3, raw_reg4, raw_reg5, raw_reg6, raw_reg7, raw_reg8, raw_reg9, raw_reg10, raw_reg11, raw_reg12, raw_reg13, raw_reg14, raw_reg15, raw_reg16, raw_reg17, raw_reg18, raw_reg19, raw_reg20, raw_reg21, raw_reg22, raw_reg23, raw_reg24, raw_reg25, raw_reg26, raw_reg27, raw_reg28, raw_reg29, raw_reg30, raw_reg31, raw_reg32, raw_reg33, raw_reg34, raw_reg35, raw_reg36, raw_reg37, raw_reg38, raw_reg39, raw_reg40, raw_reg41, raw_reg42, raw_reg43, raw_reg44, raw_reg45, raw_reg46, raw_reg47, raw_reg48, raw_reg49, raw_reg50, raw_reg51, raw_reg52, raw_reg53, raw_reg54, raw_reg55, raw_reg56, raw_reg57, raw_reg58, raw_reg59, raw_reg60, raw_reg61, raw_reg62, raw_reg63, raw_reg64 }, { _3204_, _3203_, _3202_, _3201_, _3200_, _3199_, _3198_, _3197_, _3196_, _3195_, _3194_, _3193_, _3192_, _3191_, _3190_, _3189_, _3188_, _3187_, _3186_, _3185_, _3184_, _3183_, _3182_, _3181_, _3180_, _3179_, _3178_, _3177_, _3176_, _3175_, _3174_, _3173_, _3172_, _3171_, _3170_, _3169_, _3168_, _3167_, _3166_, _3165_, _3164_, _3163_, _3162_, _3161_, _3160_, _3159_, _3158_, _3157_, _3156_, _3155_, _3154_, _3153_, _3152_, _3151_, _3150_, _3149_, _3148_, _3147_, _3146_, _3145_, _3144_, _3143_, _3142_, _3141_ });
  assign _3209_ = dp2lut_Xinfo_2[17] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5520" *) raw_reg64 : _3208_;
  assign _3210_ = dp2lut_Xinfo_2[16] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5517" *) raw_reg0 : _3209_;
  assign _0265_ = _0394_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5516" *) _3210_ : lut_X_data_20;
  function [15:0] _7082_;
    input [15:0] a;
    input [1023:0] b;
    input [63:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5498|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5241" *)
    (* parallel_case *)
    casez (s)
      64'b???????????????????????????????????????????????????????????????1:
        _7082_ = b[15:0];
      64'b??????????????????????????????????????????????????????????????1?:
        _7082_ = b[31:16];
      64'b?????????????????????????????????????????????????????????????1??:
        _7082_ = b[47:32];
      64'b????????????????????????????????????????????????????????????1???:
        _7082_ = b[63:48];
      64'b???????????????????????????????????????????????????????????1????:
        _7082_ = b[79:64];
      64'b??????????????????????????????????????????????????????????1?????:
        _7082_ = b[95:80];
      64'b?????????????????????????????????????????????????????????1??????:
        _7082_ = b[111:96];
      64'b????????????????????????????????????????????????????????1???????:
        _7082_ = b[127:112];
      64'b???????????????????????????????????????????????????????1????????:
        _7082_ = b[143:128];
      64'b??????????????????????????????????????????????????????1?????????:
        _7082_ = b[159:144];
      64'b?????????????????????????????????????????????????????1??????????:
        _7082_ = b[175:160];
      64'b????????????????????????????????????????????????????1???????????:
        _7082_ = b[191:176];
      64'b???????????????????????????????????????????????????1????????????:
        _7082_ = b[207:192];
      64'b??????????????????????????????????????????????????1?????????????:
        _7082_ = b[223:208];
      64'b?????????????????????????????????????????????????1??????????????:
        _7082_ = b[239:224];
      64'b????????????????????????????????????????????????1???????????????:
        _7082_ = b[255:240];
      64'b???????????????????????????????????????????????1????????????????:
        _7082_ = b[271:256];
      64'b??????????????????????????????????????????????1?????????????????:
        _7082_ = b[287:272];
      64'b?????????????????????????????????????????????1??????????????????:
        _7082_ = b[303:288];
      64'b????????????????????????????????????????????1???????????????????:
        _7082_ = b[319:304];
      64'b???????????????????????????????????????????1????????????????????:
        _7082_ = b[335:320];
      64'b??????????????????????????????????????????1?????????????????????:
        _7082_ = b[351:336];
      64'b?????????????????????????????????????????1??????????????????????:
        _7082_ = b[367:352];
      64'b????????????????????????????????????????1???????????????????????:
        _7082_ = b[383:368];
      64'b???????????????????????????????????????1????????????????????????:
        _7082_ = b[399:384];
      64'b??????????????????????????????????????1?????????????????????????:
        _7082_ = b[415:400];
      64'b?????????????????????????????????????1??????????????????????????:
        _7082_ = b[431:416];
      64'b????????????????????????????????????1???????????????????????????:
        _7082_ = b[447:432];
      64'b???????????????????????????????????1????????????????????????????:
        _7082_ = b[463:448];
      64'b??????????????????????????????????1?????????????????????????????:
        _7082_ = b[479:464];
      64'b?????????????????????????????????1??????????????????????????????:
        _7082_ = b[495:480];
      64'b????????????????????????????????1???????????????????????????????:
        _7082_ = b[511:496];
      64'b???????????????????????????????1????????????????????????????????:
        _7082_ = b[527:512];
      64'b??????????????????????????????1?????????????????????????????????:
        _7082_ = b[543:528];
      64'b?????????????????????????????1??????????????????????????????????:
        _7082_ = b[559:544];
      64'b????????????????????????????1???????????????????????????????????:
        _7082_ = b[575:560];
      64'b???????????????????????????1????????????????????????????????????:
        _7082_ = b[591:576];
      64'b??????????????????????????1?????????????????????????????????????:
        _7082_ = b[607:592];
      64'b?????????????????????????1??????????????????????????????????????:
        _7082_ = b[623:608];
      64'b????????????????????????1???????????????????????????????????????:
        _7082_ = b[639:624];
      64'b???????????????????????1????????????????????????????????????????:
        _7082_ = b[655:640];
      64'b??????????????????????1?????????????????????????????????????????:
        _7082_ = b[671:656];
      64'b?????????????????????1??????????????????????????????????????????:
        _7082_ = b[687:672];
      64'b????????????????????1???????????????????????????????????????????:
        _7082_ = b[703:688];
      64'b???????????????????1????????????????????????????????????????????:
        _7082_ = b[719:704];
      64'b??????????????????1?????????????????????????????????????????????:
        _7082_ = b[735:720];
      64'b?????????????????1??????????????????????????????????????????????:
        _7082_ = b[751:736];
      64'b????????????????1???????????????????????????????????????????????:
        _7082_ = b[767:752];
      64'b???????????????1????????????????????????????????????????????????:
        _7082_ = b[783:768];
      64'b??????????????1?????????????????????????????????????????????????:
        _7082_ = b[799:784];
      64'b?????????????1??????????????????????????????????????????????????:
        _7082_ = b[815:800];
      64'b????????????1???????????????????????????????????????????????????:
        _7082_ = b[831:816];
      64'b???????????1????????????????????????????????????????????????????:
        _7082_ = b[847:832];
      64'b??????????1?????????????????????????????????????????????????????:
        _7082_ = b[863:848];
      64'b?????????1??????????????????????????????????????????????????????:
        _7082_ = b[879:864];
      64'b????????1???????????????????????????????????????????????????????:
        _7082_ = b[895:880];
      64'b???????1????????????????????????????????????????????????????????:
        _7082_ = b[911:896];
      64'b??????1?????????????????????????????????????????????????????????:
        _7082_ = b[927:912];
      64'b?????1??????????????????????????????????????????????????????????:
        _7082_ = b[943:928];
      64'b????1???????????????????????????????????????????????????????????:
        _7082_ = b[959:944];
      64'b???1????????????????????????????????????????????????????????????:
        _7082_ = b[975:960];
      64'b??1?????????????????????????????????????????????????????????????:
        _7082_ = b[991:976];
      64'b?1??????????????????????????????????????????????????????????????:
        _7082_ = b[1007:992];
      64'b1???????????????????????????????????????????????????????????????:
        _7082_ = b[1023:1008];
      default:
        _7082_ = a;
    endcase
  endfunction
  assign _3211_ = _7082_(raw_reg0, { raw_reg1, raw_reg2, raw_reg3, raw_reg4, raw_reg5, raw_reg6, raw_reg7, raw_reg8, raw_reg9, raw_reg10, raw_reg11, raw_reg12, raw_reg13, raw_reg14, raw_reg15, raw_reg16, raw_reg17, raw_reg18, raw_reg19, raw_reg20, raw_reg21, raw_reg22, raw_reg23, raw_reg24, raw_reg25, raw_reg26, raw_reg27, raw_reg28, raw_reg29, raw_reg30, raw_reg31, raw_reg32, raw_reg33, raw_reg34, raw_reg35, raw_reg36, raw_reg37, raw_reg38, raw_reg39, raw_reg40, raw_reg41, raw_reg42, raw_reg43, raw_reg44, raw_reg45, raw_reg46, raw_reg47, raw_reg48, raw_reg49, raw_reg50, raw_reg51, raw_reg52, raw_reg53, raw_reg54, raw_reg55, raw_reg56, raw_reg57, raw_reg58, raw_reg59, raw_reg60, raw_reg61, raw_reg62, raw_reg63, raw_reg64 }, { _3276_, _3275_, _3274_, _3273_, _3272_, _3271_, _3270_, _3269_, _3268_, _3267_, _3266_, _3265_, _3264_, _3263_, _3262_, _3261_, _3260_, _3259_, _3258_, _3257_, _3256_, _3255_, _3254_, _3253_, _3252_, _3251_, _3250_, _3249_, _3248_, _3247_, _3246_, _3245_, _3244_, _3243_, _3242_, _3241_, _3240_, _3239_, _3238_, _3237_, _3236_, _3235_, _3234_, _3233_, _3232_, _3231_, _3230_, _3229_, _3228_, _3227_, _3226_, _3225_, _3224_, _3223_, _3222_, _3221_, _3220_, _3219_, _3218_, _3217_, _3216_, _3215_, _3214_, _0416_ });
  assign _3212_ = dp2lut_X_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5498|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5241" *) 7'b1000000;
  assign _3213_ = dp2lut_X_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5494|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5241" *) 6'b111111;
  assign _3214_ = dp2lut_X_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5490|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5241" *) 6'b111110;
  assign _3215_ = dp2lut_X_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5486|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5241" *) 6'b111101;
  assign _3216_ = dp2lut_X_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5482|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5241" *) 6'b111100;
  assign _3217_ = dp2lut_X_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5478|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5241" *) 6'b111011;
  assign _3218_ = dp2lut_X_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5474|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5241" *) 6'b111010;
  assign _3219_ = dp2lut_X_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5470|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5241" *) 6'b111001;
  assign _3220_ = dp2lut_X_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5466|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5241" *) 6'b111000;
  assign _3221_ = dp2lut_X_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5462|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5241" *) 6'b110111;
  assign _3222_ = dp2lut_X_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5458|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5241" *) 6'b110110;
  assign _3223_ = dp2lut_X_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5454|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5241" *) 6'b110101;
  assign _3224_ = dp2lut_X_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5450|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5241" *) 6'b110100;
  assign _3225_ = dp2lut_X_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5446|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5241" *) 6'b110011;
  assign _3226_ = dp2lut_X_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5442|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5241" *) 6'b110010;
  assign _3227_ = dp2lut_X_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5438|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5241" *) 6'b110001;
  assign _3228_ = dp2lut_X_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5434|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5241" *) 6'b110000;
  assign _3229_ = dp2lut_X_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5430|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5241" *) 6'b101111;
  assign _3230_ = dp2lut_X_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5426|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5241" *) 6'b101110;
  assign _3231_ = dp2lut_X_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5422|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5241" *) 6'b101101;
  assign _3232_ = dp2lut_X_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5418|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5241" *) 6'b101100;
  assign _3233_ = dp2lut_X_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5414|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5241" *) 6'b101011;
  assign _3234_ = dp2lut_X_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5410|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5241" *) 6'b101010;
  assign _3235_ = dp2lut_X_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5406|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5241" *) 6'b101001;
  assign _3236_ = dp2lut_X_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5402|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5241" *) 6'b101000;
  assign _3237_ = dp2lut_X_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5398|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5241" *) 6'b100111;
  assign _3238_ = dp2lut_X_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5394|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5241" *) 6'b100110;
  assign _3239_ = dp2lut_X_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5390|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5241" *) 6'b100101;
  assign _3240_ = dp2lut_X_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5386|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5241" *) 6'b100100;
  assign _3241_ = dp2lut_X_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5382|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5241" *) 6'b100011;
  assign _3242_ = dp2lut_X_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5378|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5241" *) 6'b100010;
  assign _3243_ = dp2lut_X_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5374|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5241" *) 6'b100001;
  assign _3244_ = dp2lut_X_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5370|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5241" *) 6'b100000;
  assign _3245_ = dp2lut_X_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5366|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5241" *) 5'b11111;
  assign _3246_ = dp2lut_X_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5362|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5241" *) 5'b11110;
  assign _3247_ = dp2lut_X_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5358|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5241" *) 5'b11101;
  assign _3248_ = dp2lut_X_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5354|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5241" *) 5'b11100;
  assign _3249_ = dp2lut_X_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5350|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5241" *) 5'b11011;
  assign _3250_ = dp2lut_X_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5346|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5241" *) 5'b11010;
  assign _3251_ = dp2lut_X_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5342|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5241" *) 5'b11001;
  assign _3252_ = dp2lut_X_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5338|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5241" *) 5'b11000;
  assign _3253_ = dp2lut_X_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5334|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5241" *) 5'b10111;
  assign _3254_ = dp2lut_X_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5330|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5241" *) 5'b10110;
  assign _3255_ = dp2lut_X_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5326|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5241" *) 5'b10101;
  assign _3256_ = dp2lut_X_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5322|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5241" *) 5'b10100;
  assign _3257_ = dp2lut_X_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5318|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5241" *) 5'b10011;
  assign _3258_ = dp2lut_X_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5314|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5241" *) 5'b10010;
  assign _3259_ = dp2lut_X_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5310|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5241" *) 5'b10001;
  assign _3260_ = dp2lut_X_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5306|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5241" *) 5'b10000;
  assign _3261_ = dp2lut_X_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5302|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5241" *) 4'b1111;
  assign _3262_ = dp2lut_X_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5298|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5241" *) 4'b1110;
  assign _3263_ = dp2lut_X_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5294|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5241" *) 4'b1101;
  assign _3264_ = dp2lut_X_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5290|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5241" *) 4'b1100;
  assign _3265_ = dp2lut_X_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5286|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5241" *) 4'b1011;
  assign _3266_ = dp2lut_X_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5282|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5241" *) 4'b1010;
  assign _3267_ = dp2lut_X_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5278|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5241" *) 4'b1001;
  assign _3268_ = dp2lut_X_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5274|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5241" *) 4'b1000;
  assign _3269_ = dp2lut_X_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5270|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5241" *) 3'b111;
  assign _3270_ = dp2lut_X_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5266|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5241" *) 3'b110;
  assign _3271_ = dp2lut_X_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5262|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5241" *) 3'b101;
  assign _3272_ = dp2lut_X_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5258|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5241" *) 3'b100;
  assign _3273_ = dp2lut_X_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5254|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5241" *) 2'b11;
  assign _3274_ = dp2lut_X_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5250|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5241" *) 2'b10;
  assign _3275_ = dp2lut_X_entry_1 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5246|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5241" *) 1'b1;
  assign _3276_ = ! (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5242|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5241" *) dp2lut_X_entry_1;
  assign _3277_ = dp2lut_Xinfo_1[17] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5237" *) raw_reg64 : _3211_;
  assign _3278_ = dp2lut_Xinfo_1[16] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5234" *) raw_reg0 : _3277_;
  assign _0264_ = _0393_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5233" *) _3278_ : lut_X_data_11;
  function [15:0] _7151_;
    input [15:0] a;
    input [1023:0] b;
    input [63:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5498|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5241" *)
    (* parallel_case *)
    casez (s)
      64'b???????????????????????????????????????????????????????????????1:
        _7151_ = b[15:0];
      64'b??????????????????????????????????????????????????????????????1?:
        _7151_ = b[31:16];
      64'b?????????????????????????????????????????????????????????????1??:
        _7151_ = b[47:32];
      64'b????????????????????????????????????????????????????????????1???:
        _7151_ = b[63:48];
      64'b???????????????????????????????????????????????????????????1????:
        _7151_ = b[79:64];
      64'b??????????????????????????????????????????????????????????1?????:
        _7151_ = b[95:80];
      64'b?????????????????????????????????????????????????????????1??????:
        _7151_ = b[111:96];
      64'b????????????????????????????????????????????????????????1???????:
        _7151_ = b[127:112];
      64'b???????????????????????????????????????????????????????1????????:
        _7151_ = b[143:128];
      64'b??????????????????????????????????????????????????????1?????????:
        _7151_ = b[159:144];
      64'b?????????????????????????????????????????????????????1??????????:
        _7151_ = b[175:160];
      64'b????????????????????????????????????????????????????1???????????:
        _7151_ = b[191:176];
      64'b???????????????????????????????????????????????????1????????????:
        _7151_ = b[207:192];
      64'b??????????????????????????????????????????????????1?????????????:
        _7151_ = b[223:208];
      64'b?????????????????????????????????????????????????1??????????????:
        _7151_ = b[239:224];
      64'b????????????????????????????????????????????????1???????????????:
        _7151_ = b[255:240];
      64'b???????????????????????????????????????????????1????????????????:
        _7151_ = b[271:256];
      64'b??????????????????????????????????????????????1?????????????????:
        _7151_ = b[287:272];
      64'b?????????????????????????????????????????????1??????????????????:
        _7151_ = b[303:288];
      64'b????????????????????????????????????????????1???????????????????:
        _7151_ = b[319:304];
      64'b???????????????????????????????????????????1????????????????????:
        _7151_ = b[335:320];
      64'b??????????????????????????????????????????1?????????????????????:
        _7151_ = b[351:336];
      64'b?????????????????????????????????????????1??????????????????????:
        _7151_ = b[367:352];
      64'b????????????????????????????????????????1???????????????????????:
        _7151_ = b[383:368];
      64'b???????????????????????????????????????1????????????????????????:
        _7151_ = b[399:384];
      64'b??????????????????????????????????????1?????????????????????????:
        _7151_ = b[415:400];
      64'b?????????????????????????????????????1??????????????????????????:
        _7151_ = b[431:416];
      64'b????????????????????????????????????1???????????????????????????:
        _7151_ = b[447:432];
      64'b???????????????????????????????????1????????????????????????????:
        _7151_ = b[463:448];
      64'b??????????????????????????????????1?????????????????????????????:
        _7151_ = b[479:464];
      64'b?????????????????????????????????1??????????????????????????????:
        _7151_ = b[495:480];
      64'b????????????????????????????????1???????????????????????????????:
        _7151_ = b[511:496];
      64'b???????????????????????????????1????????????????????????????????:
        _7151_ = b[527:512];
      64'b??????????????????????????????1?????????????????????????????????:
        _7151_ = b[543:528];
      64'b?????????????????????????????1??????????????????????????????????:
        _7151_ = b[559:544];
      64'b????????????????????????????1???????????????????????????????????:
        _7151_ = b[575:560];
      64'b???????????????????????????1????????????????????????????????????:
        _7151_ = b[591:576];
      64'b??????????????????????????1?????????????????????????????????????:
        _7151_ = b[607:592];
      64'b?????????????????????????1??????????????????????????????????????:
        _7151_ = b[623:608];
      64'b????????????????????????1???????????????????????????????????????:
        _7151_ = b[639:624];
      64'b???????????????????????1????????????????????????????????????????:
        _7151_ = b[655:640];
      64'b??????????????????????1?????????????????????????????????????????:
        _7151_ = b[671:656];
      64'b?????????????????????1??????????????????????????????????????????:
        _7151_ = b[687:672];
      64'b????????????????????1???????????????????????????????????????????:
        _7151_ = b[703:688];
      64'b???????????????????1????????????????????????????????????????????:
        _7151_ = b[719:704];
      64'b??????????????????1?????????????????????????????????????????????:
        _7151_ = b[735:720];
      64'b?????????????????1??????????????????????????????????????????????:
        _7151_ = b[751:736];
      64'b????????????????1???????????????????????????????????????????????:
        _7151_ = b[767:752];
      64'b???????????????1????????????????????????????????????????????????:
        _7151_ = b[783:768];
      64'b??????????????1?????????????????????????????????????????????????:
        _7151_ = b[799:784];
      64'b?????????????1??????????????????????????????????????????????????:
        _7151_ = b[815:800];
      64'b????????????1???????????????????????????????????????????????????:
        _7151_ = b[831:816];
      64'b???????????1????????????????????????????????????????????????????:
        _7151_ = b[847:832];
      64'b??????????1?????????????????????????????????????????????????????:
        _7151_ = b[863:848];
      64'b?????????1??????????????????????????????????????????????????????:
        _7151_ = b[879:864];
      64'b????????1???????????????????????????????????????????????????????:
        _7151_ = b[895:880];
      64'b???????1????????????????????????????????????????????????????????:
        _7151_ = b[911:896];
      64'b??????1?????????????????????????????????????????????????????????:
        _7151_ = b[927:912];
      64'b?????1??????????????????????????????????????????????????????????:
        _7151_ = b[943:928];
      64'b????1???????????????????????????????????????????????????????????:
        _7151_ = b[959:944];
      64'b???1????????????????????????????????????????????????????????????:
        _7151_ = b[975:960];
      64'b??1?????????????????????????????????????????????????????????????:
        _7151_ = b[991:976];
      64'b?1??????????????????????????????????????????????????????????????:
        _7151_ = b[1007:992];
      64'b1???????????????????????????????????????????????????????????????:
        _7151_ = b[1023:1008];
      default:
        _7151_ = a;
    endcase
  endfunction
  assign _3279_ = _7151_(raw_reg0, { raw_reg1, raw_reg2, raw_reg3, raw_reg4, raw_reg5, raw_reg6, raw_reg7, raw_reg8, raw_reg9, raw_reg10, raw_reg11, raw_reg12, raw_reg13, raw_reg14, raw_reg15, raw_reg16, raw_reg17, raw_reg18, raw_reg19, raw_reg20, raw_reg21, raw_reg22, raw_reg23, raw_reg24, raw_reg25, raw_reg26, raw_reg27, raw_reg28, raw_reg29, raw_reg30, raw_reg31, raw_reg32, raw_reg33, raw_reg34, raw_reg35, raw_reg36, raw_reg37, raw_reg38, raw_reg39, raw_reg40, raw_reg41, raw_reg42, raw_reg43, raw_reg44, raw_reg45, raw_reg46, raw_reg47, raw_reg48, raw_reg49, raw_reg50, raw_reg51, raw_reg52, raw_reg53, raw_reg54, raw_reg55, raw_reg56, raw_reg57, raw_reg58, raw_reg59, raw_reg60, raw_reg61, raw_reg62, raw_reg63, raw_reg64 }, { _3275_, _3274_, _3273_, _3272_, _3271_, _3270_, _3269_, _3268_, _3267_, _3266_, _3265_, _3264_, _3263_, _3262_, _3261_, _3260_, _3259_, _3258_, _3257_, _3256_, _3255_, _3254_, _3253_, _3252_, _3251_, _3250_, _3249_, _3248_, _3247_, _3246_, _3245_, _3244_, _3243_, _3242_, _3241_, _3240_, _3239_, _3238_, _3237_, _3236_, _3235_, _3234_, _3233_, _3232_, _3231_, _3230_, _3229_, _3228_, _3227_, _3226_, _3225_, _3224_, _3223_, _3222_, _3221_, _3220_, _3219_, _3218_, _3217_, _3216_, _3215_, _3214_, _3213_, _3212_ });
  assign _3280_ = dp2lut_Xinfo_1[17] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5237" *) raw_reg64 : _3279_;
  assign _3281_ = dp2lut_Xinfo_1[16] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5234" *) raw_reg0 : _3280_;
  assign _0263_ = _0393_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5233" *) _3281_ : lut_X_data_10;
  function [15:0] _7155_;
    input [15:0] a;
    input [1023:0] b;
    input [63:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5215|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4958" *)
    (* parallel_case *)
    casez (s)
      64'b???????????????????????????????????????????????????????????????1:
        _7155_ = b[15:0];
      64'b??????????????????????????????????????????????????????????????1?:
        _7155_ = b[31:16];
      64'b?????????????????????????????????????????????????????????????1??:
        _7155_ = b[47:32];
      64'b????????????????????????????????????????????????????????????1???:
        _7155_ = b[63:48];
      64'b???????????????????????????????????????????????????????????1????:
        _7155_ = b[79:64];
      64'b??????????????????????????????????????????????????????????1?????:
        _7155_ = b[95:80];
      64'b?????????????????????????????????????????????????????????1??????:
        _7155_ = b[111:96];
      64'b????????????????????????????????????????????????????????1???????:
        _7155_ = b[127:112];
      64'b???????????????????????????????????????????????????????1????????:
        _7155_ = b[143:128];
      64'b??????????????????????????????????????????????????????1?????????:
        _7155_ = b[159:144];
      64'b?????????????????????????????????????????????????????1??????????:
        _7155_ = b[175:160];
      64'b????????????????????????????????????????????????????1???????????:
        _7155_ = b[191:176];
      64'b???????????????????????????????????????????????????1????????????:
        _7155_ = b[207:192];
      64'b??????????????????????????????????????????????????1?????????????:
        _7155_ = b[223:208];
      64'b?????????????????????????????????????????????????1??????????????:
        _7155_ = b[239:224];
      64'b????????????????????????????????????????????????1???????????????:
        _7155_ = b[255:240];
      64'b???????????????????????????????????????????????1????????????????:
        _7155_ = b[271:256];
      64'b??????????????????????????????????????????????1?????????????????:
        _7155_ = b[287:272];
      64'b?????????????????????????????????????????????1??????????????????:
        _7155_ = b[303:288];
      64'b????????????????????????????????????????????1???????????????????:
        _7155_ = b[319:304];
      64'b???????????????????????????????????????????1????????????????????:
        _7155_ = b[335:320];
      64'b??????????????????????????????????????????1?????????????????????:
        _7155_ = b[351:336];
      64'b?????????????????????????????????????????1??????????????????????:
        _7155_ = b[367:352];
      64'b????????????????????????????????????????1???????????????????????:
        _7155_ = b[383:368];
      64'b???????????????????????????????????????1????????????????????????:
        _7155_ = b[399:384];
      64'b??????????????????????????????????????1?????????????????????????:
        _7155_ = b[415:400];
      64'b?????????????????????????????????????1??????????????????????????:
        _7155_ = b[431:416];
      64'b????????????????????????????????????1???????????????????????????:
        _7155_ = b[447:432];
      64'b???????????????????????????????????1????????????????????????????:
        _7155_ = b[463:448];
      64'b??????????????????????????????????1?????????????????????????????:
        _7155_ = b[479:464];
      64'b?????????????????????????????????1??????????????????????????????:
        _7155_ = b[495:480];
      64'b????????????????????????????????1???????????????????????????????:
        _7155_ = b[511:496];
      64'b???????????????????????????????1????????????????????????????????:
        _7155_ = b[527:512];
      64'b??????????????????????????????1?????????????????????????????????:
        _7155_ = b[543:528];
      64'b?????????????????????????????1??????????????????????????????????:
        _7155_ = b[559:544];
      64'b????????????????????????????1???????????????????????????????????:
        _7155_ = b[575:560];
      64'b???????????????????????????1????????????????????????????????????:
        _7155_ = b[591:576];
      64'b??????????????????????????1?????????????????????????????????????:
        _7155_ = b[607:592];
      64'b?????????????????????????1??????????????????????????????????????:
        _7155_ = b[623:608];
      64'b????????????????????????1???????????????????????????????????????:
        _7155_ = b[639:624];
      64'b???????????????????????1????????????????????????????????????????:
        _7155_ = b[655:640];
      64'b??????????????????????1?????????????????????????????????????????:
        _7155_ = b[671:656];
      64'b?????????????????????1??????????????????????????????????????????:
        _7155_ = b[687:672];
      64'b????????????????????1???????????????????????????????????????????:
        _7155_ = b[703:688];
      64'b???????????????????1????????????????????????????????????????????:
        _7155_ = b[719:704];
      64'b??????????????????1?????????????????????????????????????????????:
        _7155_ = b[735:720];
      64'b?????????????????1??????????????????????????????????????????????:
        _7155_ = b[751:736];
      64'b????????????????1???????????????????????????????????????????????:
        _7155_ = b[767:752];
      64'b???????????????1????????????????????????????????????????????????:
        _7155_ = b[783:768];
      64'b??????????????1?????????????????????????????????????????????????:
        _7155_ = b[799:784];
      64'b?????????????1??????????????????????????????????????????????????:
        _7155_ = b[815:800];
      64'b????????????1???????????????????????????????????????????????????:
        _7155_ = b[831:816];
      64'b???????????1????????????????????????????????????????????????????:
        _7155_ = b[847:832];
      64'b??????????1?????????????????????????????????????????????????????:
        _7155_ = b[863:848];
      64'b?????????1??????????????????????????????????????????????????????:
        _7155_ = b[879:864];
      64'b????????1???????????????????????????????????????????????????????:
        _7155_ = b[895:880];
      64'b???????1????????????????????????????????????????????????????????:
        _7155_ = b[911:896];
      64'b??????1?????????????????????????????????????????????????????????:
        _7155_ = b[927:912];
      64'b?????1??????????????????????????????????????????????????????????:
        _7155_ = b[943:928];
      64'b????1???????????????????????????????????????????????????????????:
        _7155_ = b[959:944];
      64'b???1????????????????????????????????????????????????????????????:
        _7155_ = b[975:960];
      64'b??1?????????????????????????????????????????????????????????????:
        _7155_ = b[991:976];
      64'b?1??????????????????????????????????????????????????????????????:
        _7155_ = b[1007:992];
      64'b1???????????????????????????????????????????????????????????????:
        _7155_ = b[1023:1008];
      default:
        _7155_ = a;
    endcase
  endfunction
  assign _3282_ = _7155_(raw_reg0, { raw_reg1, raw_reg2, raw_reg3, raw_reg4, raw_reg5, raw_reg6, raw_reg7, raw_reg8, raw_reg9, raw_reg10, raw_reg11, raw_reg12, raw_reg13, raw_reg14, raw_reg15, raw_reg16, raw_reg17, raw_reg18, raw_reg19, raw_reg20, raw_reg21, raw_reg22, raw_reg23, raw_reg24, raw_reg25, raw_reg26, raw_reg27, raw_reg28, raw_reg29, raw_reg30, raw_reg31, raw_reg32, raw_reg33, raw_reg34, raw_reg35, raw_reg36, raw_reg37, raw_reg38, raw_reg39, raw_reg40, raw_reg41, raw_reg42, raw_reg43, raw_reg44, raw_reg45, raw_reg46, raw_reg47, raw_reg48, raw_reg49, raw_reg50, raw_reg51, raw_reg52, raw_reg53, raw_reg54, raw_reg55, raw_reg56, raw_reg57, raw_reg58, raw_reg59, raw_reg60, raw_reg61, raw_reg62, raw_reg63, raw_reg64 }, { _3347_, _3346_, _3345_, _3344_, _3343_, _3342_, _3341_, _3340_, _3339_, _3338_, _3337_, _3336_, _3335_, _3334_, _3333_, _3332_, _3331_, _3330_, _3329_, _3328_, _3327_, _3326_, _3325_, _3324_, _3323_, _3322_, _3321_, _3320_, _3319_, _3318_, _3317_, _3316_, _3315_, _3314_, _3313_, _3312_, _3311_, _3310_, _3309_, _3308_, _3307_, _3306_, _3305_, _3304_, _3303_, _3302_, _3301_, _3300_, _3299_, _3298_, _3297_, _3296_, _3295_, _3294_, _3293_, _3292_, _3291_, _3290_, _3289_, _3288_, _3287_, _3286_, _3285_, _0417_ });
  assign _3283_ = dp2lut_X_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5215|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4958" *) 7'b1000000;
  assign _3284_ = dp2lut_X_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5211|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4958" *) 6'b111111;
  assign _3285_ = dp2lut_X_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5207|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4958" *) 6'b111110;
  assign _3286_ = dp2lut_X_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5203|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4958" *) 6'b111101;
  assign _3287_ = dp2lut_X_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5199|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4958" *) 6'b111100;
  assign _3288_ = dp2lut_X_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5195|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4958" *) 6'b111011;
  assign _3289_ = dp2lut_X_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5191|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4958" *) 6'b111010;
  assign _3290_ = dp2lut_X_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5187|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4958" *) 6'b111001;
  assign _3291_ = dp2lut_X_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5183|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4958" *) 6'b111000;
  assign _3292_ = dp2lut_X_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5179|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4958" *) 6'b110111;
  assign _3293_ = dp2lut_X_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5175|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4958" *) 6'b110110;
  assign _3294_ = dp2lut_X_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5171|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4958" *) 6'b110101;
  assign _3295_ = dp2lut_X_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5167|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4958" *) 6'b110100;
  assign _3296_ = dp2lut_X_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5163|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4958" *) 6'b110011;
  assign _3297_ = dp2lut_X_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5159|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4958" *) 6'b110010;
  assign _3298_ = dp2lut_X_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5155|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4958" *) 6'b110001;
  assign _3299_ = dp2lut_X_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5151|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4958" *) 6'b110000;
  assign _3300_ = dp2lut_X_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5147|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4958" *) 6'b101111;
  assign _3301_ = dp2lut_X_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5143|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4958" *) 6'b101110;
  assign _3302_ = dp2lut_X_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5139|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4958" *) 6'b101101;
  assign _3303_ = dp2lut_X_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5135|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4958" *) 6'b101100;
  assign _3304_ = dp2lut_X_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5131|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4958" *) 6'b101011;
  assign _3305_ = dp2lut_X_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5127|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4958" *) 6'b101010;
  assign _3306_ = dp2lut_X_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5123|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4958" *) 6'b101001;
  assign _3307_ = dp2lut_X_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5119|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4958" *) 6'b101000;
  assign _3308_ = dp2lut_X_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5115|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4958" *) 6'b100111;
  assign _3309_ = dp2lut_X_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5111|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4958" *) 6'b100110;
  assign _3310_ = dp2lut_X_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5107|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4958" *) 6'b100101;
  assign _3311_ = dp2lut_X_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5103|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4958" *) 6'b100100;
  assign _3312_ = dp2lut_X_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5099|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4958" *) 6'b100011;
  assign _3313_ = dp2lut_X_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5095|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4958" *) 6'b100010;
  assign _3314_ = dp2lut_X_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5091|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4958" *) 6'b100001;
  assign _3315_ = dp2lut_X_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5087|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4958" *) 6'b100000;
  assign _3316_ = dp2lut_X_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5083|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4958" *) 5'b11111;
  assign _3317_ = dp2lut_X_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5079|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4958" *) 5'b11110;
  assign _3318_ = dp2lut_X_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5075|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4958" *) 5'b11101;
  assign _3319_ = dp2lut_X_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5071|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4958" *) 5'b11100;
  assign _3320_ = dp2lut_X_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5067|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4958" *) 5'b11011;
  assign _3321_ = dp2lut_X_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5063|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4958" *) 5'b11010;
  assign _3322_ = dp2lut_X_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5059|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4958" *) 5'b11001;
  assign _3323_ = dp2lut_X_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5055|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4958" *) 5'b11000;
  assign _3324_ = dp2lut_X_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5051|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4958" *) 5'b10111;
  assign _3325_ = dp2lut_X_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5047|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4958" *) 5'b10110;
  assign _3326_ = dp2lut_X_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5043|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4958" *) 5'b10101;
  assign _3327_ = dp2lut_X_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5039|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4958" *) 5'b10100;
  assign _3328_ = dp2lut_X_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5035|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4958" *) 5'b10011;
  assign _3329_ = dp2lut_X_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5031|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4958" *) 5'b10010;
  assign _3330_ = dp2lut_X_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5027|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4958" *) 5'b10001;
  assign _3331_ = dp2lut_X_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5023|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4958" *) 5'b10000;
  assign _3332_ = dp2lut_X_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5019|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4958" *) 4'b1111;
  assign _3333_ = dp2lut_X_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5015|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4958" *) 4'b1110;
  assign _3334_ = dp2lut_X_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5011|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4958" *) 4'b1101;
  assign _3335_ = dp2lut_X_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5007|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4958" *) 4'b1100;
  assign _3336_ = dp2lut_X_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5003|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4958" *) 4'b1011;
  assign _3337_ = dp2lut_X_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4999|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4958" *) 4'b1010;
  assign _3338_ = dp2lut_X_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4995|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4958" *) 4'b1001;
  assign _3339_ = dp2lut_X_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4991|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4958" *) 4'b1000;
  assign _3340_ = dp2lut_X_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4987|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4958" *) 3'b111;
  assign _3341_ = dp2lut_X_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4983|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4958" *) 3'b110;
  assign _3342_ = dp2lut_X_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4979|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4958" *) 3'b101;
  assign _3343_ = dp2lut_X_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4975|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4958" *) 3'b100;
  assign _3344_ = dp2lut_X_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4971|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4958" *) 2'b11;
  assign _3345_ = dp2lut_X_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4967|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4958" *) 2'b10;
  assign _3346_ = dp2lut_X_entry_0 == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4963|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4958" *) 1'b1;
  assign _3347_ = ! (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4959|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4958" *) dp2lut_X_entry_0;
  assign _3348_ = dp2lut_Xinfo_0[17] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4954" *) raw_reg64 : _3282_;
  assign _3349_ = dp2lut_Xinfo_0[16] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4951" *) raw_reg0 : _3348_;
  assign _0262_ = _0392_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4950" *) _3349_ : lut_X_data_01;
  function [15:0] _7224_;
    input [15:0] a;
    input [1023:0] b;
    input [63:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:5215|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4958" *)
    (* parallel_case *)
    casez (s)
      64'b???????????????????????????????????????????????????????????????1:
        _7224_ = b[15:0];
      64'b??????????????????????????????????????????????????????????????1?:
        _7224_ = b[31:16];
      64'b?????????????????????????????????????????????????????????????1??:
        _7224_ = b[47:32];
      64'b????????????????????????????????????????????????????????????1???:
        _7224_ = b[63:48];
      64'b???????????????????????????????????????????????????????????1????:
        _7224_ = b[79:64];
      64'b??????????????????????????????????????????????????????????1?????:
        _7224_ = b[95:80];
      64'b?????????????????????????????????????????????????????????1??????:
        _7224_ = b[111:96];
      64'b????????????????????????????????????????????????????????1???????:
        _7224_ = b[127:112];
      64'b???????????????????????????????????????????????????????1????????:
        _7224_ = b[143:128];
      64'b??????????????????????????????????????????????????????1?????????:
        _7224_ = b[159:144];
      64'b?????????????????????????????????????????????????????1??????????:
        _7224_ = b[175:160];
      64'b????????????????????????????????????????????????????1???????????:
        _7224_ = b[191:176];
      64'b???????????????????????????????????????????????????1????????????:
        _7224_ = b[207:192];
      64'b??????????????????????????????????????????????????1?????????????:
        _7224_ = b[223:208];
      64'b?????????????????????????????????????????????????1??????????????:
        _7224_ = b[239:224];
      64'b????????????????????????????????????????????????1???????????????:
        _7224_ = b[255:240];
      64'b???????????????????????????????????????????????1????????????????:
        _7224_ = b[271:256];
      64'b??????????????????????????????????????????????1?????????????????:
        _7224_ = b[287:272];
      64'b?????????????????????????????????????????????1??????????????????:
        _7224_ = b[303:288];
      64'b????????????????????????????????????????????1???????????????????:
        _7224_ = b[319:304];
      64'b???????????????????????????????????????????1????????????????????:
        _7224_ = b[335:320];
      64'b??????????????????????????????????????????1?????????????????????:
        _7224_ = b[351:336];
      64'b?????????????????????????????????????????1??????????????????????:
        _7224_ = b[367:352];
      64'b????????????????????????????????????????1???????????????????????:
        _7224_ = b[383:368];
      64'b???????????????????????????????????????1????????????????????????:
        _7224_ = b[399:384];
      64'b??????????????????????????????????????1?????????????????????????:
        _7224_ = b[415:400];
      64'b?????????????????????????????????????1??????????????????????????:
        _7224_ = b[431:416];
      64'b????????????????????????????????????1???????????????????????????:
        _7224_ = b[447:432];
      64'b???????????????????????????????????1????????????????????????????:
        _7224_ = b[463:448];
      64'b??????????????????????????????????1?????????????????????????????:
        _7224_ = b[479:464];
      64'b?????????????????????????????????1??????????????????????????????:
        _7224_ = b[495:480];
      64'b????????????????????????????????1???????????????????????????????:
        _7224_ = b[511:496];
      64'b???????????????????????????????1????????????????????????????????:
        _7224_ = b[527:512];
      64'b??????????????????????????????1?????????????????????????????????:
        _7224_ = b[543:528];
      64'b?????????????????????????????1??????????????????????????????????:
        _7224_ = b[559:544];
      64'b????????????????????????????1???????????????????????????????????:
        _7224_ = b[575:560];
      64'b???????????????????????????1????????????????????????????????????:
        _7224_ = b[591:576];
      64'b??????????????????????????1?????????????????????????????????????:
        _7224_ = b[607:592];
      64'b?????????????????????????1??????????????????????????????????????:
        _7224_ = b[623:608];
      64'b????????????????????????1???????????????????????????????????????:
        _7224_ = b[639:624];
      64'b???????????????????????1????????????????????????????????????????:
        _7224_ = b[655:640];
      64'b??????????????????????1?????????????????????????????????????????:
        _7224_ = b[671:656];
      64'b?????????????????????1??????????????????????????????????????????:
        _7224_ = b[687:672];
      64'b????????????????????1???????????????????????????????????????????:
        _7224_ = b[703:688];
      64'b???????????????????1????????????????????????????????????????????:
        _7224_ = b[719:704];
      64'b??????????????????1?????????????????????????????????????????????:
        _7224_ = b[735:720];
      64'b?????????????????1??????????????????????????????????????????????:
        _7224_ = b[751:736];
      64'b????????????????1???????????????????????????????????????????????:
        _7224_ = b[767:752];
      64'b???????????????1????????????????????????????????????????????????:
        _7224_ = b[783:768];
      64'b??????????????1?????????????????????????????????????????????????:
        _7224_ = b[799:784];
      64'b?????????????1??????????????????????????????????????????????????:
        _7224_ = b[815:800];
      64'b????????????1???????????????????????????????????????????????????:
        _7224_ = b[831:816];
      64'b???????????1????????????????????????????????????????????????????:
        _7224_ = b[847:832];
      64'b??????????1?????????????????????????????????????????????????????:
        _7224_ = b[863:848];
      64'b?????????1??????????????????????????????????????????????????????:
        _7224_ = b[879:864];
      64'b????????1???????????????????????????????????????????????????????:
        _7224_ = b[895:880];
      64'b???????1????????????????????????????????????????????????????????:
        _7224_ = b[911:896];
      64'b??????1?????????????????????????????????????????????????????????:
        _7224_ = b[927:912];
      64'b?????1??????????????????????????????????????????????????????????:
        _7224_ = b[943:928];
      64'b????1???????????????????????????????????????????????????????????:
        _7224_ = b[959:944];
      64'b???1????????????????????????????????????????????????????????????:
        _7224_ = b[975:960];
      64'b??1?????????????????????????????????????????????????????????????:
        _7224_ = b[991:976];
      64'b?1??????????????????????????????????????????????????????????????:
        _7224_ = b[1007:992];
      64'b1???????????????????????????????????????????????????????????????:
        _7224_ = b[1023:1008];
      default:
        _7224_ = a;
    endcase
  endfunction
  assign _3350_ = _7224_(raw_reg0, { raw_reg1, raw_reg2, raw_reg3, raw_reg4, raw_reg5, raw_reg6, raw_reg7, raw_reg8, raw_reg9, raw_reg10, raw_reg11, raw_reg12, raw_reg13, raw_reg14, raw_reg15, raw_reg16, raw_reg17, raw_reg18, raw_reg19, raw_reg20, raw_reg21, raw_reg22, raw_reg23, raw_reg24, raw_reg25, raw_reg26, raw_reg27, raw_reg28, raw_reg29, raw_reg30, raw_reg31, raw_reg32, raw_reg33, raw_reg34, raw_reg35, raw_reg36, raw_reg37, raw_reg38, raw_reg39, raw_reg40, raw_reg41, raw_reg42, raw_reg43, raw_reg44, raw_reg45, raw_reg46, raw_reg47, raw_reg48, raw_reg49, raw_reg50, raw_reg51, raw_reg52, raw_reg53, raw_reg54, raw_reg55, raw_reg56, raw_reg57, raw_reg58, raw_reg59, raw_reg60, raw_reg61, raw_reg62, raw_reg63, raw_reg64 }, { _3346_, _3345_, _3344_, _3343_, _3342_, _3341_, _3340_, _3339_, _3338_, _3337_, _3336_, _3335_, _3334_, _3333_, _3332_, _3331_, _3330_, _3329_, _3328_, _3327_, _3326_, _3325_, _3324_, _3323_, _3322_, _3321_, _3320_, _3319_, _3318_, _3317_, _3316_, _3315_, _3314_, _3313_, _3312_, _3311_, _3310_, _3309_, _3308_, _3307_, _3306_, _3305_, _3304_, _3303_, _3302_, _3301_, _3300_, _3299_, _3298_, _3297_, _3296_, _3295_, _3294_, _3293_, _3292_, _3291_, _3290_, _3289_, _3288_, _3287_, _3286_, _3285_, _3284_, _3283_ });
  assign _3351_ = dp2lut_Xinfo_0[17] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4954" *) raw_reg64 : _3350_;
  assign _3352_ = dp2lut_Xinfo_0[16] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4951" *) raw_reg0 : _3351_;
  assign _0261_ = _0392_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4950" *) _3352_ : lut_X_data_00;
  function [0:0] _7228_;
    input [0:0] a;
    input [3:0] b;
    input [3:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4848|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4843" *)
    (* parallel_case *)
    casez (s)
      4'b???1:
        _7228_ = b[0:0];
      4'b??1?:
        _7228_ = b[1:1];
      4'b?1??:
        _7228_ = b[2:2];
      4'b1???:
        _7228_ = b[3:3];
      default:
        _7228_ = a;
    endcase
  endfunction
  assign _0383_ = _7228_(1'b0, { reg2dp_lut_hybrid_priority, 1'b1, reg2dp_lut_uflow_priority, reg2dp_lut_oflow_priority }, { _3358_, _3356_, _3354_, _3353_ });
  assign _3353_ = { dp2lut_Xinfo_7[17:16], dp2lut_Yinfo_7[17:16] } == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4848|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4843" *) 4'b1010;
  assign _3354_ = { dp2lut_Xinfo_7[17:16], dp2lut_Yinfo_7[17:16] } == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4847|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4843" *) 3'b101;
  assign _3356_ = | (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4846|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4843" *) { _3355_[0], _3355_[1] };
  assign _3355_[0] = { dp2lut_Xinfo_7[17:16], dp2lut_Yinfo_7[17:16] } == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4846|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4843" *) 3'b100;
  assign _3355_[1] = { dp2lut_Xinfo_7[17:16], dp2lut_Yinfo_7[17:16] } == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4846|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4843" *) 4'b1000;
  assign _3358_ = | (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4844|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4843" *) { _3357_[0], _3357_[1], _3357_[2] };
  assign _3357_[0] = ! (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4844|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4843" *) { dp2lut_Xinfo_7[17:16], dp2lut_Yinfo_7[17:16] };
  assign _3357_[1] = { dp2lut_Xinfo_7[17:16], dp2lut_Yinfo_7[17:16] } == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4844|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4843" *) 3'b110;
  assign _3357_[2] = { dp2lut_Xinfo_7[17:16], dp2lut_Yinfo_7[17:16] } == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4844|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4843" *) 4'b1001;
  assign lut_Y_sel[7] = int8_en ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4842" *) _0383_ : 1'b0;
  function [0:0] _7239_;
    input [0:0] a;
    input [3:0] b;
    input [3:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4828|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4823" *)
    (* parallel_case *)
    casez (s)
      4'b???1:
        _7239_ = b[0:0];
      4'b??1?:
        _7239_ = b[1:1];
      4'b?1??:
        _7239_ = b[2:2];
      4'b1???:
        _7239_ = b[3:3];
      default:
        _7239_ = a;
    endcase
  endfunction
  assign _0382_ = _7239_(1'b0, { reg2dp_lut_hybrid_priority, 1'b1, reg2dp_lut_uflow_priority, reg2dp_lut_oflow_priority }, { _3364_, _3362_, _3360_, _3359_ });
  assign _3359_ = { dp2lut_Xinfo_6[17:16], dp2lut_Yinfo_6[17:16] } == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4828|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4823" *) 4'b1010;
  assign _3360_ = { dp2lut_Xinfo_6[17:16], dp2lut_Yinfo_6[17:16] } == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4827|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4823" *) 3'b101;
  assign _3362_ = | (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4826|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4823" *) { _3361_[0], _3361_[1] };
  assign _3361_[0] = { dp2lut_Xinfo_6[17:16], dp2lut_Yinfo_6[17:16] } == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4826|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4823" *) 3'b100;
  assign _3361_[1] = { dp2lut_Xinfo_6[17:16], dp2lut_Yinfo_6[17:16] } == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4826|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4823" *) 4'b1000;
  assign _3364_ = | (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4824|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4823" *) { _3363_[0], _3363_[1], _3363_[2] };
  assign _3363_[0] = ! (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4824|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4823" *) { dp2lut_Xinfo_6[17:16], dp2lut_Yinfo_6[17:16] };
  assign _3363_[1] = { dp2lut_Xinfo_6[17:16], dp2lut_Yinfo_6[17:16] } == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4824|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4823" *) 3'b110;
  assign _3363_[2] = { dp2lut_Xinfo_6[17:16], dp2lut_Yinfo_6[17:16] } == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4824|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4823" *) 4'b1001;
  assign lut_Y_sel[6] = int8_en ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4822" *) _0382_ : 1'b0;
  function [0:0] _7250_;
    input [0:0] a;
    input [3:0] b;
    input [3:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4808|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4803" *)
    (* parallel_case *)
    casez (s)
      4'b???1:
        _7250_ = b[0:0];
      4'b??1?:
        _7250_ = b[1:1];
      4'b?1??:
        _7250_ = b[2:2];
      4'b1???:
        _7250_ = b[3:3];
      default:
        _7250_ = a;
    endcase
  endfunction
  assign _0381_ = _7250_(1'b0, { reg2dp_lut_hybrid_priority, 1'b1, reg2dp_lut_uflow_priority, reg2dp_lut_oflow_priority }, { _3370_, _3368_, _3366_, _3365_ });
  assign _3365_ = { dp2lut_Xinfo_5[17:16], dp2lut_Yinfo_5[17:16] } == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4808|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4803" *) 4'b1010;
  assign _3366_ = { dp2lut_Xinfo_5[17:16], dp2lut_Yinfo_5[17:16] } == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4807|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4803" *) 3'b101;
  assign _3368_ = | (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4806|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4803" *) { _3367_[0], _3367_[1] };
  assign _3367_[0] = { dp2lut_Xinfo_5[17:16], dp2lut_Yinfo_5[17:16] } == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4806|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4803" *) 3'b100;
  assign _3367_[1] = { dp2lut_Xinfo_5[17:16], dp2lut_Yinfo_5[17:16] } == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4806|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4803" *) 4'b1000;
  assign _3370_ = | (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4804|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4803" *) { _3369_[0], _3369_[1], _3369_[2] };
  assign _3369_[0] = ! (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4804|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4803" *) { dp2lut_Xinfo_5[17:16], dp2lut_Yinfo_5[17:16] };
  assign _3369_[1] = { dp2lut_Xinfo_5[17:16], dp2lut_Yinfo_5[17:16] } == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4804|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4803" *) 3'b110;
  assign _3369_[2] = { dp2lut_Xinfo_5[17:16], dp2lut_Yinfo_5[17:16] } == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4804|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4803" *) 4'b1001;
  assign lut_Y_sel[5] = int8_en ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4802" *) _0381_ : 1'b0;
  function [0:0] _7261_;
    input [0:0] a;
    input [3:0] b;
    input [3:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4788|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4783" *)
    (* parallel_case *)
    casez (s)
      4'b???1:
        _7261_ = b[0:0];
      4'b??1?:
        _7261_ = b[1:1];
      4'b?1??:
        _7261_ = b[2:2];
      4'b1???:
        _7261_ = b[3:3];
      default:
        _7261_ = a;
    endcase
  endfunction
  assign _0380_ = _7261_(1'b0, { reg2dp_lut_hybrid_priority, 1'b1, reg2dp_lut_uflow_priority, reg2dp_lut_oflow_priority }, { _3376_, _3374_, _3372_, _3371_ });
  assign _3371_ = { dp2lut_Xinfo_4[17:16], dp2lut_Yinfo_4[17:16] } == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4788|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4783" *) 4'b1010;
  assign _3372_ = { dp2lut_Xinfo_4[17:16], dp2lut_Yinfo_4[17:16] } == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4787|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4783" *) 3'b101;
  assign _3374_ = | (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4786|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4783" *) { _3373_[0], _3373_[1] };
  assign _3373_[0] = { dp2lut_Xinfo_4[17:16], dp2lut_Yinfo_4[17:16] } == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4786|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4783" *) 3'b100;
  assign _3373_[1] = { dp2lut_Xinfo_4[17:16], dp2lut_Yinfo_4[17:16] } == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4786|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4783" *) 4'b1000;
  assign _3376_ = | (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4784|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4783" *) { _3375_[0], _3375_[1], _3375_[2] };
  assign _3375_[0] = ! (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4784|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4783" *) { dp2lut_Xinfo_4[17:16], dp2lut_Yinfo_4[17:16] };
  assign _3375_[1] = { dp2lut_Xinfo_4[17:16], dp2lut_Yinfo_4[17:16] } == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4784|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4783" *) 3'b110;
  assign _3375_[2] = { dp2lut_Xinfo_4[17:16], dp2lut_Yinfo_4[17:16] } == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4784|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4783" *) 4'b1001;
  assign lut_Y_sel[4] = int8_en ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4782" *) _0380_ : 1'b0;
  function [0:0] _7272_;
    input [0:0] a;
    input [3:0] b;
    input [3:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4770|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4765" *)
    (* parallel_case *)
    casez (s)
      4'b???1:
        _7272_ = b[0:0];
      4'b??1?:
        _7272_ = b[1:1];
      4'b?1??:
        _7272_ = b[2:2];
      4'b1???:
        _7272_ = b[3:3];
      default:
        _7272_ = a;
    endcase
  endfunction
  assign lut_Y_sel[3] = _7272_(1'b0, { reg2dp_lut_hybrid_priority, 1'b1, reg2dp_lut_uflow_priority, reg2dp_lut_oflow_priority }, { _3382_, _3380_, _3378_, _3377_ });
  assign _3377_ = { dp2lut_Xinfo_3[17:16], dp2lut_Yinfo_3[17:16] } == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4770|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4765" *) 4'b1010;
  assign _3378_ = { dp2lut_Xinfo_3[17:16], dp2lut_Yinfo_3[17:16] } == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4769|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4765" *) 3'b101;
  assign _3380_ = | (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4768|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4765" *) { _3379_[0], _3379_[1] };
  assign _3379_[0] = { dp2lut_Xinfo_3[17:16], dp2lut_Yinfo_3[17:16] } == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4768|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4765" *) 3'b100;
  assign _3379_[1] = { dp2lut_Xinfo_3[17:16], dp2lut_Yinfo_3[17:16] } == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4768|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4765" *) 4'b1000;
  assign _3382_ = | (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4766|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4765" *) { _3381_[0], _3381_[1], _3381_[2] };
  assign _3381_[0] = ! (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4766|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4765" *) { dp2lut_Xinfo_3[17:16], dp2lut_Yinfo_3[17:16] };
  assign _3381_[1] = { dp2lut_Xinfo_3[17:16], dp2lut_Yinfo_3[17:16] } == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4766|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4765" *) 3'b110;
  assign _3381_[2] = { dp2lut_Xinfo_3[17:16], dp2lut_Yinfo_3[17:16] } == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4766|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4765" *) 4'b1001;
  function [0:0] _7282_;
    input [0:0] a;
    input [3:0] b;
    input [3:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4754|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4749" *)
    (* parallel_case *)
    casez (s)
      4'b???1:
        _7282_ = b[0:0];
      4'b??1?:
        _7282_ = b[1:1];
      4'b?1??:
        _7282_ = b[2:2];
      4'b1???:
        _7282_ = b[3:3];
      default:
        _7282_ = a;
    endcase
  endfunction
  assign lut_Y_sel[2] = _7282_(1'b0, { reg2dp_lut_hybrid_priority, 1'b1, reg2dp_lut_uflow_priority, reg2dp_lut_oflow_priority }, { _3388_, _3386_, _3384_, _3383_ });
  assign _3383_ = { dp2lut_Xinfo_2[17:16], dp2lut_Yinfo_2[17:16] } == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4754|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4749" *) 4'b1010;
  assign _3384_ = { dp2lut_Xinfo_2[17:16], dp2lut_Yinfo_2[17:16] } == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4753|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4749" *) 3'b101;
  assign _3386_ = | (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4752|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4749" *) { _3385_[0], _3385_[1] };
  assign _3385_[0] = { dp2lut_Xinfo_2[17:16], dp2lut_Yinfo_2[17:16] } == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4752|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4749" *) 3'b100;
  assign _3385_[1] = { dp2lut_Xinfo_2[17:16], dp2lut_Yinfo_2[17:16] } == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4752|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4749" *) 4'b1000;
  assign _3388_ = | (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4750|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4749" *) { _3387_[0], _3387_[1], _3387_[2] };
  assign _3387_[0] = ! (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4750|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4749" *) { dp2lut_Xinfo_2[17:16], dp2lut_Yinfo_2[17:16] };
  assign _3387_[1] = { dp2lut_Xinfo_2[17:16], dp2lut_Yinfo_2[17:16] } == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4750|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4749" *) 3'b110;
  assign _3387_[2] = { dp2lut_Xinfo_2[17:16], dp2lut_Yinfo_2[17:16] } == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4750|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4749" *) 4'b1001;
  function [0:0] _7292_;
    input [0:0] a;
    input [3:0] b;
    input [3:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4738|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4733" *)
    (* parallel_case *)
    casez (s)
      4'b???1:
        _7292_ = b[0:0];
      4'b??1?:
        _7292_ = b[1:1];
      4'b?1??:
        _7292_ = b[2:2];
      4'b1???:
        _7292_ = b[3:3];
      default:
        _7292_ = a;
    endcase
  endfunction
  assign lut_Y_sel[1] = _7292_(1'b0, { reg2dp_lut_hybrid_priority, 1'b1, reg2dp_lut_uflow_priority, reg2dp_lut_oflow_priority }, { _3394_, _3392_, _3390_, _3389_ });
  assign _3389_ = { dp2lut_Xinfo_1[17:16], dp2lut_Yinfo_1[17:16] } == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4738|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4733" *) 4'b1010;
  assign _3390_ = { dp2lut_Xinfo_1[17:16], dp2lut_Yinfo_1[17:16] } == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4737|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4733" *) 3'b101;
  assign _3392_ = | (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4736|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4733" *) { _3391_[0], _3391_[1] };
  assign _3391_[0] = { dp2lut_Xinfo_1[17:16], dp2lut_Yinfo_1[17:16] } == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4736|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4733" *) 3'b100;
  assign _3391_[1] = { dp2lut_Xinfo_1[17:16], dp2lut_Yinfo_1[17:16] } == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4736|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4733" *) 4'b1000;
  assign _3394_ = | (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4734|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4733" *) { _3393_[0], _3393_[1], _3393_[2] };
  assign _3393_[0] = ! (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4734|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4733" *) { dp2lut_Xinfo_1[17:16], dp2lut_Yinfo_1[17:16] };
  assign _3393_[1] = { dp2lut_Xinfo_1[17:16], dp2lut_Yinfo_1[17:16] } == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4734|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4733" *) 3'b110;
  assign _3393_[2] = { dp2lut_Xinfo_1[17:16], dp2lut_Yinfo_1[17:16] } == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4734|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4733" *) 4'b1001;
  function [0:0] _7302_;
    input [0:0] a;
    input [3:0] b;
    input [3:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4722|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4717" *)
    (* parallel_case *)
    casez (s)
      4'b???1:
        _7302_ = b[0:0];
      4'b??1?:
        _7302_ = b[1:1];
      4'b?1??:
        _7302_ = b[2:2];
      4'b1???:
        _7302_ = b[3:3];
      default:
        _7302_ = a;
    endcase
  endfunction
  assign lut_Y_sel[0] = _7302_(1'b0, { reg2dp_lut_hybrid_priority, 1'b1, reg2dp_lut_uflow_priority, reg2dp_lut_oflow_priority }, { _3400_, _3398_, _3396_, _3395_ });
  assign _3395_ = { dp2lut_Xinfo_0[17:16], dp2lut_Yinfo_0[17:16] } == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4722|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4717" *) 4'b1010;
  assign _3396_ = { dp2lut_Xinfo_0[17:16], dp2lut_Yinfo_0[17:16] } == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4721|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4717" *) 3'b101;
  assign _3398_ = | (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4720|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4717" *) { _3397_[0], _3397_[1] };
  assign _3397_[0] = { dp2lut_Xinfo_0[17:16], dp2lut_Yinfo_0[17:16] } == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4720|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4717" *) 3'b100;
  assign _3397_[1] = { dp2lut_Xinfo_0[17:16], dp2lut_Yinfo_0[17:16] } == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4720|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4717" *) 4'b1000;
  assign _3400_ = | (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4718|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4717" *) { _3399_[0], _3399_[1], _3399_[2] };
  assign _3399_[0] = ! (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4718|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4717" *) { dp2lut_Xinfo_0[17:16], dp2lut_Yinfo_0[17:16] };
  assign _3399_[1] = { dp2lut_Xinfo_0[17:16], dp2lut_Yinfo_0[17:16] } == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4718|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4717" *) 3'b110;
  assign _3399_[2] = { dp2lut_Xinfo_0[17:16], dp2lut_Yinfo_0[17:16] } == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4718|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4717" *) 4'b1001;
  function [0:0] _7312_;
    input [0:0] a;
    input [3:0] b;
    input [3:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4704|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4699" *)
    (* parallel_case *)
    casez (s)
      4'b???1:
        _7312_ = b[0:0];
      4'b??1?:
        _7312_ = b[1:1];
      4'b?1??:
        _7312_ = b[2:2];
      4'b1???:
        _7312_ = b[3:3];
      default:
        _7312_ = a;
    endcase
  endfunction
  assign _0379_ = _7312_(1'b0, { _0677_, 1'b1, _0678_, _0679_ }, { _3358_, _3402_, _3354_, _3353_ });
  assign _3402_ = | (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4701|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4699" *) { _3401_[0], _3401_[1] };
  assign _3401_[0] = { dp2lut_Xinfo_7[17:16], dp2lut_Yinfo_7[17:16] } == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4701|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4699" *) 1'b1;
  assign _3401_[1] = { dp2lut_Xinfo_7[17:16], dp2lut_Yinfo_7[17:16] } == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4701|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4699" *) 2'b10;
  assign lut_X_sel[7] = int8_en ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4698" *) _0379_ : 1'b0;
  function [0:0] _7317_;
    input [0:0] a;
    input [3:0] b;
    input [3:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4684|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4679" *)
    (* parallel_case *)
    casez (s)
      4'b???1:
        _7317_ = b[0:0];
      4'b??1?:
        _7317_ = b[1:1];
      4'b?1??:
        _7317_ = b[2:2];
      4'b1???:
        _7317_ = b[3:3];
      default:
        _7317_ = a;
    endcase
  endfunction
  assign _0378_ = _7317_(1'b0, { _0677_, 1'b1, _0678_, _0679_ }, { _3364_, _3404_, _3360_, _3359_ });
  assign _3404_ = | (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4681|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4679" *) { _3403_[0], _3403_[1] };
  assign _3403_[0] = { dp2lut_Xinfo_6[17:16], dp2lut_Yinfo_6[17:16] } == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4681|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4679" *) 1'b1;
  assign _3403_[1] = { dp2lut_Xinfo_6[17:16], dp2lut_Yinfo_6[17:16] } == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4681|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4679" *) 2'b10;
  assign lut_X_sel[6] = int8_en ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4678" *) _0378_ : 1'b0;
  function [0:0] _7322_;
    input [0:0] a;
    input [3:0] b;
    input [3:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4664|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4659" *)
    (* parallel_case *)
    casez (s)
      4'b???1:
        _7322_ = b[0:0];
      4'b??1?:
        _7322_ = b[1:1];
      4'b?1??:
        _7322_ = b[2:2];
      4'b1???:
        _7322_ = b[3:3];
      default:
        _7322_ = a;
    endcase
  endfunction
  assign _0377_ = _7322_(1'b0, { _0677_, 1'b1, _0678_, _0679_ }, { _3370_, _3406_, _3366_, _3365_ });
  assign _3406_ = | (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4661|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4659" *) { _3405_[0], _3405_[1] };
  assign _3405_[0] = { dp2lut_Xinfo_5[17:16], dp2lut_Yinfo_5[17:16] } == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4661|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4659" *) 1'b1;
  assign _3405_[1] = { dp2lut_Xinfo_5[17:16], dp2lut_Yinfo_5[17:16] } == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4661|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4659" *) 2'b10;
  assign lut_X_sel[5] = int8_en ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4658" *) _0377_ : 1'b0;
  function [0:0] _7327_;
    input [0:0] a;
    input [3:0] b;
    input [3:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4644|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4639" *)
    (* parallel_case *)
    casez (s)
      4'b???1:
        _7327_ = b[0:0];
      4'b??1?:
        _7327_ = b[1:1];
      4'b?1??:
        _7327_ = b[2:2];
      4'b1???:
        _7327_ = b[3:3];
      default:
        _7327_ = a;
    endcase
  endfunction
  assign _0376_ = _7327_(1'b0, { _0677_, 1'b1, _0678_, _0679_ }, { _3376_, _3408_, _3372_, _3371_ });
  assign _3408_ = | (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4641|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4639" *) { _3407_[0], _3407_[1] };
  assign _3407_[0] = { dp2lut_Xinfo_4[17:16], dp2lut_Yinfo_4[17:16] } == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4641|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4639" *) 1'b1;
  assign _3407_[1] = { dp2lut_Xinfo_4[17:16], dp2lut_Yinfo_4[17:16] } == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4641|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4639" *) 2'b10;
  assign lut_X_sel[4] = int8_en ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4638" *) _0376_ : 1'b0;
  function [0:0] _7332_;
    input [0:0] a;
    input [3:0] b;
    input [3:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4626|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4621" *)
    (* parallel_case *)
    casez (s)
      4'b???1:
        _7332_ = b[0:0];
      4'b??1?:
        _7332_ = b[1:1];
      4'b?1??:
        _7332_ = b[2:2];
      4'b1???:
        _7332_ = b[3:3];
      default:
        _7332_ = a;
    endcase
  endfunction
  assign lut_X_sel[3] = _7332_(1'b0, { _0677_, 1'b1, _0678_, _0679_ }, { _3382_, _3410_, _3378_, _3377_ });
  assign _3410_ = | (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4623|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4621" *) { _3409_[0], _3409_[1] };
  assign _3409_[0] = { dp2lut_Xinfo_3[17:16], dp2lut_Yinfo_3[17:16] } == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4623|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4621" *) 1'b1;
  assign _3409_[1] = { dp2lut_Xinfo_3[17:16], dp2lut_Yinfo_3[17:16] } == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4623|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4621" *) 2'b10;
  function [0:0] _7336_;
    input [0:0] a;
    input [3:0] b;
    input [3:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4610|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4605" *)
    (* parallel_case *)
    casez (s)
      4'b???1:
        _7336_ = b[0:0];
      4'b??1?:
        _7336_ = b[1:1];
      4'b?1??:
        _7336_ = b[2:2];
      4'b1???:
        _7336_ = b[3:3];
      default:
        _7336_ = a;
    endcase
  endfunction
  assign lut_X_sel[2] = _7336_(1'b0, { _0677_, 1'b1, _0678_, _0679_ }, { _3388_, _3412_, _3384_, _3383_ });
  assign _3412_ = | (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4607|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4605" *) { _3411_[0], _3411_[1] };
  assign _3411_[0] = { dp2lut_Xinfo_2[17:16], dp2lut_Yinfo_2[17:16] } == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4607|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4605" *) 1'b1;
  assign _3411_[1] = { dp2lut_Xinfo_2[17:16], dp2lut_Yinfo_2[17:16] } == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4607|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4605" *) 2'b10;
  function [0:0] _7340_;
    input [0:0] a;
    input [3:0] b;
    input [3:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4594|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4589" *)
    (* parallel_case *)
    casez (s)
      4'b???1:
        _7340_ = b[0:0];
      4'b??1?:
        _7340_ = b[1:1];
      4'b?1??:
        _7340_ = b[2:2];
      4'b1???:
        _7340_ = b[3:3];
      default:
        _7340_ = a;
    endcase
  endfunction
  assign lut_X_sel[1] = _7340_(1'b0, { _0677_, 1'b1, _0678_, _0679_ }, { _3394_, _3414_, _3390_, _3389_ });
  assign _3414_ = | (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4591|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4589" *) { _3413_[0], _3413_[1] };
  assign _3413_[0] = { dp2lut_Xinfo_1[17:16], dp2lut_Yinfo_1[17:16] } == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4591|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4589" *) 1'b1;
  assign _3413_[1] = { dp2lut_Xinfo_1[17:16], dp2lut_Yinfo_1[17:16] } == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4591|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4589" *) 2'b10;
  function [0:0] _7344_;
    input [0:0] a;
    input [3:0] b;
    input [3:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4578|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4573" *)
    (* parallel_case *)
    casez (s)
      4'b???1:
        _7344_ = b[0:0];
      4'b??1?:
        _7344_ = b[1:1];
      4'b?1??:
        _7344_ = b[2:2];
      4'b1???:
        _7344_ = b[3:3];
      default:
        _7344_ = a;
    endcase
  endfunction
  assign lut_X_sel[0] = _7344_(1'b0, { _0677_, 1'b1, _0678_, _0679_ }, { _3400_, _3416_, _3396_, _3395_ });
  assign _3416_ = | (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4575|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4573" *) { _3415_[0], _3415_[1] };
  assign _3415_[0] = { dp2lut_Xinfo_0[17:16], dp2lut_Yinfo_0[17:16] } == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4575|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4573" *) 1'b1;
  assign _3415_[1] = { dp2lut_Xinfo_0[17:16], dp2lut_Yinfo_0[17:16] } == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4575|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4573" *) 2'b10;
  function [15:0] _7348_;
    input [15:0] a;
    input [4095:0] b;
    input [255:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4547|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4034" *)
    (* parallel_case *)
    casez (s)
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1:
        _7348_ = b[15:0];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?:
        _7348_ = b[31:16];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??:
        _7348_ = b[47:32];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???:
        _7348_ = b[63:48];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????:
        _7348_ = b[79:64];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????:
        _7348_ = b[95:80];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????:
        _7348_ = b[111:96];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????:
        _7348_ = b[127:112];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????:
        _7348_ = b[143:128];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????:
        _7348_ = b[159:144];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????:
        _7348_ = b[175:160];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????:
        _7348_ = b[191:176];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????:
        _7348_ = b[207:192];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????:
        _7348_ = b[223:208];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????:
        _7348_ = b[239:224];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????:
        _7348_ = b[255:240];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????:
        _7348_ = b[271:256];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????:
        _7348_ = b[287:272];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????:
        _7348_ = b[303:288];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????:
        _7348_ = b[319:304];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????:
        _7348_ = b[335:320];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????:
        _7348_ = b[351:336];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????:
        _7348_ = b[367:352];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????:
        _7348_ = b[383:368];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????:
        _7348_ = b[399:384];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????:
        _7348_ = b[415:400];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????:
        _7348_ = b[431:416];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????:
        _7348_ = b[447:432];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????:
        _7348_ = b[463:448];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????:
        _7348_ = b[479:464];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????:
        _7348_ = b[495:480];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????:
        _7348_ = b[511:496];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????:
        _7348_ = b[527:512];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????:
        _7348_ = b[543:528];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????:
        _7348_ = b[559:544];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????:
        _7348_ = b[575:560];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????:
        _7348_ = b[591:576];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????:
        _7348_ = b[607:592];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????:
        _7348_ = b[623:608];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????:
        _7348_ = b[639:624];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????:
        _7348_ = b[655:640];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????:
        _7348_ = b[671:656];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????:
        _7348_ = b[687:672];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????:
        _7348_ = b[703:688];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????:
        _7348_ = b[719:704];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????:
        _7348_ = b[735:720];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????:
        _7348_ = b[751:736];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????:
        _7348_ = b[767:752];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????:
        _7348_ = b[783:768];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????:
        _7348_ = b[799:784];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????:
        _7348_ = b[815:800];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????:
        _7348_ = b[831:816];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????:
        _7348_ = b[847:832];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????:
        _7348_ = b[863:848];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????:
        _7348_ = b[879:864];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????:
        _7348_ = b[895:880];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????:
        _7348_ = b[911:896];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????:
        _7348_ = b[927:912];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????:
        _7348_ = b[943:928];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????:
        _7348_ = b[959:944];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????:
        _7348_ = b[975:960];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????:
        _7348_ = b[991:976];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????:
        _7348_ = b[1007:992];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????:
        _7348_ = b[1023:1008];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????:
        _7348_ = b[1039:1024];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????:
        _7348_ = b[1055:1040];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????:
        _7348_ = b[1071:1056];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????:
        _7348_ = b[1087:1072];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????:
        _7348_ = b[1103:1088];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????:
        _7348_ = b[1119:1104];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????:
        _7348_ = b[1135:1120];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????:
        _7348_ = b[1151:1136];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????:
        _7348_ = b[1167:1152];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????:
        _7348_ = b[1183:1168];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????:
        _7348_ = b[1199:1184];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????:
        _7348_ = b[1215:1200];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????:
        _7348_ = b[1231:1216];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????:
        _7348_ = b[1247:1232];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????:
        _7348_ = b[1263:1248];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????:
        _7348_ = b[1279:1264];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????:
        _7348_ = b[1295:1280];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????:
        _7348_ = b[1311:1296];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????:
        _7348_ = b[1327:1312];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????:
        _7348_ = b[1343:1328];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????:
        _7348_ = b[1359:1344];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????:
        _7348_ = b[1375:1360];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????:
        _7348_ = b[1391:1376];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????:
        _7348_ = b[1407:1392];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????:
        _7348_ = b[1423:1408];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????:
        _7348_ = b[1439:1424];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????:
        _7348_ = b[1455:1440];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????:
        _7348_ = b[1471:1456];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????:
        _7348_ = b[1487:1472];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????:
        _7348_ = b[1503:1488];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????:
        _7348_ = b[1519:1504];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????:
        _7348_ = b[1535:1520];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????:
        _7348_ = b[1551:1536];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????:
        _7348_ = b[1567:1552];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????:
        _7348_ = b[1583:1568];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????:
        _7348_ = b[1599:1584];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????:
        _7348_ = b[1615:1600];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????:
        _7348_ = b[1631:1616];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????:
        _7348_ = b[1647:1632];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????:
        _7348_ = b[1663:1648];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _7348_ = b[1679:1664];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _7348_ = b[1695:1680];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _7348_ = b[1711:1696];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _7348_ = b[1727:1712];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _7348_ = b[1743:1728];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _7348_ = b[1759:1744];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _7348_ = b[1775:1760];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _7348_ = b[1791:1776];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _7348_ = b[1807:1792];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _7348_ = b[1823:1808];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _7348_ = b[1839:1824];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _7348_ = b[1855:1840];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _7348_ = b[1871:1856];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _7348_ = b[1887:1872];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _7348_ = b[1903:1888];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _7348_ = b[1919:1904];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _7348_ = b[1935:1920];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _7348_ = b[1951:1936];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _7348_ = b[1967:1952];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _7348_ = b[1983:1968];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _7348_ = b[1999:1984];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _7348_ = b[2015:2000];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _7348_ = b[2031:2016];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _7348_ = b[2047:2032];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _7348_ = b[2063:2048];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _7348_ = b[2079:2064];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _7348_ = b[2095:2080];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _7348_ = b[2111:2096];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _7348_ = b[2127:2112];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _7348_ = b[2143:2128];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _7348_ = b[2159:2144];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _7348_ = b[2175:2160];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _7348_ = b[2191:2176];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _7348_ = b[2207:2192];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _7348_ = b[2223:2208];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _7348_ = b[2239:2224];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _7348_ = b[2255:2240];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _7348_ = b[2271:2256];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _7348_ = b[2287:2272];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _7348_ = b[2303:2288];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _7348_ = b[2319:2304];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _7348_ = b[2335:2320];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _7348_ = b[2351:2336];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _7348_ = b[2367:2352];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _7348_ = b[2383:2368];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _7348_ = b[2399:2384];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _7348_ = b[2415:2400];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _7348_ = b[2431:2416];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _7348_ = b[2447:2432];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _7348_ = b[2463:2448];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _7348_ = b[2479:2464];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _7348_ = b[2495:2480];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _7348_ = b[2511:2496];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _7348_ = b[2527:2512];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _7348_ = b[2543:2528];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _7348_ = b[2559:2544];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _7348_ = b[2575:2560];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _7348_ = b[2591:2576];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _7348_ = b[2607:2592];
      256'b????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _7348_ = b[2623:2608];
      256'b???????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _7348_ = b[2639:2624];
      256'b??????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _7348_ = b[2655:2640];
      256'b?????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _7348_ = b[2671:2656];
      256'b????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _7348_ = b[2687:2672];
      256'b???????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _7348_ = b[2703:2688];
      256'b??????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _7348_ = b[2719:2704];
      256'b?????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _7348_ = b[2735:2720];
      256'b????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _7348_ = b[2751:2736];
      256'b???????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _7348_ = b[2767:2752];
      256'b??????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _7348_ = b[2783:2768];
      256'b?????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _7348_ = b[2799:2784];
      256'b????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _7348_ = b[2815:2800];
      256'b???????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _7348_ = b[2831:2816];
      256'b??????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _7348_ = b[2847:2832];
      256'b?????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _7348_ = b[2863:2848];
      256'b????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _7348_ = b[2879:2864];
      256'b???????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _7348_ = b[2895:2880];
      256'b??????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _7348_ = b[2911:2896];
      256'b?????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _7348_ = b[2927:2912];
      256'b????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _7348_ = b[2943:2928];
      256'b???????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _7348_ = b[2959:2944];
      256'b??????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _7348_ = b[2975:2960];
      256'b?????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _7348_ = b[2991:2976];
      256'b????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _7348_ = b[3007:2992];
      256'b???????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _7348_ = b[3023:3008];
      256'b??????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _7348_ = b[3039:3024];
      256'b?????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _7348_ = b[3055:3040];
      256'b????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _7348_ = b[3071:3056];
      256'b???????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _7348_ = b[3087:3072];
      256'b??????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _7348_ = b[3103:3088];
      256'b?????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _7348_ = b[3119:3104];
      256'b????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _7348_ = b[3135:3120];
      256'b???????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _7348_ = b[3151:3136];
      256'b??????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _7348_ = b[3167:3152];
      256'b?????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _7348_ = b[3183:3168];
      256'b????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _7348_ = b[3199:3184];
      256'b???????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _7348_ = b[3215:3200];
      256'b??????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _7348_ = b[3231:3216];
      256'b?????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _7348_ = b[3247:3232];
      256'b????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _7348_ = b[3263:3248];
      256'b???????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _7348_ = b[3279:3264];
      256'b??????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _7348_ = b[3295:3280];
      256'b?????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _7348_ = b[3311:3296];
      256'b????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _7348_ = b[3327:3312];
      256'b???????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _7348_ = b[3343:3328];
      256'b??????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _7348_ = b[3359:3344];
      256'b?????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _7348_ = b[3375:3360];
      256'b????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _7348_ = b[3391:3376];
      256'b???????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _7348_ = b[3407:3392];
      256'b??????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _7348_ = b[3423:3408];
      256'b?????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _7348_ = b[3439:3424];
      256'b????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _7348_ = b[3455:3440];
      256'b???????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _7348_ = b[3471:3456];
      256'b??????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _7348_ = b[3487:3472];
      256'b?????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _7348_ = b[3503:3488];
      256'b????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _7348_ = b[3519:3504];
      256'b???????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _7348_ = b[3535:3520];
      256'b??????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _7348_ = b[3551:3536];
      256'b?????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _7348_ = b[3567:3552];
      256'b????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _7348_ = b[3583:3568];
      256'b???????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _7348_ = b[3599:3584];
      256'b??????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _7348_ = b[3615:3600];
      256'b?????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _7348_ = b[3631:3616];
      256'b????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _7348_ = b[3647:3632];
      256'b???????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _7348_ = b[3663:3648];
      256'b??????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _7348_ = b[3679:3664];
      256'b?????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _7348_ = b[3695:3680];
      256'b????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _7348_ = b[3711:3696];
      256'b???????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _7348_ = b[3727:3712];
      256'b??????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _7348_ = b[3743:3728];
      256'b?????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _7348_ = b[3759:3744];
      256'b????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _7348_ = b[3775:3760];
      256'b???????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _7348_ = b[3791:3776];
      256'b??????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _7348_ = b[3807:3792];
      256'b?????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _7348_ = b[3823:3808];
      256'b????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _7348_ = b[3839:3824];
      256'b???????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _7348_ = b[3855:3840];
      256'b??????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _7348_ = b[3871:3856];
      256'b?????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _7348_ = b[3887:3872];
      256'b????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _7348_ = b[3903:3888];
      256'b???????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _7348_ = b[3919:3904];
      256'b??????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _7348_ = b[3935:3920];
      256'b?????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _7348_ = b[3951:3936];
      256'b????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _7348_ = b[3967:3952];
      256'b???????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _7348_ = b[3983:3968];
      256'b??????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _7348_ = b[3999:3984];
      256'b?????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _7348_ = b[4015:4000];
      256'b????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _7348_ = b[4031:4016];
      256'b???1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _7348_ = b[4047:4032];
      256'b??1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _7348_ = b[4063:4048];
      256'b?1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _7348_ = b[4079:4064];
      256'b1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _7348_ = b[4095:4080];
      default:
        _7348_ = a;
    endcase
  endfunction
  assign _0000_ = _7348_(density_reg0, { density_reg1, density_reg2, density_reg3, density_reg4, density_reg5, density_reg6, density_reg7, density_reg8, density_reg9, density_reg10, density_reg11, density_reg12, density_reg13, density_reg14, density_reg15, density_reg16, density_reg17, density_reg18, density_reg19, density_reg20, density_reg21, density_reg22, density_reg23, density_reg24, density_reg25, density_reg26, density_reg27, density_reg28, density_reg29, density_reg30, density_reg31, density_reg32, density_reg33, density_reg34, density_reg35, density_reg36, density_reg37, density_reg38, density_reg39, density_reg40, density_reg41, density_reg42, density_reg43, density_reg44, density_reg45, density_reg46, density_reg47, density_reg48, density_reg49, density_reg50, density_reg51, density_reg52, density_reg53, density_reg54, density_reg55, density_reg56, density_reg57, density_reg58, density_reg59, density_reg60, density_reg61, density_reg62, density_reg63, density_reg64, density_reg65, density_reg66, density_reg67, density_reg68, density_reg69, density_reg70, density_reg71, density_reg72, density_reg73, density_reg74, density_reg75, density_reg76, density_reg77, density_reg78, density_reg79, density_reg80, density_reg81, density_reg82, density_reg83, density_reg84, density_reg85, density_reg86, density_reg87, density_reg88, density_reg89, density_reg90, density_reg91, density_reg92, density_reg93, density_reg94, density_reg95, density_reg96, density_reg97, density_reg98, density_reg99, density_reg100, density_reg101, density_reg102, density_reg103, density_reg104, density_reg105, density_reg106, density_reg107, density_reg108, density_reg109, density_reg110, density_reg111, density_reg112, density_reg113, density_reg114, density_reg115, density_reg116, density_reg117, density_reg118, density_reg119, density_reg120, density_reg121, density_reg122, density_reg123, density_reg124, density_reg125, density_reg126, density_reg127, density_reg128, density_reg129, density_reg130, density_reg131, density_reg132, density_reg133, density_reg134, density_reg135, density_reg136, density_reg137, density_reg138, density_reg139, density_reg140, density_reg141, density_reg142, density_reg143, density_reg144, density_reg145, density_reg146, density_reg147, density_reg148, density_reg149, density_reg150, density_reg151, density_reg152, density_reg153, density_reg154, density_reg155, density_reg156, density_reg157, density_reg158, density_reg159, density_reg160, density_reg161, density_reg162, density_reg163, density_reg164, density_reg165, density_reg166, density_reg167, density_reg168, density_reg169, density_reg170, density_reg171, density_reg172, density_reg173, density_reg174, density_reg175, density_reg176, density_reg177, density_reg178, density_reg179, density_reg180, density_reg181, density_reg182, density_reg183, density_reg184, density_reg185, density_reg186, density_reg187, density_reg188, density_reg189, density_reg190, density_reg191, density_reg192, density_reg193, density_reg194, density_reg195, density_reg196, density_reg197, density_reg198, density_reg199, density_reg200, density_reg201, density_reg202, density_reg203, density_reg204, density_reg205, density_reg206, density_reg207, density_reg208, density_reg209, density_reg210, density_reg211, density_reg212, density_reg213, density_reg214, density_reg215, density_reg216, density_reg217, density_reg218, density_reg219, density_reg220, density_reg221, density_reg222, density_reg223, density_reg224, density_reg225, density_reg226, density_reg227, density_reg228, density_reg229, density_reg230, density_reg231, density_reg232, density_reg233, density_reg234, density_reg235, density_reg236, density_reg237, density_reg238, density_reg239, density_reg240, density_reg241, density_reg242, density_reg243, density_reg244, density_reg245, density_reg246, density_reg247, density_reg248, density_reg249, density_reg250, density_reg251, density_reg252, density_reg253, density_reg254, density_reg255, density_reg256 }, { _0452_, _0453_, _0454_, _0455_, _0456_, _0457_, _0458_, _0459_, _0460_, _0461_, _0462_, _0463_, _0464_, _0465_, _0466_, _0467_, _0468_, _0469_, _0470_, _0471_, _0472_, _0473_, _0474_, _0475_, _0476_, _0477_, _0478_, _0479_, _0480_, _0481_, _0482_, _0483_, _0419_, _0420_, _0421_, _0422_, _0423_, _0424_, _0425_, _0426_, _0427_, _0428_, _0429_, _0430_, _0431_, _0432_, _0433_, _0434_, _0435_, _0436_, _0437_, _0438_, _0439_, _0440_, _0441_, _0442_, _0443_, _0444_, _0445_, _0446_, _0447_, _0448_, _0449_, _0450_, _0484_, _0485_, _0486_, _0487_, _0488_, _0489_, _0490_, _0491_, _0492_, _0493_, _0494_, _0495_, _0496_, _0497_, _0498_, _0499_, _0500_, _0501_, _0502_, _0503_, _0504_, _0505_, _0506_, _0507_, _0508_, _0509_, _0510_, _0511_, _0512_, _0513_, _0514_, _0515_, _0516_, _0517_, _0518_, _0519_, _0520_, _0521_, _0522_, _0523_, _0524_, _0525_, _0526_, _0527_, _0528_, _0529_, _0530_, _0531_, _0532_, _0533_, _0534_, _0535_, _0536_, _0537_, _0538_, _0539_, _0540_, _0541_, _0542_, _0543_, _0544_, _0545_, _0546_, _0547_, _0548_, _0549_, _0550_, _0551_, _0552_, _0553_, _0554_, _0555_, _0556_, _0557_, _0558_, _0559_, _0560_, _0561_, _0562_, _0563_, _0564_, _0565_, _0566_, _0567_, _0568_, _0569_, _0570_, _0571_, _0572_, _0573_, _0574_, _0575_, _0576_, _0577_, _0578_, _0579_, _0580_, _0581_, _0582_, _0583_, _0584_, _0585_, _0586_, _0587_, _0588_, _0589_, _0590_, _0591_, _0592_, _0593_, _0594_, _0595_, _0596_, _0597_, _0598_, _0599_, _0600_, _0601_, _0602_, _0603_, _0604_, _0605_, _0606_, _0607_, _0608_, _0609_, _0610_, _0611_, _0612_, _0613_, _0614_, _0615_, _0616_, _0617_, _0618_, _0619_, _0620_, _0621_, _0622_, _0623_, _0624_, _0625_, _0626_, _0627_, _0628_, _0629_, _0630_, _0631_, _0632_, _0633_, _0634_, _0635_, _0636_, _0637_, _0638_, _0639_, _0640_, _0641_, _0642_, _0643_, _0644_, _0645_, _0646_, _0647_, _0648_, _0649_, _0650_, _0651_, _0652_, _0653_, _0654_, _0655_, _0656_, _0657_, _0658_, _0659_, _0660_, _0661_, _0662_, _0663_, _0664_, _0665_, _0666_, _0667_, _0668_, _0669_, _0670_, _0671_, _0672_, _0673_, _0674_, _0675_ });
  function [15:0] _7349_;
    input [15:0] a;
    input [1023:0] b;
    input [63:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4024|./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3895" *)
    (* parallel_case *)
    casez (s)
      64'b???????????????????????????????????????????????????????????????1:
        _7349_ = b[15:0];
      64'b??????????????????????????????????????????????????????????????1?:
        _7349_ = b[31:16];
      64'b?????????????????????????????????????????????????????????????1??:
        _7349_ = b[47:32];
      64'b????????????????????????????????????????????????????????????1???:
        _7349_ = b[63:48];
      64'b???????????????????????????????????????????????????????????1????:
        _7349_ = b[79:64];
      64'b??????????????????????????????????????????????????????????1?????:
        _7349_ = b[95:80];
      64'b?????????????????????????????????????????????????????????1??????:
        _7349_ = b[111:96];
      64'b????????????????????????????????????????????????????????1???????:
        _7349_ = b[127:112];
      64'b???????????????????????????????????????????????????????1????????:
        _7349_ = b[143:128];
      64'b??????????????????????????????????????????????????????1?????????:
        _7349_ = b[159:144];
      64'b?????????????????????????????????????????????????????1??????????:
        _7349_ = b[175:160];
      64'b????????????????????????????????????????????????????1???????????:
        _7349_ = b[191:176];
      64'b???????????????????????????????????????????????????1????????????:
        _7349_ = b[207:192];
      64'b??????????????????????????????????????????????????1?????????????:
        _7349_ = b[223:208];
      64'b?????????????????????????????????????????????????1??????????????:
        _7349_ = b[239:224];
      64'b????????????????????????????????????????????????1???????????????:
        _7349_ = b[255:240];
      64'b???????????????????????????????????????????????1????????????????:
        _7349_ = b[271:256];
      64'b??????????????????????????????????????????????1?????????????????:
        _7349_ = b[287:272];
      64'b?????????????????????????????????????????????1??????????????????:
        _7349_ = b[303:288];
      64'b????????????????????????????????????????????1???????????????????:
        _7349_ = b[319:304];
      64'b???????????????????????????????????????????1????????????????????:
        _7349_ = b[335:320];
      64'b??????????????????????????????????????????1?????????????????????:
        _7349_ = b[351:336];
      64'b?????????????????????????????????????????1??????????????????????:
        _7349_ = b[367:352];
      64'b????????????????????????????????????????1???????????????????????:
        _7349_ = b[383:368];
      64'b???????????????????????????????????????1????????????????????????:
        _7349_ = b[399:384];
      64'b??????????????????????????????????????1?????????????????????????:
        _7349_ = b[415:400];
      64'b?????????????????????????????????????1??????????????????????????:
        _7349_ = b[431:416];
      64'b????????????????????????????????????1???????????????????????????:
        _7349_ = b[447:432];
      64'b???????????????????????????????????1????????????????????????????:
        _7349_ = b[463:448];
      64'b??????????????????????????????????1?????????????????????????????:
        _7349_ = b[479:464];
      64'b?????????????????????????????????1??????????????????????????????:
        _7349_ = b[495:480];
      64'b????????????????????????????????1???????????????????????????????:
        _7349_ = b[511:496];
      64'b???????????????????????????????1????????????????????????????????:
        _7349_ = b[527:512];
      64'b??????????????????????????????1?????????????????????????????????:
        _7349_ = b[543:528];
      64'b?????????????????????????????1??????????????????????????????????:
        _7349_ = b[559:544];
      64'b????????????????????????????1???????????????????????????????????:
        _7349_ = b[575:560];
      64'b???????????????????????????1????????????????????????????????????:
        _7349_ = b[591:576];
      64'b??????????????????????????1?????????????????????????????????????:
        _7349_ = b[607:592];
      64'b?????????????????????????1??????????????????????????????????????:
        _7349_ = b[623:608];
      64'b????????????????????????1???????????????????????????????????????:
        _7349_ = b[639:624];
      64'b???????????????????????1????????????????????????????????????????:
        _7349_ = b[655:640];
      64'b??????????????????????1?????????????????????????????????????????:
        _7349_ = b[671:656];
      64'b?????????????????????1??????????????????????????????????????????:
        _7349_ = b[687:672];
      64'b????????????????????1???????????????????????????????????????????:
        _7349_ = b[703:688];
      64'b???????????????????1????????????????????????????????????????????:
        _7349_ = b[719:704];
      64'b??????????????????1?????????????????????????????????????????????:
        _7349_ = b[735:720];
      64'b?????????????????1??????????????????????????????????????????????:
        _7349_ = b[751:736];
      64'b????????????????1???????????????????????????????????????????????:
        _7349_ = b[767:752];
      64'b???????????????1????????????????????????????????????????????????:
        _7349_ = b[783:768];
      64'b??????????????1?????????????????????????????????????????????????:
        _7349_ = b[799:784];
      64'b?????????????1??????????????????????????????????????????????????:
        _7349_ = b[815:800];
      64'b????????????1???????????????????????????????????????????????????:
        _7349_ = b[831:816];
      64'b???????????1????????????????????????????????????????????????????:
        _7349_ = b[847:832];
      64'b??????????1?????????????????????????????????????????????????????:
        _7349_ = b[863:848];
      64'b?????????1??????????????????????????????????????????????????????:
        _7349_ = b[879:864];
      64'b????????1???????????????????????????????????????????????????????:
        _7349_ = b[895:880];
      64'b???????1????????????????????????????????????????????????????????:
        _7349_ = b[911:896];
      64'b??????1?????????????????????????????????????????????????????????:
        _7349_ = b[927:912];
      64'b?????1??????????????????????????????????????????????????????????:
        _7349_ = b[943:928];
      64'b????1???????????????????????????????????????????????????????????:
        _7349_ = b[959:944];
      64'b???1????????????????????????????????????????????????????????????:
        _7349_ = b[975:960];
      64'b??1?????????????????????????????????????????????????????????????:
        _7349_ = b[991:976];
      64'b?1??????????????????????????????????????????????????????????????:
        _7349_ = b[1007:992];
      64'b1???????????????????????????????????????????????????????????????:
        _7349_ = b[1023:1008];
      default:
        _7349_ = a;
    endcase
  endfunction
  assign _0310_ = _7349_(raw_reg0, { raw_reg1, raw_reg2, raw_reg3, raw_reg4, raw_reg5, raw_reg6, raw_reg7, raw_reg8, raw_reg9, raw_reg10, raw_reg11, raw_reg12, raw_reg13, raw_reg14, raw_reg15, raw_reg16, raw_reg17, raw_reg18, raw_reg19, raw_reg20, raw_reg21, raw_reg22, raw_reg23, raw_reg24, raw_reg25, raw_reg26, raw_reg27, raw_reg28, raw_reg29, raw_reg30, raw_reg31, raw_reg32, raw_reg33, raw_reg34, raw_reg35, raw_reg36, raw_reg37, raw_reg38, raw_reg39, raw_reg40, raw_reg41, raw_reg42, raw_reg43, raw_reg44, raw_reg45, raw_reg46, raw_reg47, raw_reg48, raw_reg49, raw_reg50, raw_reg51, raw_reg52, raw_reg53, raw_reg54, raw_reg55, raw_reg56, raw_reg57, raw_reg58, raw_reg59, raw_reg60, raw_reg61, raw_reg62, raw_reg63, raw_reg64 }, { _0452_, _0453_, _0454_, _0455_, _0456_, _0457_, _0458_, _0459_, _0460_, _0461_, _0462_, _0463_, _0464_, _0465_, _0466_, _0467_, _0468_, _0469_, _0470_, _0471_, _0472_, _0473_, _0474_, _0475_, _0476_, _0477_, _0478_, _0479_, _0480_, _0481_, _0482_, _0483_, _0419_, _0420_, _0421_, _0422_, _0423_, _0424_, _0425_, _0426_, _0427_, _0428_, _0429_, _0430_, _0431_, _0432_, _0433_, _0434_, _0435_, _0436_, _0437_, _0438_, _0439_, _0440_, _0441_, _0442_, _0443_, _0444_, _0445_, _0446_, _0447_, _0448_, _0449_, _0450_ });
  assign _3417_ = _0675_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3883" *) reg2dp_lut_data : density_reg256;
  assign _0174_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3882" *) _3417_ : density_reg256;
  assign _3418_ = _0674_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3873" *) reg2dp_lut_data : density_reg255;
  assign _0173_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3872" *) _3418_ : density_reg255;
  assign _3419_ = _0673_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3863" *) reg2dp_lut_data : density_reg254;
  assign _0172_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3862" *) _3419_ : density_reg254;
  assign _3420_ = _0672_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3853" *) reg2dp_lut_data : density_reg253;
  assign _0171_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3852" *) _3420_ : density_reg253;
  assign _3421_ = _0671_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3843" *) reg2dp_lut_data : density_reg252;
  assign _0170_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3842" *) _3421_ : density_reg252;
  assign _3422_ = _0670_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3833" *) reg2dp_lut_data : density_reg251;
  assign _0169_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3832" *) _3422_ : density_reg251;
  assign _3423_ = _0669_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3823" *) reg2dp_lut_data : density_reg250;
  assign _0168_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3822" *) _3423_ : density_reg250;
  assign _3424_ = _0668_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3813" *) reg2dp_lut_data : density_reg249;
  assign _0166_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3812" *) _3424_ : density_reg249;
  assign _3425_ = _0667_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3803" *) reg2dp_lut_data : density_reg248;
  assign _0165_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3802" *) _3425_ : density_reg248;
  assign _3426_ = _0666_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3793" *) reg2dp_lut_data : density_reg247;
  assign _0164_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3792" *) _3426_ : density_reg247;
  assign _3427_ = _0665_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3783" *) reg2dp_lut_data : density_reg246;
  assign _0163_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3782" *) _3427_ : density_reg246;
  assign _3428_ = _0664_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3773" *) reg2dp_lut_data : density_reg245;
  assign _0162_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3772" *) _3428_ : density_reg245;
  assign _3429_ = _0663_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3763" *) reg2dp_lut_data : density_reg244;
  assign _0161_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3762" *) _3429_ : density_reg244;
  assign _3430_ = _0662_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3753" *) reg2dp_lut_data : density_reg243;
  assign _0160_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3752" *) _3430_ : density_reg243;
  assign _3431_ = _0661_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3743" *) reg2dp_lut_data : density_reg242;
  assign _0159_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3742" *) _3431_ : density_reg242;
  assign _3432_ = _0660_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3733" *) reg2dp_lut_data : density_reg241;
  assign _0158_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3732" *) _3432_ : density_reg241;
  assign _3433_ = _0659_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3723" *) reg2dp_lut_data : density_reg240;
  assign _0157_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3722" *) _3433_ : density_reg240;
  assign _3434_ = _0658_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3713" *) reg2dp_lut_data : density_reg239;
  assign _0155_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3712" *) _3434_ : density_reg239;
  assign _3435_ = _0657_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3703" *) reg2dp_lut_data : density_reg238;
  assign _0154_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3702" *) _3435_ : density_reg238;
  assign _3436_ = _0656_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3693" *) reg2dp_lut_data : density_reg237;
  assign _0153_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3692" *) _3436_ : density_reg237;
  assign _3437_ = _0655_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3683" *) reg2dp_lut_data : density_reg236;
  assign _0152_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3682" *) _3437_ : density_reg236;
  assign _3438_ = _0654_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3673" *) reg2dp_lut_data : density_reg235;
  assign _0151_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3672" *) _3438_ : density_reg235;
  assign _3439_ = _0653_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3663" *) reg2dp_lut_data : density_reg234;
  assign _0150_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3662" *) _3439_ : density_reg234;
  assign _3440_ = _0652_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3653" *) reg2dp_lut_data : density_reg233;
  assign _0149_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3652" *) _3440_ : density_reg233;
  assign _3441_ = _0651_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3643" *) reg2dp_lut_data : density_reg232;
  assign _0148_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3642" *) _3441_ : density_reg232;
  assign _3442_ = _0650_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3633" *) reg2dp_lut_data : density_reg231;
  assign _0147_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3632" *) _3442_ : density_reg231;
  assign _3443_ = _0649_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3623" *) reg2dp_lut_data : density_reg230;
  assign _0146_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3622" *) _3443_ : density_reg230;
  assign _3444_ = _0648_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3613" *) reg2dp_lut_data : density_reg229;
  assign _0144_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3612" *) _3444_ : density_reg229;
  assign _3445_ = _0647_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3603" *) reg2dp_lut_data : density_reg228;
  assign _0143_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3602" *) _3445_ : density_reg228;
  assign _3446_ = _0646_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3593" *) reg2dp_lut_data : density_reg227;
  assign _0142_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3592" *) _3446_ : density_reg227;
  assign _3447_ = _0645_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3583" *) reg2dp_lut_data : density_reg226;
  assign _0141_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3582" *) _3447_ : density_reg226;
  assign _3448_ = _0644_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3573" *) reg2dp_lut_data : density_reg225;
  assign _0140_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3572" *) _3448_ : density_reg225;
  assign _3449_ = _0643_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3563" *) reg2dp_lut_data : density_reg224;
  assign _0139_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3562" *) _3449_ : density_reg224;
  assign _3450_ = _0642_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3553" *) reg2dp_lut_data : density_reg223;
  assign _0138_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3552" *) _3450_ : density_reg223;
  assign _3451_ = _0641_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3543" *) reg2dp_lut_data : density_reg222;
  assign _0137_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3542" *) _3451_ : density_reg222;
  assign _3452_ = _0640_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3533" *) reg2dp_lut_data : density_reg221;
  assign _0136_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3532" *) _3452_ : density_reg221;
  assign _3453_ = _0639_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3523" *) reg2dp_lut_data : density_reg220;
  assign _0135_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3522" *) _3453_ : density_reg220;
  assign _3454_ = _0638_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3513" *) reg2dp_lut_data : density_reg219;
  assign _0133_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3512" *) _3454_ : density_reg219;
  assign _3455_ = _0637_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3503" *) reg2dp_lut_data : density_reg218;
  assign _0132_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3502" *) _3455_ : density_reg218;
  assign _3456_ = _0636_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3493" *) reg2dp_lut_data : density_reg217;
  assign _0131_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3492" *) _3456_ : density_reg217;
  assign _3457_ = _0635_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3483" *) reg2dp_lut_data : density_reg216;
  assign _0130_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3482" *) _3457_ : density_reg216;
  assign _3458_ = _0634_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3473" *) reg2dp_lut_data : density_reg215;
  assign _0129_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3472" *) _3458_ : density_reg215;
  assign _3459_ = _0633_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3463" *) reg2dp_lut_data : density_reg214;
  assign _0128_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3462" *) _3459_ : density_reg214;
  assign _3460_ = _0632_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3453" *) reg2dp_lut_data : density_reg213;
  assign _0127_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3452" *) _3460_ : density_reg213;
  assign _3461_ = _0631_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3443" *) reg2dp_lut_data : density_reg212;
  assign _0126_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3442" *) _3461_ : density_reg212;
  assign _3462_ = _0630_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3433" *) reg2dp_lut_data : density_reg211;
  assign _0125_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3432" *) _3462_ : density_reg211;
  assign _3463_ = _0629_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3423" *) reg2dp_lut_data : density_reg210;
  assign _0124_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3422" *) _3463_ : density_reg210;
  assign _3464_ = _0628_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3413" *) reg2dp_lut_data : density_reg209;
  assign _0122_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3412" *) _3464_ : density_reg209;
  assign _3465_ = _0627_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3403" *) reg2dp_lut_data : density_reg208;
  assign _0121_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3402" *) _3465_ : density_reg208;
  assign _3466_ = _0626_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3393" *) reg2dp_lut_data : density_reg207;
  assign _0120_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3392" *) _3466_ : density_reg207;
  assign _3467_ = _0625_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3383" *) reg2dp_lut_data : density_reg206;
  assign _0119_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3382" *) _3467_ : density_reg206;
  assign _3468_ = _0624_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3373" *) reg2dp_lut_data : density_reg205;
  assign _0118_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3372" *) _3468_ : density_reg205;
  assign _3469_ = _0623_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3363" *) reg2dp_lut_data : density_reg204;
  assign _0117_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3362" *) _3469_ : density_reg204;
  assign _3470_ = _0622_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3353" *) reg2dp_lut_data : density_reg203;
  assign _0116_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3352" *) _3470_ : density_reg203;
  assign _3471_ = _0621_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3343" *) reg2dp_lut_data : density_reg202;
  assign _0115_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3342" *) _3471_ : density_reg202;
  assign _3472_ = _0620_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3333" *) reg2dp_lut_data : density_reg201;
  assign _0114_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3332" *) _3472_ : density_reg201;
  assign _3473_ = _0619_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3323" *) reg2dp_lut_data : density_reg200;
  assign _0113_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3322" *) _3473_ : density_reg200;
  assign _3474_ = _0618_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3313" *) reg2dp_lut_data : density_reg199;
  assign _0110_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3312" *) _3474_ : density_reg199;
  assign _3475_ = _0617_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3303" *) reg2dp_lut_data : density_reg198;
  assign _0109_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3302" *) _3475_ : density_reg198;
  assign _3476_ = _0616_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3293" *) reg2dp_lut_data : density_reg197;
  assign _0108_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3292" *) _3476_ : density_reg197;
  assign _3477_ = _0615_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3283" *) reg2dp_lut_data : density_reg196;
  assign _0107_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3282" *) _3477_ : density_reg196;
  assign _3478_ = _0614_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3273" *) reg2dp_lut_data : density_reg195;
  assign _0106_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3272" *) _3478_ : density_reg195;
  assign _3479_ = _0613_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3263" *) reg2dp_lut_data : density_reg194;
  assign _0105_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3262" *) _3479_ : density_reg194;
  assign _3480_ = _0612_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3253" *) reg2dp_lut_data : density_reg193;
  assign _0104_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3252" *) _3480_ : density_reg193;
  assign _3481_ = _0611_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3243" *) reg2dp_lut_data : density_reg192;
  assign _0103_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3242" *) _3481_ : density_reg192;
  assign _3482_ = _0610_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3233" *) reg2dp_lut_data : density_reg191;
  assign _0102_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3232" *) _3482_ : density_reg191;
  assign _3483_ = _0609_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3223" *) reg2dp_lut_data : density_reg190;
  assign _0101_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3222" *) _3483_ : density_reg190;
  assign _3484_ = _0608_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3213" *) reg2dp_lut_data : density_reg189;
  assign _0099_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3212" *) _3484_ : density_reg189;
  assign _3485_ = _0607_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3203" *) reg2dp_lut_data : density_reg188;
  assign _0098_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3202" *) _3485_ : density_reg188;
  assign _3486_ = _0606_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3193" *) reg2dp_lut_data : density_reg187;
  assign _0097_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3192" *) _3486_ : density_reg187;
  assign _3487_ = _0605_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3183" *) reg2dp_lut_data : density_reg186;
  assign _0096_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3182" *) _3487_ : density_reg186;
  assign _3488_ = _0604_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3173" *) reg2dp_lut_data : density_reg185;
  assign _0095_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3172" *) _3488_ : density_reg185;
  assign _3489_ = _0603_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3163" *) reg2dp_lut_data : density_reg184;
  assign _0094_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3162" *) _3489_ : density_reg184;
  assign _3490_ = _0602_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3153" *) reg2dp_lut_data : density_reg183;
  assign _0093_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3152" *) _3490_ : density_reg183;
  assign _3491_ = _0601_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3143" *) reg2dp_lut_data : density_reg182;
  assign _0092_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3142" *) _3491_ : density_reg182;
  assign _3492_ = _0600_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3133" *) reg2dp_lut_data : density_reg181;
  assign _0091_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3132" *) _3492_ : density_reg181;
  assign _3493_ = _0599_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3123" *) reg2dp_lut_data : density_reg180;
  assign _0090_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3122" *) _3493_ : density_reg180;
  assign _3494_ = _0598_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3113" *) reg2dp_lut_data : density_reg179;
  assign _0088_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3112" *) _3494_ : density_reg179;
  assign _3495_ = _0597_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3103" *) reg2dp_lut_data : density_reg178;
  assign _0087_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3102" *) _3495_ : density_reg178;
  assign _3496_ = _0596_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3093" *) reg2dp_lut_data : density_reg177;
  assign _0086_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3092" *) _3496_ : density_reg177;
  assign _3497_ = _0595_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3083" *) reg2dp_lut_data : density_reg176;
  assign _0085_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3082" *) _3497_ : density_reg176;
  assign _3498_ = _0594_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3073" *) reg2dp_lut_data : density_reg175;
  assign _0084_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3072" *) _3498_ : density_reg175;
  assign _3499_ = _0593_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3063" *) reg2dp_lut_data : density_reg174;
  assign _0083_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3062" *) _3499_ : density_reg174;
  assign _3500_ = _0592_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3053" *) reg2dp_lut_data : density_reg173;
  assign _0082_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3052" *) _3500_ : density_reg173;
  assign _3501_ = _0591_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3043" *) reg2dp_lut_data : density_reg172;
  assign _0081_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3042" *) _3501_ : density_reg172;
  assign _3502_ = _0590_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3033" *) reg2dp_lut_data : density_reg171;
  assign _0080_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3032" *) _3502_ : density_reg171;
  assign _3503_ = _0589_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3023" *) reg2dp_lut_data : density_reg170;
  assign _0079_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3022" *) _3503_ : density_reg170;
  assign _3504_ = _0588_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3013" *) reg2dp_lut_data : density_reg169;
  assign _0077_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3012" *) _3504_ : density_reg169;
  assign _3505_ = _0587_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3003" *) reg2dp_lut_data : density_reg168;
  assign _0076_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:3002" *) _3505_ : density_reg168;
  assign _3506_ = _0586_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2993" *) reg2dp_lut_data : density_reg167;
  assign _0075_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2992" *) _3506_ : density_reg167;
  assign _3507_ = _0585_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2983" *) reg2dp_lut_data : density_reg166;
  assign _0074_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2982" *) _3507_ : density_reg166;
  assign _3508_ = _0584_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2973" *) reg2dp_lut_data : density_reg165;
  assign _0073_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2972" *) _3508_ : density_reg165;
  assign _3509_ = _0583_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2963" *) reg2dp_lut_data : density_reg164;
  assign _0072_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2962" *) _3509_ : density_reg164;
  assign _3510_ = _0582_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2953" *) reg2dp_lut_data : density_reg163;
  assign _0071_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2952" *) _3510_ : density_reg163;
  assign _3511_ = _0581_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2943" *) reg2dp_lut_data : density_reg162;
  assign _0070_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2942" *) _3511_ : density_reg162;
  assign _3512_ = _0580_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2933" *) reg2dp_lut_data : density_reg161;
  assign _0069_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2932" *) _3512_ : density_reg161;
  assign _3513_ = _0579_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2923" *) reg2dp_lut_data : density_reg160;
  assign _0068_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2922" *) _3513_ : density_reg160;
  assign _3514_ = _0578_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2913" *) reg2dp_lut_data : density_reg159;
  assign _0066_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2912" *) _3514_ : density_reg159;
  assign _3515_ = _0577_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2903" *) reg2dp_lut_data : density_reg158;
  assign _0065_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2902" *) _3515_ : density_reg158;
  assign _3516_ = _0576_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2893" *) reg2dp_lut_data : density_reg157;
  assign _0064_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2892" *) _3516_ : density_reg157;
  assign _3517_ = _0575_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2883" *) reg2dp_lut_data : density_reg156;
  assign _0063_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2882" *) _3517_ : density_reg156;
  assign _3518_ = _0574_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2873" *) reg2dp_lut_data : density_reg155;
  assign _0062_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2872" *) _3518_ : density_reg155;
  assign _3519_ = _0573_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2863" *) reg2dp_lut_data : density_reg154;
  assign _0061_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2862" *) _3519_ : density_reg154;
  assign _3520_ = _0572_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2853" *) reg2dp_lut_data : density_reg153;
  assign _0060_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2852" *) _3520_ : density_reg153;
  assign _3521_ = _0571_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2843" *) reg2dp_lut_data : density_reg152;
  assign _0059_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2842" *) _3521_ : density_reg152;
  assign _3522_ = _0570_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2833" *) reg2dp_lut_data : density_reg151;
  assign _0058_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2832" *) _3522_ : density_reg151;
  assign _3523_ = _0569_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2823" *) reg2dp_lut_data : density_reg150;
  assign _0057_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2822" *) _3523_ : density_reg150;
  assign _3524_ = _0568_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2813" *) reg2dp_lut_data : density_reg149;
  assign _0055_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2812" *) _3524_ : density_reg149;
  assign _3525_ = _0567_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2803" *) reg2dp_lut_data : density_reg148;
  assign _0054_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2802" *) _3525_ : density_reg148;
  assign _3526_ = _0566_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2793" *) reg2dp_lut_data : density_reg147;
  assign _0053_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2792" *) _3526_ : density_reg147;
  assign _3527_ = _0565_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2783" *) reg2dp_lut_data : density_reg146;
  assign _0052_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2782" *) _3527_ : density_reg146;
  assign _3528_ = _0564_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2773" *) reg2dp_lut_data : density_reg145;
  assign _0051_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2772" *) _3528_ : density_reg145;
  assign _3529_ = _0563_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2763" *) reg2dp_lut_data : density_reg144;
  assign _0050_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2762" *) _3529_ : density_reg144;
  assign _3530_ = _0562_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2753" *) reg2dp_lut_data : density_reg143;
  assign _0049_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2752" *) _3530_ : density_reg143;
  assign _3531_ = _0561_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2743" *) reg2dp_lut_data : density_reg142;
  assign _0048_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2742" *) _3531_ : density_reg142;
  assign _3532_ = _0560_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2733" *) reg2dp_lut_data : density_reg141;
  assign _0047_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2732" *) _3532_ : density_reg141;
  assign _3533_ = _0559_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2723" *) reg2dp_lut_data : density_reg140;
  assign _0046_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2722" *) _3533_ : density_reg140;
  assign _3534_ = _0558_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2713" *) reg2dp_lut_data : density_reg139;
  assign _0044_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2712" *) _3534_ : density_reg139;
  assign _3535_ = _0557_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2703" *) reg2dp_lut_data : density_reg138;
  assign _0043_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2702" *) _3535_ : density_reg138;
  assign _3536_ = _0556_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2693" *) reg2dp_lut_data : density_reg137;
  assign _0042_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2692" *) _3536_ : density_reg137;
  assign _3537_ = _0555_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2683" *) reg2dp_lut_data : density_reg136;
  assign _0041_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2682" *) _3537_ : density_reg136;
  assign _3538_ = _0554_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2673" *) reg2dp_lut_data : density_reg135;
  assign _0040_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2672" *) _3538_ : density_reg135;
  assign _3539_ = _0553_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2663" *) reg2dp_lut_data : density_reg134;
  assign _0039_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2662" *) _3539_ : density_reg134;
  assign _3540_ = _0552_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2653" *) reg2dp_lut_data : density_reg133;
  assign _0038_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2652" *) _3540_ : density_reg133;
  assign _3541_ = _0551_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2643" *) reg2dp_lut_data : density_reg132;
  assign _0037_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2642" *) _3541_ : density_reg132;
  assign _3542_ = _0550_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2633" *) reg2dp_lut_data : density_reg131;
  assign _0036_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2632" *) _3542_ : density_reg131;
  assign _3543_ = _0549_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2623" *) reg2dp_lut_data : density_reg130;
  assign _0035_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2622" *) _3543_ : density_reg130;
  assign _3544_ = _0548_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2613" *) reg2dp_lut_data : density_reg129;
  assign _0033_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2612" *) _3544_ : density_reg129;
  assign _3545_ = _0547_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2603" *) reg2dp_lut_data : density_reg128;
  assign _0032_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2602" *) _3545_ : density_reg128;
  assign _3546_ = _0546_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2593" *) reg2dp_lut_data : density_reg127;
  assign _0031_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2592" *) _3546_ : density_reg127;
  assign _3547_ = _0545_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2583" *) reg2dp_lut_data : density_reg126;
  assign _0030_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2582" *) _3547_ : density_reg126;
  assign _3548_ = _0544_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2573" *) reg2dp_lut_data : density_reg125;
  assign _0029_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2572" *) _3548_ : density_reg125;
  assign _3549_ = _0543_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2563" *) reg2dp_lut_data : density_reg124;
  assign _0028_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2562" *) _3549_ : density_reg124;
  assign _3550_ = _0542_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2553" *) reg2dp_lut_data : density_reg123;
  assign _0027_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2552" *) _3550_ : density_reg123;
  assign _3551_ = _0541_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2543" *) reg2dp_lut_data : density_reg122;
  assign _0026_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2542" *) _3551_ : density_reg122;
  assign _3552_ = _0540_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2533" *) reg2dp_lut_data : density_reg121;
  assign _0025_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2532" *) _3552_ : density_reg121;
  assign _3553_ = _0539_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2523" *) reg2dp_lut_data : density_reg120;
  assign _0024_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2522" *) _3553_ : density_reg120;
  assign _3554_ = _0538_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2513" *) reg2dp_lut_data : density_reg119;
  assign _0022_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2512" *) _3554_ : density_reg119;
  assign _3555_ = _0537_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2503" *) reg2dp_lut_data : density_reg118;
  assign _0021_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2502" *) _3555_ : density_reg118;
  assign _3556_ = _0536_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2493" *) reg2dp_lut_data : density_reg117;
  assign _0020_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2492" *) _3556_ : density_reg117;
  assign _3557_ = _0535_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2483" *) reg2dp_lut_data : density_reg116;
  assign _0019_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2482" *) _3557_ : density_reg116;
  assign _3558_ = _0534_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2473" *) reg2dp_lut_data : density_reg115;
  assign _0018_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2472" *) _3558_ : density_reg115;
  assign _3559_ = _0533_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2463" *) reg2dp_lut_data : density_reg114;
  assign _0017_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2462" *) _3559_ : density_reg114;
  assign _3560_ = _0532_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2453" *) reg2dp_lut_data : density_reg113;
  assign _0016_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2452" *) _3560_ : density_reg113;
  assign _3561_ = _0531_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2443" *) reg2dp_lut_data : density_reg112;
  assign _0015_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2442" *) _3561_ : density_reg112;
  assign _3562_ = _0530_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2433" *) reg2dp_lut_data : density_reg111;
  assign _0014_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2432" *) _3562_ : density_reg111;
  assign _3563_ = _0529_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2423" *) reg2dp_lut_data : density_reg110;
  assign _0013_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2422" *) _3563_ : density_reg110;
  assign _3564_ = _0528_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2413" *) reg2dp_lut_data : density_reg109;
  assign _0011_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2412" *) _3564_ : density_reg109;
  assign _3565_ = _0527_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2403" *) reg2dp_lut_data : density_reg108;
  assign _0010_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2402" *) _3565_ : density_reg108;
  assign _3566_ = _0526_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2393" *) reg2dp_lut_data : density_reg107;
  assign _0009_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2392" *) _3566_ : density_reg107;
  assign _3567_ = _0525_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2383" *) reg2dp_lut_data : density_reg106;
  assign _0008_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2382" *) _3567_ : density_reg106;
  assign _3568_ = _0524_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2373" *) reg2dp_lut_data : density_reg105;
  assign _0007_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2372" *) _3568_ : density_reg105;
  assign _3569_ = _0523_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2363" *) reg2dp_lut_data : density_reg104;
  assign _0006_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2362" *) _3569_ : density_reg104;
  assign _3570_ = _0522_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2353" *) reg2dp_lut_data : density_reg103;
  assign _0005_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2352" *) _3570_ : density_reg103;
  assign _3571_ = _0521_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2343" *) reg2dp_lut_data : density_reg102;
  assign _0004_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2342" *) _3571_ : density_reg102;
  assign _3572_ = _0520_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2333" *) reg2dp_lut_data : density_reg101;
  assign _0003_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2332" *) _3572_ : density_reg101;
  assign _3573_ = _0519_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2323" *) reg2dp_lut_data : density_reg100;
  assign _0002_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2322" *) _3573_ : density_reg100;
  assign _3574_ = _0518_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2313" *) reg2dp_lut_data : density_reg99;
  assign _0256_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2312" *) _3574_ : density_reg99;
  assign _3575_ = _0517_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2303" *) reg2dp_lut_data : density_reg98;
  assign _0255_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2302" *) _3575_ : density_reg98;
  assign _3576_ = _0516_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2293" *) reg2dp_lut_data : density_reg97;
  assign _0254_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2292" *) _3576_ : density_reg97;
  assign _3577_ = _0515_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2283" *) reg2dp_lut_data : density_reg96;
  assign _0253_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2282" *) _3577_ : density_reg96;
  assign _3578_ = _0514_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2273" *) reg2dp_lut_data : density_reg95;
  assign _0252_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2272" *) _3578_ : density_reg95;
  assign _3579_ = _0513_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2263" *) reg2dp_lut_data : density_reg94;
  assign _0251_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2262" *) _3579_ : density_reg94;
  assign _3580_ = _0512_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2253" *) reg2dp_lut_data : density_reg93;
  assign _0250_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2252" *) _3580_ : density_reg93;
  assign _3581_ = _0511_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2243" *) reg2dp_lut_data : density_reg92;
  assign _0249_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2242" *) _3581_ : density_reg92;
  assign _3582_ = _0510_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2233" *) reg2dp_lut_data : density_reg91;
  assign _0248_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2232" *) _3582_ : density_reg91;
  assign _3583_ = _0509_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2223" *) reg2dp_lut_data : density_reg90;
  assign _0247_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2222" *) _3583_ : density_reg90;
  assign _3584_ = _0508_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2213" *) reg2dp_lut_data : density_reg89;
  assign _0245_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2212" *) _3584_ : density_reg89;
  assign _3585_ = _0507_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2203" *) reg2dp_lut_data : density_reg88;
  assign _0244_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2202" *) _3585_ : density_reg88;
  assign _3586_ = _0506_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2193" *) reg2dp_lut_data : density_reg87;
  assign _0243_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2192" *) _3586_ : density_reg87;
  assign _3587_ = _0505_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2183" *) reg2dp_lut_data : density_reg86;
  assign _0242_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2182" *) _3587_ : density_reg86;
  assign _3588_ = _0504_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2173" *) reg2dp_lut_data : density_reg85;
  assign _0241_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2172" *) _3588_ : density_reg85;
  assign _3589_ = _0503_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2163" *) reg2dp_lut_data : density_reg84;
  assign _0240_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2162" *) _3589_ : density_reg84;
  assign _3590_ = _0502_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2153" *) reg2dp_lut_data : density_reg83;
  assign _0239_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2152" *) _3590_ : density_reg83;
  assign _3591_ = _0501_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2143" *) reg2dp_lut_data : density_reg82;
  assign _0238_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2142" *) _3591_ : density_reg82;
  assign _3592_ = _0500_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2133" *) reg2dp_lut_data : density_reg81;
  assign _0237_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2132" *) _3592_ : density_reg81;
  assign _3593_ = _0499_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2123" *) reg2dp_lut_data : density_reg80;
  assign _0236_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2122" *) _3593_ : density_reg80;
  assign _3594_ = _0498_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2113" *) reg2dp_lut_data : density_reg79;
  assign _0234_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2112" *) _3594_ : density_reg79;
  assign _3595_ = _0497_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2103" *) reg2dp_lut_data : density_reg78;
  assign _0233_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2102" *) _3595_ : density_reg78;
  assign _3596_ = _0496_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2093" *) reg2dp_lut_data : density_reg77;
  assign _0232_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2092" *) _3596_ : density_reg77;
  assign _3597_ = _0495_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2083" *) reg2dp_lut_data : density_reg76;
  assign _0231_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2082" *) _3597_ : density_reg76;
  assign _3598_ = _0494_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2073" *) reg2dp_lut_data : density_reg75;
  assign _0230_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2072" *) _3598_ : density_reg75;
  assign _3599_ = _0493_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2063" *) reg2dp_lut_data : density_reg74;
  assign _0229_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2062" *) _3599_ : density_reg74;
  assign _3600_ = _0492_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2053" *) reg2dp_lut_data : density_reg73;
  assign _0228_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2052" *) _3600_ : density_reg73;
  assign _3601_ = _0491_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2043" *) reg2dp_lut_data : density_reg72;
  assign _0227_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2042" *) _3601_ : density_reg72;
  assign _3602_ = _0490_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2033" *) reg2dp_lut_data : density_reg71;
  assign _0226_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2032" *) _3602_ : density_reg71;
  assign _3603_ = _0489_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2023" *) reg2dp_lut_data : density_reg70;
  assign _0225_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2022" *) _3603_ : density_reg70;
  assign _3604_ = _0488_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2013" *) reg2dp_lut_data : density_reg69;
  assign _0223_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2012" *) _3604_ : density_reg69;
  assign _3605_ = _0487_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2003" *) reg2dp_lut_data : density_reg68;
  assign _0222_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:2002" *) _3605_ : density_reg68;
  assign _3606_ = _0486_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1993" *) reg2dp_lut_data : density_reg67;
  assign _0221_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1992" *) _3606_ : density_reg67;
  assign _3607_ = _0485_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1983" *) reg2dp_lut_data : density_reg66;
  assign _0220_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1982" *) _3607_ : density_reg66;
  assign _3608_ = _0484_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1973" *) reg2dp_lut_data : density_reg65;
  assign _0219_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1972" *) _3608_ : density_reg65;
  assign _3609_ = _0450_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1963" *) reg2dp_lut_data : density_reg64;
  assign _0218_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1962" *) _3609_ : density_reg64;
  assign _3610_ = _0449_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1953" *) reg2dp_lut_data : density_reg63;
  assign _0217_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1952" *) _3610_ : density_reg63;
  assign _3611_ = _0448_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1943" *) reg2dp_lut_data : density_reg62;
  assign _0216_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1942" *) _3611_ : density_reg62;
  assign _3612_ = _0447_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1933" *) reg2dp_lut_data : density_reg61;
  assign _0215_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1932" *) _3612_ : density_reg61;
  assign _3613_ = _0446_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1923" *) reg2dp_lut_data : density_reg60;
  assign _0214_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1922" *) _3613_ : density_reg60;
  assign _3614_ = _0445_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1913" *) reg2dp_lut_data : density_reg59;
  assign _0212_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1912" *) _3614_ : density_reg59;
  assign _3615_ = _0444_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1903" *) reg2dp_lut_data : density_reg58;
  assign _0211_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1902" *) _3615_ : density_reg58;
  assign _3616_ = _0443_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1893" *) reg2dp_lut_data : density_reg57;
  assign _0210_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1892" *) _3616_ : density_reg57;
  assign _3617_ = _0442_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1883" *) reg2dp_lut_data : density_reg56;
  assign _0209_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1882" *) _3617_ : density_reg56;
  assign _3618_ = _0441_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1873" *) reg2dp_lut_data : density_reg55;
  assign _0208_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1872" *) _3618_ : density_reg55;
  assign _3619_ = _0440_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1863" *) reg2dp_lut_data : density_reg54;
  assign _0207_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1862" *) _3619_ : density_reg54;
  assign _3620_ = _0439_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1853" *) reg2dp_lut_data : density_reg53;
  assign _0206_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1852" *) _3620_ : density_reg53;
  assign _3621_ = _0438_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1843" *) reg2dp_lut_data : density_reg52;
  assign _0205_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1842" *) _3621_ : density_reg52;
  assign _3622_ = _0437_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1833" *) reg2dp_lut_data : density_reg51;
  assign _0204_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1832" *) _3622_ : density_reg51;
  assign _3623_ = _0436_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1823" *) reg2dp_lut_data : density_reg50;
  assign _0203_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1822" *) _3623_ : density_reg50;
  assign _3624_ = _0435_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1813" *) reg2dp_lut_data : density_reg49;
  assign _0201_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1812" *) _3624_ : density_reg49;
  assign _3625_ = _0434_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1803" *) reg2dp_lut_data : density_reg48;
  assign _0200_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1802" *) _3625_ : density_reg48;
  assign _3626_ = _0433_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1793" *) reg2dp_lut_data : density_reg47;
  assign _0199_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1792" *) _3626_ : density_reg47;
  assign _3627_ = _0432_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1783" *) reg2dp_lut_data : density_reg46;
  assign _0198_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1782" *) _3627_ : density_reg46;
  assign _3628_ = _0431_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1773" *) reg2dp_lut_data : density_reg45;
  assign _0197_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1772" *) _3628_ : density_reg45;
  assign _3629_ = _0430_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1763" *) reg2dp_lut_data : density_reg44;
  assign _0196_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1762" *) _3629_ : density_reg44;
  assign _3630_ = _0429_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1753" *) reg2dp_lut_data : density_reg43;
  assign _0195_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1752" *) _3630_ : density_reg43;
  assign _3631_ = _0428_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1743" *) reg2dp_lut_data : density_reg42;
  assign _0194_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1742" *) _3631_ : density_reg42;
  assign _3632_ = _0427_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1733" *) reg2dp_lut_data : density_reg41;
  assign _0193_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1732" *) _3632_ : density_reg41;
  assign _3633_ = _0426_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1723" *) reg2dp_lut_data : density_reg40;
  assign _0192_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1722" *) _3633_ : density_reg40;
  assign _3634_ = _0425_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1713" *) reg2dp_lut_data : density_reg39;
  assign _0190_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1712" *) _3634_ : density_reg39;
  assign _3635_ = _0424_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1703" *) reg2dp_lut_data : density_reg38;
  assign _0189_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1702" *) _3635_ : density_reg38;
  assign _3636_ = _0423_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1693" *) reg2dp_lut_data : density_reg37;
  assign _0188_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1692" *) _3636_ : density_reg37;
  assign _3637_ = _0422_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1683" *) reg2dp_lut_data : density_reg36;
  assign _0187_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1682" *) _3637_ : density_reg36;
  assign _3638_ = _0421_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1673" *) reg2dp_lut_data : density_reg35;
  assign _0186_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1672" *) _3638_ : density_reg35;
  assign _3639_ = _0420_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1663" *) reg2dp_lut_data : density_reg34;
  assign _0185_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1662" *) _3639_ : density_reg34;
  assign _3640_ = _0419_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1653" *) reg2dp_lut_data : density_reg33;
  assign _0184_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1652" *) _3640_ : density_reg33;
  assign _3641_ = _0483_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1643" *) reg2dp_lut_data : density_reg32;
  assign _0183_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1642" *) _3641_ : density_reg32;
  assign _3642_ = _0482_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1633" *) reg2dp_lut_data : density_reg31;
  assign _0182_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1632" *) _3642_ : density_reg31;
  assign _3643_ = _0481_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1623" *) reg2dp_lut_data : density_reg30;
  assign _0181_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1622" *) _3643_ : density_reg30;
  assign _3644_ = _0480_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1613" *) reg2dp_lut_data : density_reg29;
  assign _0179_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1612" *) _3644_ : density_reg29;
  assign _3645_ = _0479_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1603" *) reg2dp_lut_data : density_reg28;
  assign _0178_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1602" *) _3645_ : density_reg28;
  assign _3646_ = _0478_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1593" *) reg2dp_lut_data : density_reg27;
  assign _0177_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1592" *) _3646_ : density_reg27;
  assign _3647_ = _0477_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1583" *) reg2dp_lut_data : density_reg26;
  assign _0176_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1582" *) _3647_ : density_reg26;
  assign _3648_ = _0476_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1573" *) reg2dp_lut_data : density_reg25;
  assign _0175_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1572" *) _3648_ : density_reg25;
  assign _3649_ = _0475_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1563" *) reg2dp_lut_data : density_reg24;
  assign _0167_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1562" *) _3649_ : density_reg24;
  assign _3650_ = _0474_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1553" *) reg2dp_lut_data : density_reg23;
  assign _0156_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1552" *) _3650_ : density_reg23;
  assign _3651_ = _0473_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1543" *) reg2dp_lut_data : density_reg22;
  assign _0145_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1542" *) _3651_ : density_reg22;
  assign _3652_ = _0472_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1533" *) reg2dp_lut_data : density_reg21;
  assign _0134_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1532" *) _3652_ : density_reg21;
  assign _3653_ = _0471_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1523" *) reg2dp_lut_data : density_reg20;
  assign _0123_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1522" *) _3653_ : density_reg20;
  assign _3654_ = _0470_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1513" *) reg2dp_lut_data : density_reg19;
  assign _0111_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1512" *) _3654_ : density_reg19;
  assign _3655_ = _0469_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1503" *) reg2dp_lut_data : density_reg18;
  assign _0100_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1502" *) _3655_ : density_reg18;
  assign _3656_ = _0468_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1493" *) reg2dp_lut_data : density_reg17;
  assign _0089_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1492" *) _3656_ : density_reg17;
  assign _3657_ = _0467_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1483" *) reg2dp_lut_data : density_reg16;
  assign _0078_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1482" *) _3657_ : density_reg16;
  assign _3658_ = _0466_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1473" *) reg2dp_lut_data : density_reg15;
  assign _0067_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1472" *) _3658_ : density_reg15;
  assign _3659_ = _0465_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1463" *) reg2dp_lut_data : density_reg14;
  assign _0056_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1462" *) _3659_ : density_reg14;
  assign _3660_ = _0464_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1453" *) reg2dp_lut_data : density_reg13;
  assign _0045_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1452" *) _3660_ : density_reg13;
  assign _3661_ = _0463_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1443" *) reg2dp_lut_data : density_reg12;
  assign _0034_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1442" *) _3661_ : density_reg12;
  assign _3662_ = _0462_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1433" *) reg2dp_lut_data : density_reg11;
  assign _0023_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1432" *) _3662_ : density_reg11;
  assign _3663_ = _0461_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1423" *) reg2dp_lut_data : density_reg10;
  assign _0012_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1422" *) _3663_ : density_reg10;
  assign _3664_ = _0460_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1413" *) reg2dp_lut_data : density_reg9;
  assign _0257_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1412" *) _3664_ : density_reg9;
  assign _3665_ = _0459_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1403" *) reg2dp_lut_data : density_reg8;
  assign _0246_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1402" *) _3665_ : density_reg8;
  assign _3666_ = _0458_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1393" *) reg2dp_lut_data : density_reg7;
  assign _0235_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1392" *) _3666_ : density_reg7;
  assign _3667_ = _0457_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1383" *) reg2dp_lut_data : density_reg6;
  assign _0224_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1382" *) _3667_ : density_reg6;
  assign _3668_ = _0456_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1373" *) reg2dp_lut_data : density_reg5;
  assign _0213_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1372" *) _3668_ : density_reg5;
  assign _3669_ = _0455_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1363" *) reg2dp_lut_data : density_reg4;
  assign _0202_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1362" *) _3669_ : density_reg4;
  assign _3670_ = _0454_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1353" *) reg2dp_lut_data : density_reg3;
  assign _0191_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1352" *) _3670_ : density_reg3;
  assign _3671_ = _0453_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1343" *) reg2dp_lut_data : density_reg2;
  assign _0180_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1342" *) _3671_ : density_reg2;
  assign _3672_ = _0452_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1333" *) reg2dp_lut_data : density_reg1;
  assign _0112_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1332" *) _3672_ : density_reg1;
  assign _3673_ = _0451_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1323" *) reg2dp_lut_data : density_reg0;
  assign _0001_ = _0389_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1322" *) _3673_ : density_reg0;
  assign _3674_ = _0450_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1312" *) reg2dp_lut_data : raw_reg64;
  assign _0371_ = _0384_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1311" *) _3674_ : raw_reg64;
  assign _3675_ = _0449_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1302" *) reg2dp_lut_data : raw_reg63;
  assign _0370_ = _0384_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1301" *) _3675_ : raw_reg63;
  assign _3676_ = _0448_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1292" *) reg2dp_lut_data : raw_reg62;
  assign _0369_ = _0384_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1291" *) _3676_ : raw_reg62;
  assign _3677_ = _0447_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1282" *) reg2dp_lut_data : raw_reg61;
  assign _0368_ = _0384_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1281" *) _3677_ : raw_reg61;
  assign _3678_ = _0446_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1272" *) reg2dp_lut_data : raw_reg60;
  assign _0367_ = _0384_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1271" *) _3678_ : raw_reg60;
  assign _3679_ = _0445_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1262" *) reg2dp_lut_data : raw_reg59;
  assign _0365_ = _0384_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1261" *) _3679_ : raw_reg59;
  assign _3680_ = _0444_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1252" *) reg2dp_lut_data : raw_reg58;
  assign _0364_ = _0384_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1251" *) _3680_ : raw_reg58;
  assign _3681_ = _0443_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1242" *) reg2dp_lut_data : raw_reg57;
  assign _0363_ = _0384_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1241" *) _3681_ : raw_reg57;
  assign _3682_ = _0442_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1232" *) reg2dp_lut_data : raw_reg56;
  assign _0362_ = _0384_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1231" *) _3682_ : raw_reg56;
  assign _3683_ = _0441_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1222" *) reg2dp_lut_data : raw_reg55;
  assign _0361_ = _0384_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1221" *) _3683_ : raw_reg55;
  assign _3684_ = _0440_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1212" *) reg2dp_lut_data : raw_reg54;
  assign _0360_ = _0384_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1211" *) _3684_ : raw_reg54;
  assign _3685_ = _0439_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1202" *) reg2dp_lut_data : raw_reg53;
  assign _0359_ = _0384_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1201" *) _3685_ : raw_reg53;
  assign _3686_ = _0438_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1192" *) reg2dp_lut_data : raw_reg52;
  assign _0358_ = _0384_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1191" *) _3686_ : raw_reg52;
  assign _3687_ = _0437_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1182" *) reg2dp_lut_data : raw_reg51;
  assign _0357_ = _0384_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1181" *) _3687_ : raw_reg51;
  assign _3688_ = _0436_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1172" *) reg2dp_lut_data : raw_reg50;
  assign _0356_ = _0384_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1171" *) _3688_ : raw_reg50;
  assign _3689_ = _0435_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1162" *) reg2dp_lut_data : raw_reg49;
  assign _0354_ = _0384_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1161" *) _3689_ : raw_reg49;
  assign _3690_ = _0434_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1152" *) reg2dp_lut_data : raw_reg48;
  assign _0353_ = _0384_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1151" *) _3690_ : raw_reg48;
  assign _3691_ = _0433_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1142" *) reg2dp_lut_data : raw_reg47;
  assign _0352_ = _0384_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1141" *) _3691_ : raw_reg47;
  assign _3692_ = _0432_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1132" *) reg2dp_lut_data : raw_reg46;
  assign _0351_ = _0384_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1131" *) _3692_ : raw_reg46;
  assign _3693_ = _0431_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1122" *) reg2dp_lut_data : raw_reg45;
  assign _0350_ = _0384_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1121" *) _3693_ : raw_reg45;
  assign _3694_ = _0430_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1112" *) reg2dp_lut_data : raw_reg44;
  assign _0349_ = _0384_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1111" *) _3694_ : raw_reg44;
  assign _3695_ = _0429_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1102" *) reg2dp_lut_data : raw_reg43;
  assign _0348_ = _0384_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1101" *) _3695_ : raw_reg43;
  assign _3696_ = _0428_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1092" *) reg2dp_lut_data : raw_reg42;
  assign _0347_ = _0384_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1091" *) _3696_ : raw_reg42;
  assign _3697_ = _0427_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1082" *) reg2dp_lut_data : raw_reg41;
  assign _0346_ = _0384_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1081" *) _3697_ : raw_reg41;
  assign _3698_ = _0426_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1072" *) reg2dp_lut_data : raw_reg40;
  assign _0345_ = _0384_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1071" *) _3698_ : raw_reg40;
  assign _3699_ = _0425_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1062" *) reg2dp_lut_data : raw_reg39;
  assign _0343_ = _0384_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1061" *) _3699_ : raw_reg39;
  assign _3700_ = _0424_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1052" *) reg2dp_lut_data : raw_reg38;
  assign _0342_ = _0384_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1051" *) _3700_ : raw_reg38;
  assign _3701_ = _0423_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1042" *) reg2dp_lut_data : raw_reg37;
  assign _0341_ = _0384_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1041" *) _3701_ : raw_reg37;
  assign _3702_ = _0422_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1032" *) reg2dp_lut_data : raw_reg36;
  assign _0340_ = _0384_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1031" *) _3702_ : raw_reg36;
  assign _3703_ = _0421_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1022" *) reg2dp_lut_data : raw_reg35;
  assign _0339_ = _0384_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1021" *) _3703_ : raw_reg35;
  assign _3704_ = _0420_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1012" *) reg2dp_lut_data : raw_reg34;
  assign _0338_ = _0384_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1011" *) _3704_ : raw_reg34;
  assign _3705_ = _0419_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1002" *) reg2dp_lut_data : raw_reg33;
  assign _0337_ = _0384_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:1001" *) _3705_ : raw_reg33;
  assign _3706_ = _0483_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:992" *) reg2dp_lut_data : raw_reg32;
  assign _0336_ = _0384_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:991" *) _3706_ : raw_reg32;
  assign _3707_ = _0482_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:982" *) reg2dp_lut_data : raw_reg31;
  assign _0335_ = _0384_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:981" *) _3707_ : raw_reg31;
  assign _3708_ = _0481_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:972" *) reg2dp_lut_data : raw_reg30;
  assign _0334_ = _0384_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:971" *) _3708_ : raw_reg30;
  assign _3709_ = _0480_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:962" *) reg2dp_lut_data : raw_reg29;
  assign _0332_ = _0384_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:961" *) _3709_ : raw_reg29;
  assign _3710_ = _0479_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:952" *) reg2dp_lut_data : raw_reg28;
  assign _0331_ = _0384_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:951" *) _3710_ : raw_reg28;
  assign _3711_ = _0478_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:942" *) reg2dp_lut_data : raw_reg27;
  assign _0330_ = _0384_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:941" *) _3711_ : raw_reg27;
  assign _3712_ = _0477_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:932" *) reg2dp_lut_data : raw_reg26;
  assign _0329_ = _0384_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:931" *) _3712_ : raw_reg26;
  assign _3713_ = _0476_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:922" *) reg2dp_lut_data : raw_reg25;
  assign _0328_ = _0384_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:921" *) _3713_ : raw_reg25;
  assign _3714_ = _0475_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:912" *) reg2dp_lut_data : raw_reg24;
  assign _0327_ = _0384_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:911" *) _3714_ : raw_reg24;
  assign _3715_ = _0474_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:902" *) reg2dp_lut_data : raw_reg23;
  assign _0326_ = _0384_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:901" *) _3715_ : raw_reg23;
  assign _3716_ = _0473_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:892" *) reg2dp_lut_data : raw_reg22;
  assign _0325_ = _0384_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:891" *) _3716_ : raw_reg22;
  assign _3717_ = _0472_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:882" *) reg2dp_lut_data : raw_reg21;
  assign _0324_ = _0384_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:881" *) _3717_ : raw_reg21;
  assign _3718_ = _0471_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:872" *) reg2dp_lut_data : raw_reg20;
  assign _0323_ = _0384_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:871" *) _3718_ : raw_reg20;
  assign _3719_ = _0470_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:862" *) reg2dp_lut_data : raw_reg19;
  assign _0321_ = _0384_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:861" *) _3719_ : raw_reg19;
  assign _3720_ = _0469_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:852" *) reg2dp_lut_data : raw_reg18;
  assign _0320_ = _0384_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:851" *) _3720_ : raw_reg18;
  assign _3721_ = _0468_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:842" *) reg2dp_lut_data : raw_reg17;
  assign _0319_ = _0384_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:841" *) _3721_ : raw_reg17;
  assign _3722_ = _0467_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:832" *) reg2dp_lut_data : raw_reg16;
  assign _0318_ = _0384_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:831" *) _3722_ : raw_reg16;
  assign _3723_ = _0466_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:822" *) reg2dp_lut_data : raw_reg15;
  assign _0317_ = _0384_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:821" *) _3723_ : raw_reg15;
  assign _3724_ = _0465_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:812" *) reg2dp_lut_data : raw_reg14;
  assign _0316_ = _0384_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:811" *) _3724_ : raw_reg14;
  assign _3725_ = _0464_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:802" *) reg2dp_lut_data : raw_reg13;
  assign _0315_ = _0384_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:801" *) _3725_ : raw_reg13;
  assign _3726_ = _0463_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:792" *) reg2dp_lut_data : raw_reg12;
  assign _0314_ = _0384_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:791" *) _3726_ : raw_reg12;
  assign _3727_ = _0462_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:782" *) reg2dp_lut_data : raw_reg11;
  assign _0313_ = _0384_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:781" *) _3727_ : raw_reg11;
  assign _3728_ = _0461_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:772" *) reg2dp_lut_data : raw_reg10;
  assign _0312_ = _0384_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:771" *) _3728_ : raw_reg10;
  assign _3729_ = _0460_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:762" *) reg2dp_lut_data : raw_reg9;
  assign _0375_ = _0384_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:761" *) _3729_ : raw_reg9;
  assign _3730_ = _0459_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:752" *) reg2dp_lut_data : raw_reg8;
  assign _0374_ = _0384_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:751" *) _3730_ : raw_reg8;
  assign _3731_ = _0458_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:742" *) reg2dp_lut_data : raw_reg7;
  assign _0373_ = _0384_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:741" *) _3731_ : raw_reg7;
  assign _3732_ = _0457_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:732" *) reg2dp_lut_data : raw_reg6;
  assign _0372_ = _0384_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:731" *) _3732_ : raw_reg6;
  assign _3733_ = _0456_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:722" *) reg2dp_lut_data : raw_reg5;
  assign _0366_ = _0384_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:721" *) _3733_ : raw_reg5;
  assign _3734_ = _0455_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:712" *) reg2dp_lut_data : raw_reg4;
  assign _0355_ = _0384_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:711" *) _3734_ : raw_reg4;
  assign _3735_ = _0454_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:702" *) reg2dp_lut_data : raw_reg3;
  assign _0344_ = _0384_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:701" *) _3735_ : raw_reg3;
  assign _3736_ = _0453_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:692" *) reg2dp_lut_data : raw_reg2;
  assign _0333_ = _0384_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:691" *) _3736_ : raw_reg2;
  assign _3737_ = _0452_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:682" *) reg2dp_lut_data : raw_reg1;
  assign _0322_ = _0384_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:681" *) _3737_ : raw_reg1;
  assign _3738_ = _0451_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:672" *) reg2dp_lut_data : raw_reg0;
  assign _0311_ = _0384_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:671" *) _3738_ : raw_reg0;
  assign fp_lut_prdy_f = & (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:16761" *) { FMcvt_in_rdy[0], FMcvt_in_rdy[1], FMcvt_in_rdy[2], FMcvt_in_rdy[3] };
  assign _3739_ = & (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:16763" *) { FMcvt_in_rdy[1], FMcvt_in_rdy[2], FMcvt_in_rdy[3] };
  assign _3740_ = & (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:16764" *) { FMcvt_in_rdy[0], FMcvt_in_rdy[2], FMcvt_in_rdy[3] };
  assign _3741_ = & (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:16765" *) { FMcvt_in_rdy[0], FMcvt_in_rdy[1], FMcvt_in_rdy[3] };
  assign _3742_ = & (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:16766" *) { FMcvt_in_rdy[0], FMcvt_in_rdy[1], FMcvt_in_rdy[2] };
  assign _3743_ = & (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:16863" *) { FMcvt_out_vld[1], FMcvt_out_vld[2], FMcvt_out_vld[3] };
  assign _3744_ = & (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:16864" *) { FMcvt_out_vld[0], FMcvt_out_vld[2], FMcvt_out_vld[3] };
  assign _3745_ = & (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:16865" *) { FMcvt_out_vld[0], FMcvt_out_vld[1], FMcvt_out_vld[3] };
  assign _3746_ = & (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:16866" *) { FMcvt_out_vld[0], FMcvt_out_vld[1], FMcvt_out_vld[2] };
  assign fp_out_vld = & (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:16867" *) { FMcvt_out_vld[0], FMcvt_out_vld[1], FMcvt_out_vld[2], FMcvt_out_vld[3] };
  assign _3747_ = lutY_sel[0] ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:16716" *) lut_Y_data_00 : 16'b0000000000000000;
  assign lutX_data_00 = lutX_sel[0] ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:16716" *) lut_X_data_00 : _3747_;
  assign _3748_ = lutY_sel[0] ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:16717" *) lut_Y_data_01 : 16'b0000000000000000;
  assign lutX_data_01 = lutX_sel[0] ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:16717" *) lut_X_data_01 : _3748_;
  assign _3749_ = lutY_sel[0] ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:16718" *) lut_Y_info_0[15:0] : 16'b0000000000000000;
  assign lutX_info_0 = lutX_sel[0] ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:16718" *) lut_X_info_0[15:0] : _3749_;
  assign _3750_ = lutY_sel[1] ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:16719" *) lut_Y_data_10 : 16'b0000000000000000;
  assign lutX_data_10 = lutX_sel[1] ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:16719" *) lut_X_data_10 : _3750_;
  assign _3751_ = lutY_sel[1] ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:16720" *) lut_Y_data_11 : 16'b0000000000000000;
  assign lutX_data_11 = lutX_sel[1] ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:16720" *) lut_X_data_11 : _3751_;
  assign _3752_ = lutY_sel[1] ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:16721" *) lut_Y_info_1[15:0] : 16'b0000000000000000;
  assign lutX_info_1 = lutX_sel[1] ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:16721" *) lut_X_info_1[15:0] : _3752_;
  assign _3753_ = lutY_sel[2] ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:16722" *) lut_Y_data_20 : 16'b0000000000000000;
  assign lutX_data_20 = lutX_sel[2] ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:16722" *) lut_X_data_20 : _3753_;
  assign _3754_ = lutY_sel[2] ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:16723" *) lut_Y_data_21 : 16'b0000000000000000;
  assign lutX_data_21 = lutX_sel[2] ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:16723" *) lut_X_data_21 : _3754_;
  assign _3755_ = lutY_sel[2] ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:16724" *) lut_Y_info_2[15:0] : 16'b0000000000000000;
  assign lutX_info_2 = lutX_sel[2] ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:16724" *) lut_X_info_2[15:0] : _3755_;
  assign _3756_ = lutY_sel[3] ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:16725" *) lut_Y_data_30 : 16'b0000000000000000;
  assign lutX_data_30 = lutX_sel[3] ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:16725" *) lut_X_data_30 : _3756_;
  assign _3757_ = lutY_sel[3] ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:16726" *) lut_Y_data_31 : 16'b0000000000000000;
  assign lutX_data_31 = lutX_sel[3] ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:16726" *) lut_X_data_31 : _3757_;
  assign _3758_ = lutY_sel[3] ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:16727" *) lut_Y_info_3[15:0] : 16'b0000000000000000;
  assign lutX_info_3 = lutX_sel[3] ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:16727" *) lut_X_info_3[15:0] : _3758_;
  assign _3759_ = lutY_sel[4] ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:16728" *) lut_Y_data_40 : 16'b0000000000000000;
  assign lutX_data_40 = lutX_sel[4] ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:16728" *) lut_X_data_40 : _3759_;
  assign _3760_ = lutY_sel[4] ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:16729" *) lut_Y_data_41 : 16'b0000000000000000;
  assign lutX_data_41 = lutX_sel[4] ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:16729" *) lut_X_data_41 : _3760_;
  assign _3761_ = lutY_sel[4] ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:16730" *) lut_Y_info_4[15:0] : 16'b0000000000000000;
  assign lutX_info_4 = lutX_sel[4] ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:16730" *) lut_X_info_4[15:0] : _3761_;
  assign _3762_ = lutY_sel[5] ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:16731" *) lut_Y_data_50 : 16'b0000000000000000;
  assign lutX_data_50 = lutX_sel[5] ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:16731" *) lut_X_data_50 : _3762_;
  assign _3763_ = lutY_sel[5] ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:16732" *) lut_Y_data_51 : 16'b0000000000000000;
  assign lutX_data_51 = lutX_sel[5] ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:16732" *) lut_X_data_51 : _3763_;
  assign _3764_ = lutY_sel[5] ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:16733" *) lut_Y_info_5[15:0] : 16'b0000000000000000;
  assign lutX_info_5 = lutX_sel[5] ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:16733" *) lut_X_info_5[15:0] : _3764_;
  assign _3765_ = lutY_sel[6] ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:16734" *) lut_Y_data_60 : 16'b0000000000000000;
  assign lutX_data_60 = lutX_sel[6] ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:16734" *) lut_X_data_60 : _3765_;
  assign _3766_ = lutY_sel[6] ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:16735" *) lut_Y_data_61 : 16'b0000000000000000;
  assign lutX_data_61 = lutX_sel[6] ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:16735" *) lut_X_data_61 : _3766_;
  assign _3767_ = lutY_sel[6] ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:16736" *) lut_Y_info_6[15:0] : 16'b0000000000000000;
  assign lutX_info_6 = lutX_sel[6] ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:16736" *) lut_X_info_6[15:0] : _3767_;
  assign _3768_ = lutY_sel[7] ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:16737" *) lut_Y_data_70 : 16'b0000000000000000;
  assign lutX_data_70 = lutX_sel[7] ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:16737" *) lut_X_data_70 : _3768_;
  assign _3769_ = lutY_sel[7] ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:16738" *) lut_Y_data_71 : 16'b0000000000000000;
  assign lutX_data_71 = lutX_sel[7] ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:16738" *) lut_X_data_71 : _3769_;
  assign _3770_ = lutY_sel[7] ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:16739" *) lut_Y_info_7[15:0] : 16'b0000000000000000;
  assign lutX_info_7 = lutX_sel[7] ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:16739" *) lut_X_info_7[15:0] : _3770_;
  assign lut_prdy = fp16_en_f ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:16757" *) fp_lut_prdy_f : lut2intp_prdy;
  assign fp_lut_pvld_f = fp16_en_f ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:16762" *) lut_pvld_f : 1'b0;
  assign fp_out_prdy = fp16_en_f ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:16868" *) lut2intp_prdy : 1'b1;
  assign lut2intp_pvld = fp16_en_f ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:16872" *) fp_out_vld : lut_pvld_f;
  assign dp2reg_lut_data = reg2dp_lut_table_id ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:4553" *) density_out : raw_out;
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:16767" *)
  fp_format_cvt u_fp_format_cvt_0 (
    .FMcvt_in_rdy(FMcvt_in_rdy[0]),
    .FMcvt_in_vld(FMcvt_in_vld[0]),
    .FMcvt_out_rdy(FMcvt_out_rdy[0]),
    .FMcvt_out_vld(FMcvt_out_vld[0]),
    .fp16to17_in_X0(lutX_data_00),
    .fp16to17_out_X0(lut_X_dat_00_fp17),
    .fp16to32_in_X0(lutX_data_00),
    .fp16to32_in_X1(lutX_data_01),
    .fp16to32_out_X0(lut_X_dat_00),
    .fp16to32_out_X1(lut_X_dat_01),
    .lut_X_info_in(lut_X_info_0[17:16]),
    .lut_X_info_out(lut_X_inf_0[18:17]),
    .lut_X_sel_in(lutX_sel[0]),
    .lut_X_sel_out(lutX_sel_o[0]),
    .lut_Y_info_in(lut_Y_info_0[17:16]),
    .lut_Y_info_out(lut_X_inf_0[20:19]),
    .lut_Y_sel_in(lutY_sel[0]),
    .lut_Y_sel_out(lutY_sel_o[0]),
    .nvdla_core_clk(nvdla_op_gated_clk_fp16),
    .nvdla_core_rstn(nvdla_core_rstn),
    .uint16tofp17_Xin(lutX_info_0),
    .uint16tofp17_Xout(lut_X_inf_0[16:0])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:16791" *)
  fp_format_cvt u_fp_format_cvt_1 (
    .FMcvt_in_rdy(FMcvt_in_rdy[1]),
    .FMcvt_in_vld(FMcvt_in_vld[1]),
    .FMcvt_out_rdy(FMcvt_out_rdy[1]),
    .FMcvt_out_vld(FMcvt_out_vld[1]),
    .fp16to17_in_X0(lutX_data_10),
    .fp16to17_out_X0(lut_X_dat_10_fp17),
    .fp16to32_in_X0(lutX_data_10),
    .fp16to32_in_X1(lutX_data_11),
    .fp16to32_out_X0(lut_X_dat_10),
    .fp16to32_out_X1(lut_X_dat_11),
    .lut_X_info_in(lut_X_info_1[17:16]),
    .lut_X_info_out(lut_X_inf_1[18:17]),
    .lut_X_sel_in(lutX_sel[1]),
    .lut_X_sel_out(lutX_sel_o[1]),
    .lut_Y_info_in(lut_Y_info_1[17:16]),
    .lut_Y_info_out(lut_X_inf_1[20:19]),
    .lut_Y_sel_in(lutY_sel[1]),
    .lut_Y_sel_out(lutY_sel_o[1]),
    .nvdla_core_clk(nvdla_op_gated_clk_fp16),
    .nvdla_core_rstn(nvdla_core_rstn),
    .uint16tofp17_Xin(lutX_info_1),
    .uint16tofp17_Xout(lut_X_inf_1[16:0])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:16815" *)
  fp_format_cvt u_fp_format_cvt_2 (
    .FMcvt_in_rdy(FMcvt_in_rdy[2]),
    .FMcvt_in_vld(FMcvt_in_vld[2]),
    .FMcvt_out_rdy(FMcvt_out_rdy[2]),
    .FMcvt_out_vld(FMcvt_out_vld[2]),
    .fp16to17_in_X0(lutX_data_20),
    .fp16to17_out_X0(lut_X_dat_20_fp17),
    .fp16to32_in_X0(lutX_data_20),
    .fp16to32_in_X1(lutX_data_21),
    .fp16to32_out_X0(lut_X_dat_20),
    .fp16to32_out_X1(lut_X_dat_21),
    .lut_X_info_in(lut_X_info_2[17:16]),
    .lut_X_info_out(lut_X_inf_2[18:17]),
    .lut_X_sel_in(lutX_sel[2]),
    .lut_X_sel_out(lutX_sel_o[2]),
    .lut_Y_info_in(lut_Y_info_2[17:16]),
    .lut_Y_info_out(lut_X_inf_2[20:19]),
    .lut_Y_sel_in(lutY_sel[2]),
    .lut_Y_sel_out(lutY_sel_o[2]),
    .nvdla_core_clk(nvdla_op_gated_clk_fp16),
    .nvdla_core_rstn(nvdla_core_rstn),
    .uint16tofp17_Xin(lutX_info_2),
    .uint16tofp17_Xout(lut_X_inf_2[16:0])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_DP_lut.v:16839" *)
  fp_format_cvt u_fp_format_cvt_3 (
    .FMcvt_in_rdy(FMcvt_in_rdy[3]),
    .FMcvt_in_vld(FMcvt_in_vld[3]),
    .FMcvt_out_rdy(FMcvt_out_rdy[3]),
    .FMcvt_out_vld(FMcvt_out_vld[3]),
    .fp16to17_in_X0(lutX_data_30),
    .fp16to17_out_X0(lut_X_dat_30_fp17),
    .fp16to32_in_X0(lutX_data_30),
    .fp16to32_in_X1(lutX_data_31),
    .fp16to32_out_X0(lut_X_dat_30),
    .fp16to32_out_X1(lut_X_dat_31),
    .lut_X_info_in(lut_X_info_3[17:16]),
    .lut_X_info_out(lut_X_inf_3[18:17]),
    .lut_X_sel_in(lutX_sel[3]),
    .lut_X_sel_out(lutX_sel_o[3]),
    .lut_Y_info_in(lut_Y_info_3[17:16]),
    .lut_Y_info_out(lut_X_inf_3[20:19]),
    .lut_Y_sel_in(lutY_sel[3]),
    .lut_Y_sel_out(lutY_sel_o[3]),
    .nvdla_core_clk(nvdla_op_gated_clk_fp16),
    .nvdla_core_rstn(nvdla_core_rstn),
    .uint16tofp17_Xin(lutX_info_3),
    .uint16tofp17_Xout(lut_X_inf_3[16:0])
  );
  assign both_hybrid_sel = reg2dp_lut_hybrid_priority;
  assign both_of_sel = reg2dp_lut_oflow_priority;
  assign both_uf_sel = reg2dp_lut_uflow_priority;
  assign dp2lut_prdy = dp2lut_prdy_f;
endmodule
