module S(clk, in, out);
  wire [7:0] _000_;
  wire _001_;
  wire _002_;
  wire _003_;
  wire _004_;
  wire _005_;
  wire _006_;
  wire _007_;
  wire _008_;
  wire _009_;
  wire _010_;
  wire _011_;
  wire _012_;
  wire _013_;
  wire _014_;
  wire _015_;
  wire _016_;
  wire _017_;
  wire _018_;
  wire _019_;
  wire _020_;
  wire _021_;
  wire _022_;
  wire _023_;
  wire _024_;
  wire _025_;
  wire _026_;
  wire _027_;
  wire _028_;
  wire _029_;
  wire _030_;
  wire _031_;
  wire _032_;
  wire _033_;
  wire _034_;
  wire _035_;
  wire _036_;
  wire _037_;
  wire _038_;
  wire _039_;
  wire _040_;
  wire _041_;
  wire _042_;
  wire _043_;
  wire _044_;
  wire _045_;
  wire _046_;
  wire _047_;
  wire _048_;
  wire _049_;
  wire _050_;
  wire _051_;
  wire _052_;
  wire _053_;
  wire _054_;
  wire _055_;
  wire _056_;
  wire _057_;
  wire _058_;
  wire _059_;
  wire _060_;
  wire _061_;
  wire _062_;
  wire _063_;
  wire _064_;
  wire _065_;
  wire _066_;
  wire _067_;
  wire _068_;
  wire _069_;
  wire _070_;
  wire _071_;
  wire _072_;
  wire _073_;
  wire _074_;
  wire _075_;
  wire _076_;
  wire _077_;
  wire _078_;
  wire _079_;
  wire _080_;
  wire _081_;
  wire _082_;
  wire _083_;
  wire _084_;
  wire _085_;
  wire _086_;
  wire _087_;
  wire _088_;
  wire _089_;
  wire _090_;
  wire _091_;
  wire _092_;
  wire _093_;
  wire _094_;
  wire _095_;
  wire _096_;
  wire _097_;
  wire _098_;
  wire _099_;
  wire _100_;
  wire _101_;
  wire _102_;
  wire _103_;
  wire _104_;
  wire _105_;
  wire _106_;
  wire _107_;
  wire _108_;
  wire _109_;
  wire _110_;
  wire _111_;
  wire _112_;
  wire _113_;
  wire _114_;
  wire _115_;
  wire _116_;
  wire _117_;
  wire _118_;
  wire _119_;
  wire _120_;
  wire _121_;
  wire _122_;
  wire _123_;
  wire _124_;
  wire _125_;
  wire _126_;
  wire _127_;
  wire _128_;
  wire _129_;
  wire _130_;
  wire _131_;
  wire _132_;
  wire _133_;
  wire _134_;
  wire _135_;
  wire _136_;
  wire _137_;
  wire _138_;
  wire _139_;
  wire _140_;
  wire _141_;
  wire _142_;
  wire _143_;
  wire _144_;
  wire _145_;
  wire _146_;
  wire _147_;
  wire _148_;
  wire _149_;
  wire _150_;
  wire _151_;
  wire _152_;
  wire _153_;
  wire _154_;
  wire _155_;
  wire _156_;
  wire _157_;
  wire _158_;
  wire _159_;
  wire _160_;
  wire _161_;
  wire _162_;
  wire _163_;
  wire _164_;
  wire _165_;
  wire _166_;
  wire _167_;
  wire _168_;
  wire _169_;
  wire _170_;
  wire _171_;
  wire _172_;
  wire _173_;
  wire _174_;
  wire _175_;
  wire _176_;
  wire _177_;
  wire _178_;
  wire _179_;
  wire _180_;
  wire _181_;
  wire _182_;
  wire _183_;
  wire _184_;
  wire _185_;
  wire _186_;
  wire _187_;
  wire _188_;
  wire _189_;
  wire _190_;
  wire _191_;
  wire _192_;
  wire _193_;
  wire _194_;
  wire _195_;
  wire _196_;
  wire _197_;
  wire _198_;
  wire _199_;
  wire _200_;
  wire _201_;
  wire _202_;
  wire _203_;
  wire _204_;
  wire _205_;
  wire _206_;
  wire _207_;
  wire _208_;
  wire _209_;
  wire _210_;
  wire _211_;
  wire _212_;
  wire _213_;
  wire _214_;
  wire _215_;
  wire _216_;
  wire _217_;
  wire _218_;
  wire _219_;
  wire _220_;
  wire _221_;
  wire _222_;
  wire _223_;
  wire _224_;
  wire _225_;
  wire _226_;
  wire _227_;
  wire _228_;
  wire _229_;
  wire _230_;
  wire _231_;
  wire _232_;
  wire _233_;
  wire _234_;
  wire _235_;
  wire _236_;
  wire _237_;
  wire _238_;
  wire _239_;
  wire _240_;
  wire _241_;
  wire _242_;
  wire _243_;
  wire _244_;
  wire _245_;
  wire _246_;
  wire _247_;
  wire _248_;
  wire _249_;
  wire _250_;
  wire _251_;
  wire _252_;
  wire _253_;
  wire _254_;
  wire _255_;
  input clk;
  input [7:0] in;
  output [7:0] out;
  reg [7:0] out;
  always @(posedge clk)
    out <= _000_;
  function [7:0] _257_;
    input [7:0] a;
    input [2039:0] b;
    input [254:0] s;
    casez (s) // synopsys parallel_case
      255'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1:
        _257_ = b[7:0];
      255'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?:
        _257_ = b[15:8];
      255'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??:
        _257_ = b[23:16];
      255'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???:
        _257_ = b[31:24];
      255'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????:
        _257_ = b[39:32];
      255'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????:
        _257_ = b[47:40];
      255'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????:
        _257_ = b[55:48];
      255'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????:
        _257_ = b[63:56];
      255'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????:
        _257_ = b[71:64];
      255'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????:
        _257_ = b[79:72];
      255'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????:
        _257_ = b[87:80];
      255'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????:
        _257_ = b[95:88];
      255'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????:
        _257_ = b[103:96];
      255'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????:
        _257_ = b[111:104];
      255'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????:
        _257_ = b[119:112];
      255'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????:
        _257_ = b[127:120];
      255'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????:
        _257_ = b[135:128];
      255'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????:
        _257_ = b[143:136];
      255'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????:
        _257_ = b[151:144];
      255'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????:
        _257_ = b[159:152];
      255'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????:
        _257_ = b[167:160];
      255'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????:
        _257_ = b[175:168];
      255'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????:
        _257_ = b[183:176];
      255'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????:
        _257_ = b[191:184];
      255'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????:
        _257_ = b[199:192];
      255'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????:
        _257_ = b[207:200];
      255'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????:
        _257_ = b[215:208];
      255'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????:
        _257_ = b[223:216];
      255'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????:
        _257_ = b[231:224];
      255'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????:
        _257_ = b[239:232];
      255'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????:
        _257_ = b[247:240];
      255'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????:
        _257_ = b[255:248];
      255'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????:
        _257_ = b[263:256];
      255'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????:
        _257_ = b[271:264];
      255'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????:
        _257_ = b[279:272];
      255'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????:
        _257_ = b[287:280];
      255'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????:
        _257_ = b[295:288];
      255'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????:
        _257_ = b[303:296];
      255'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????:
        _257_ = b[311:304];
      255'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????:
        _257_ = b[319:312];
      255'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????:
        _257_ = b[327:320];
      255'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????:
        _257_ = b[335:328];
      255'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????:
        _257_ = b[343:336];
      255'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????:
        _257_ = b[351:344];
      255'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????:
        _257_ = b[359:352];
      255'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????:
        _257_ = b[367:360];
      255'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????:
        _257_ = b[375:368];
      255'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????:
        _257_ = b[383:376];
      255'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????:
        _257_ = b[391:384];
      255'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????:
        _257_ = b[399:392];
      255'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????:
        _257_ = b[407:400];
      255'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????:
        _257_ = b[415:408];
      255'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????:
        _257_ = b[423:416];
      255'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????:
        _257_ = b[431:424];
      255'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????:
        _257_ = b[439:432];
      255'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????:
        _257_ = b[447:440];
      255'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????:
        _257_ = b[455:448];
      255'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????:
        _257_ = b[463:456];
      255'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????:
        _257_ = b[471:464];
      255'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????:
        _257_ = b[479:472];
      255'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????:
        _257_ = b[487:480];
      255'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????:
        _257_ = b[495:488];
      255'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????:
        _257_ = b[503:496];
      255'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????:
        _257_ = b[511:504];
      255'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????:
        _257_ = b[519:512];
      255'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????:
        _257_ = b[527:520];
      255'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????:
        _257_ = b[535:528];
      255'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????:
        _257_ = b[543:536];
      255'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????:
        _257_ = b[551:544];
      255'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????:
        _257_ = b[559:552];
      255'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????:
        _257_ = b[567:560];
      255'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????:
        _257_ = b[575:568];
      255'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????:
        _257_ = b[583:576];
      255'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????:
        _257_ = b[591:584];
      255'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????:
        _257_ = b[599:592];
      255'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????:
        _257_ = b[607:600];
      255'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????:
        _257_ = b[615:608];
      255'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????:
        _257_ = b[623:616];
      255'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????:
        _257_ = b[631:624];
      255'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????:
        _257_ = b[639:632];
      255'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????:
        _257_ = b[647:640];
      255'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????:
        _257_ = b[655:648];
      255'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????:
        _257_ = b[663:656];
      255'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????:
        _257_ = b[671:664];
      255'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????:
        _257_ = b[679:672];
      255'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????:
        _257_ = b[687:680];
      255'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????:
        _257_ = b[695:688];
      255'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????:
        _257_ = b[703:696];
      255'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????:
        _257_ = b[711:704];
      255'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????:
        _257_ = b[719:712];
      255'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????:
        _257_ = b[727:720];
      255'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????:
        _257_ = b[735:728];
      255'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????:
        _257_ = b[743:736];
      255'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????:
        _257_ = b[751:744];
      255'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????:
        _257_ = b[759:752];
      255'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????:
        _257_ = b[767:760];
      255'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????:
        _257_ = b[775:768];
      255'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????:
        _257_ = b[783:776];
      255'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????:
        _257_ = b[791:784];
      255'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????:
        _257_ = b[799:792];
      255'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????:
        _257_ = b[807:800];
      255'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????:
        _257_ = b[815:808];
      255'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????:
        _257_ = b[823:816];
      255'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????:
        _257_ = b[831:824];
      255'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _257_ = b[839:832];
      255'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _257_ = b[847:840];
      255'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _257_ = b[855:848];
      255'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _257_ = b[863:856];
      255'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _257_ = b[871:864];
      255'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _257_ = b[879:872];
      255'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _257_ = b[887:880];
      255'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _257_ = b[895:888];
      255'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _257_ = b[903:896];
      255'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _257_ = b[911:904];
      255'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _257_ = b[919:912];
      255'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _257_ = b[927:920];
      255'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _257_ = b[935:928];
      255'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _257_ = b[943:936];
      255'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _257_ = b[951:944];
      255'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _257_ = b[959:952];
      255'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _257_ = b[967:960];
      255'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _257_ = b[975:968];
      255'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _257_ = b[983:976];
      255'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _257_ = b[991:984];
      255'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _257_ = b[999:992];
      255'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _257_ = b[1007:1000];
      255'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _257_ = b[1015:1008];
      255'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _257_ = b[1023:1016];
      255'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _257_ = b[1031:1024];
      255'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _257_ = b[1039:1032];
      255'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _257_ = b[1047:1040];
      255'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _257_ = b[1055:1048];
      255'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _257_ = b[1063:1056];
      255'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _257_ = b[1071:1064];
      255'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _257_ = b[1079:1072];
      255'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _257_ = b[1087:1080];
      255'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _257_ = b[1095:1088];
      255'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _257_ = b[1103:1096];
      255'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _257_ = b[1111:1104];
      255'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _257_ = b[1119:1112];
      255'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _257_ = b[1127:1120];
      255'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _257_ = b[1135:1128];
      255'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _257_ = b[1143:1136];
      255'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _257_ = b[1151:1144];
      255'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _257_ = b[1159:1152];
      255'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _257_ = b[1167:1160];
      255'b????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _257_ = b[1175:1168];
      255'b???????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _257_ = b[1183:1176];
      255'b??????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _257_ = b[1191:1184];
      255'b?????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _257_ = b[1199:1192];
      255'b????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _257_ = b[1207:1200];
      255'b???????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _257_ = b[1215:1208];
      255'b??????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _257_ = b[1223:1216];
      255'b?????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _257_ = b[1231:1224];
      255'b????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _257_ = b[1239:1232];
      255'b???????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _257_ = b[1247:1240];
      255'b??????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _257_ = b[1255:1248];
      255'b?????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _257_ = b[1263:1256];
      255'b????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _257_ = b[1271:1264];
      255'b???????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _257_ = b[1279:1272];
      255'b??????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _257_ = b[1287:1280];
      255'b?????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _257_ = b[1295:1288];
      255'b????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _257_ = b[1303:1296];
      255'b???????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _257_ = b[1311:1304];
      255'b??????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _257_ = b[1319:1312];
      255'b?????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _257_ = b[1327:1320];
      255'b????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _257_ = b[1335:1328];
      255'b???????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _257_ = b[1343:1336];
      255'b??????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _257_ = b[1351:1344];
      255'b?????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _257_ = b[1359:1352];
      255'b????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _257_ = b[1367:1360];
      255'b???????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _257_ = b[1375:1368];
      255'b??????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _257_ = b[1383:1376];
      255'b?????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _257_ = b[1391:1384];
      255'b????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _257_ = b[1399:1392];
      255'b???????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _257_ = b[1407:1400];
      255'b??????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _257_ = b[1415:1408];
      255'b?????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _257_ = b[1423:1416];
      255'b????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _257_ = b[1431:1424];
      255'b???????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _257_ = b[1439:1432];
      255'b??????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _257_ = b[1447:1440];
      255'b?????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _257_ = b[1455:1448];
      255'b????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _257_ = b[1463:1456];
      255'b???????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _257_ = b[1471:1464];
      255'b??????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _257_ = b[1479:1472];
      255'b?????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _257_ = b[1487:1480];
      255'b????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _257_ = b[1495:1488];
      255'b???????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _257_ = b[1503:1496];
      255'b??????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _257_ = b[1511:1504];
      255'b?????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _257_ = b[1519:1512];
      255'b????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _257_ = b[1527:1520];
      255'b???????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _257_ = b[1535:1528];
      255'b??????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _257_ = b[1543:1536];
      255'b?????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _257_ = b[1551:1544];
      255'b????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _257_ = b[1559:1552];
      255'b???????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _257_ = b[1567:1560];
      255'b??????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _257_ = b[1575:1568];
      255'b?????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _257_ = b[1583:1576];
      255'b????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _257_ = b[1591:1584];
      255'b???????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _257_ = b[1599:1592];
      255'b??????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _257_ = b[1607:1600];
      255'b?????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _257_ = b[1615:1608];
      255'b????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _257_ = b[1623:1616];
      255'b???????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _257_ = b[1631:1624];
      255'b??????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _257_ = b[1639:1632];
      255'b?????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _257_ = b[1647:1640];
      255'b????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _257_ = b[1655:1648];
      255'b???????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _257_ = b[1663:1656];
      255'b??????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _257_ = b[1671:1664];
      255'b?????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _257_ = b[1679:1672];
      255'b????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _257_ = b[1687:1680];
      255'b???????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _257_ = b[1695:1688];
      255'b??????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _257_ = b[1703:1696];
      255'b?????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _257_ = b[1711:1704];
      255'b????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _257_ = b[1719:1712];
      255'b???????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _257_ = b[1727:1720];
      255'b??????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _257_ = b[1735:1728];
      255'b?????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _257_ = b[1743:1736];
      255'b????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _257_ = b[1751:1744];
      255'b???????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _257_ = b[1759:1752];
      255'b??????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _257_ = b[1767:1760];
      255'b?????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _257_ = b[1775:1768];
      255'b????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _257_ = b[1783:1776];
      255'b???????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _257_ = b[1791:1784];
      255'b??????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _257_ = b[1799:1792];
      255'b?????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _257_ = b[1807:1800];
      255'b????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _257_ = b[1815:1808];
      255'b???????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _257_ = b[1823:1816];
      255'b??????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _257_ = b[1831:1824];
      255'b?????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _257_ = b[1839:1832];
      255'b????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _257_ = b[1847:1840];
      255'b???????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _257_ = b[1855:1848];
      255'b??????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _257_ = b[1863:1856];
      255'b?????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _257_ = b[1871:1864];
      255'b????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _257_ = b[1879:1872];
      255'b???????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _257_ = b[1887:1880];
      255'b??????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _257_ = b[1895:1888];
      255'b?????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _257_ = b[1903:1896];
      255'b????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _257_ = b[1911:1904];
      255'b???????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _257_ = b[1919:1912];
      255'b??????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _257_ = b[1927:1920];
      255'b?????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _257_ = b[1935:1928];
      255'b????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _257_ = b[1943:1936];
      255'b???????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _257_ = b[1951:1944];
      255'b??????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _257_ = b[1959:1952];
      255'b?????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _257_ = b[1967:1960];
      255'b????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _257_ = b[1975:1968];
      255'b???????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _257_ = b[1983:1976];
      255'b??????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _257_ = b[1991:1984];
      255'b?????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _257_ = b[1999:1992];
      255'b????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _257_ = b[2007:2000];
      255'b???1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _257_ = b[2015:2008];
      255'b??1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _257_ = b[2023:2016];
      255'b?1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _257_ = b[2031:2024];
      255'b1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _257_ = b[2039:2032];
      default:
        _257_ = a;
    endcase
  endfunction
  assign _000_ = _257_(8'b01100011, 2040'b011111000111011101111011111100100110101101101111110001010011000000000001011001110010101111111110110101111010101101110110110010101000001011001001011111011111101001011001010001111111000010101101110101001010001010101111100111001010010001110010110000001011011111111101100100110010011000110110001111111111011111001100001101001010010111100101111100010111000111011000001100010001010100000100110001110010001111000011000110001001011000000101100110100000011100010010100000001110001011101011001001111011001001110101000010011000001100101100000110100001101101101110010110101010000001010010001110111101011010110011001010011110001100101111100001000101001111010001000000001110110100100000111111001011000101011011011010101100101110111110001110010100101001001100010110001100111111010000111011111010101011111011010000110100110100110011100001010100010111111001000000100111111101010000001111001001111110101000010100011010001101000000100011111001001010011101001110001111010110111100101101101101101000100001000100001111111111110011110100101100110100001100000100111110110001011111100101110100010000010111110001001010011101111110001111010110010001011101000110010111001101100000100000010100111111011100001000100010101010010000100010000100011011101110101110000001010011011110010111100000101111011011111000000011001000111010000010100100100100000110001001000101110011000010110100111010110001100010100100011001010111100100011110011110011111001000001101110110110110001101110101010100111010101001011011000101011011110100111010100110010101111010101011100000100010111010011110000010010100101110000111001010011010110100110001101110100011011101011101000001111101001011101111011000101110001010011100000011111010110101011001100100100000000011111101100000111001100001001101010101011110111001100001101100000100011101100111101110000111111000100110000001000101101001110110011000111010010100100110110001111010000111111010011100111001010101001010001101111110001100101000011000100100001101101111111110011001000010011010000100000110011001001011010000111110110000010101001011101100010110, { _255_, _254_, _253_, _252_, _251_, _250_, _249_, _248_, _247_, _246_, _245_, _244_, _243_, _242_, _241_, _240_, _239_, _238_, _237_, _236_, _235_, _234_, _233_, _232_, _231_, _230_, _229_, _228_, _227_, _226_, _225_, _224_, _223_, _222_, _221_, _220_, _219_, _218_, _217_, _216_, _215_, _214_, _213_, _212_, _211_, _210_, _209_, _208_, _207_, _206_, _205_, _204_, _203_, _202_, _201_, _200_, _199_, _198_, _197_, _196_, _195_, _194_, _193_, _192_, _191_, _190_, _189_, _188_, _187_, _186_, _185_, _184_, _183_, _182_, _181_, _180_, _179_, _178_, _177_, _176_, _175_, _174_, _173_, _172_, _171_, _170_, _169_, _168_, _167_, _166_, _165_, _164_, _163_, _162_, _161_, _160_, _159_, _158_, _157_, _156_, _155_, _154_, _153_, _152_, _151_, _150_, _149_, _148_, _147_, _146_, _145_, _144_, _143_, _142_, _141_, _140_, _139_, _138_, _137_, _136_, _135_, _134_, _133_, _132_, _131_, _130_, _129_, _128_, _127_, _126_, _125_, _124_, _123_, _122_, _121_, _120_, _119_, _118_, _117_, _116_, _115_, _114_, _113_, _112_, _111_, _110_, _109_, _108_, _107_, _106_, _105_, _104_, _103_, _102_, _101_, _100_, _099_, _098_, _097_, _096_, _095_, _094_, _093_, _092_, _091_, _090_, _089_, _088_, _087_, _086_, _085_, _084_, _083_, _082_, _081_, _080_, _079_, _078_, _077_, _076_, _075_, _074_, _073_, _072_, _071_, _070_, _069_, _068_, _067_, _066_, _065_, _064_, _063_, _062_, _061_, _060_, _059_, _058_, _057_, _056_, _055_, _054_, _053_, _052_, _051_, _050_, _049_, _048_, _047_, _046_, _045_, _044_, _043_, _042_, _041_, _040_, _039_, _038_, _037_, _036_, _035_, _034_, _033_, _032_, _031_, _030_, _029_, _028_, _027_, _026_, _025_, _024_, _023_, _022_, _021_, _020_, _019_, _018_, _017_, _016_, _015_, _014_, _013_, _012_, _011_, _010_, _009_, _008_, _007_, _006_, _005_, _004_, _003_, _002_, _001_ });
  assign _001_ = in == 8'b11111111;
  assign _002_ = in == 8'b11111110;
  assign _003_ = in == 8'b11111101;
  assign _004_ = in == 8'b11111100;
  assign _005_ = in == 8'b11111011;
  assign _006_ = in == 8'b11111010;
  assign _007_ = in == 8'b11111001;
  assign _008_ = in == 8'b11111000;
  assign _009_ = in == 8'b11110111;
  assign _010_ = in == 8'b11110110;
  assign _011_ = in == 8'b11110101;
  assign _012_ = in == 8'b11110100;
  assign _013_ = in == 8'b11110011;
  assign _014_ = in == 8'b11110010;
  assign _015_ = in == 8'b11110001;
  assign _016_ = in == 8'b11110000;
  assign _017_ = in == 8'b11101111;
  assign _018_ = in == 8'b11101110;
  assign _019_ = in == 8'b11101101;
  assign _020_ = in == 8'b11101100;
  assign _021_ = in == 8'b11101011;
  assign _022_ = in == 8'b11101010;
  assign _023_ = in == 8'b11101001;
  assign _024_ = in == 8'b11101000;
  assign _025_ = in == 8'b11100111;
  assign _026_ = in == 8'b11100110;
  assign _027_ = in == 8'b11100101;
  assign _028_ = in == 8'b11100100;
  assign _029_ = in == 8'b11100011;
  assign _030_ = in == 8'b11100010;
  assign _031_ = in == 8'b11100001;
  assign _032_ = in == 8'b11100000;
  assign _033_ = in == 8'b11011111;
  assign _034_ = in == 8'b11011110;
  assign _035_ = in == 8'b11011101;
  assign _036_ = in == 8'b11011100;
  assign _037_ = in == 8'b11011011;
  assign _038_ = in == 8'b11011010;
  assign _039_ = in == 8'b11011001;
  assign _040_ = in == 8'b11011000;
  assign _041_ = in == 8'b11010111;
  assign _042_ = in == 8'b11010110;
  assign _043_ = in == 8'b11010101;
  assign _044_ = in == 8'b11010100;
  assign _045_ = in == 8'b11010011;
  assign _046_ = in == 8'b11010010;
  assign _047_ = in == 8'b11010001;
  assign _048_ = in == 8'b11010000;
  assign _049_ = in == 8'b11001111;
  assign _050_ = in == 8'b11001110;
  assign _051_ = in == 8'b11001101;
  assign _052_ = in == 8'b11001100;
  assign _053_ = in == 8'b11001011;
  assign _054_ = in == 8'b11001010;
  assign _055_ = in == 8'b11001001;
  assign _056_ = in == 8'b11001000;
  assign _057_ = in == 8'b11000111;
  assign _058_ = in == 8'b11000110;
  assign _059_ = in == 8'b11000101;
  assign _060_ = in == 8'b11000100;
  assign _061_ = in == 8'b11000011;
  assign _062_ = in == 8'b11000010;
  assign _063_ = in == 8'b11000001;
  assign _064_ = in == 8'b11000000;
  assign _065_ = in == 8'b10111111;
  assign _066_ = in == 8'b10111110;
  assign _067_ = in == 8'b10111101;
  assign _068_ = in == 8'b10111100;
  assign _069_ = in == 8'b10111011;
  assign _070_ = in == 8'b10111010;
  assign _071_ = in == 8'b10111001;
  assign _072_ = in == 8'b10111000;
  assign _073_ = in == 8'b10110111;
  assign _074_ = in == 8'b10110110;
  assign _075_ = in == 8'b10110101;
  assign _076_ = in == 8'b10110100;
  assign _077_ = in == 8'b10110011;
  assign _078_ = in == 8'b10110010;
  assign _079_ = in == 8'b10110001;
  assign _080_ = in == 8'b10110000;
  assign _081_ = in == 8'b10101111;
  assign _082_ = in == 8'b10101110;
  assign _083_ = in == 8'b10101101;
  assign _084_ = in == 8'b10101100;
  assign _085_ = in == 8'b10101011;
  assign _086_ = in == 8'b10101010;
  assign _087_ = in == 8'b10101001;
  assign _088_ = in == 8'b10101000;
  assign _089_ = in == 8'b10100111;
  assign _090_ = in == 8'b10100110;
  assign _091_ = in == 8'b10100101;
  assign _092_ = in == 8'b10100100;
  assign _093_ = in == 8'b10100011;
  assign _094_ = in == 8'b10100010;
  assign _095_ = in == 8'b10100001;
  assign _096_ = in == 8'b10100000;
  assign _097_ = in == 8'b10011111;
  assign _098_ = in == 8'b10011110;
  assign _099_ = in == 8'b10011101;
  assign _100_ = in == 8'b10011100;
  assign _101_ = in == 8'b10011011;
  assign _102_ = in == 8'b10011010;
  assign _103_ = in == 8'b10011001;
  assign _104_ = in == 8'b10011000;
  assign _105_ = in == 8'b10010111;
  assign _106_ = in == 8'b10010110;
  assign _107_ = in == 8'b10010101;
  assign _108_ = in == 8'b10010100;
  assign _109_ = in == 8'b10010011;
  assign _110_ = in == 8'b10010010;
  assign _111_ = in == 8'b10010001;
  assign _112_ = in == 8'b10010000;
  assign _113_ = in == 8'b10001111;
  assign _114_ = in == 8'b10001110;
  assign _115_ = in == 8'b10001101;
  assign _116_ = in == 8'b10001100;
  assign _117_ = in == 8'b10001011;
  assign _118_ = in == 8'b10001010;
  assign _119_ = in == 8'b10001001;
  assign _120_ = in == 8'b10001000;
  assign _121_ = in == 8'b10000111;
  assign _122_ = in == 8'b10000110;
  assign _123_ = in == 8'b10000101;
  assign _124_ = in == 8'b10000100;
  assign _125_ = in == 8'b10000011;
  assign _126_ = in == 8'b10000010;
  assign _127_ = in == 8'b10000001;
  assign _128_ = in == 8'b10000000;
  assign _129_ = in == 7'b1111111;
  assign _130_ = in == 7'b1111110;
  assign _131_ = in == 7'b1111101;
  assign _132_ = in == 7'b1111100;
  assign _133_ = in == 7'b1111011;
  assign _134_ = in == 7'b1111010;
  assign _135_ = in == 7'b1111001;
  assign _136_ = in == 7'b1111000;
  assign _137_ = in == 7'b1110111;
  assign _138_ = in == 7'b1110110;
  assign _139_ = in == 7'b1110101;
  assign _140_ = in == 7'b1110100;
  assign _141_ = in == 7'b1110011;
  assign _142_ = in == 7'b1110010;
  assign _143_ = in == 7'b1110001;
  assign _144_ = in == 7'b1110000;
  assign _145_ = in == 7'b1101111;
  assign _146_ = in == 7'b1101110;
  assign _147_ = in == 7'b1101101;
  assign _148_ = in == 7'b1101100;
  assign _149_ = in == 7'b1101011;
  assign _150_ = in == 7'b1101010;
  assign _151_ = in == 7'b1101001;
  assign _152_ = in == 7'b1101000;
  assign _153_ = in == 7'b1100111;
  assign _154_ = in == 7'b1100110;
  assign _155_ = in == 7'b1100101;
  assign _156_ = in == 7'b1100100;
  assign _157_ = in == 7'b1100011;
  assign _158_ = in == 7'b1100010;
  assign _159_ = in == 7'b1100001;
  assign _160_ = in == 7'b1100000;
  assign _161_ = in == 7'b1011111;
  assign _162_ = in == 7'b1011110;
  assign _163_ = in == 7'b1011101;
  assign _164_ = in == 7'b1011100;
  assign _165_ = in == 7'b1011011;
  assign _166_ = in == 7'b1011010;
  assign _167_ = in == 7'b1011001;
  assign _168_ = in == 7'b1011000;
  assign _169_ = in == 7'b1010111;
  assign _170_ = in == 7'b1010110;
  assign _171_ = in == 7'b1010101;
  assign _172_ = in == 7'b1010100;
  assign _173_ = in == 7'b1010011;
  assign _174_ = in == 7'b1010010;
  assign _175_ = in == 7'b1010001;
  assign _176_ = in == 7'b1010000;
  assign _177_ = in == 7'b1001111;
  assign _178_ = in == 7'b1001110;
  assign _179_ = in == 7'b1001101;
  assign _180_ = in == 7'b1001100;
  assign _181_ = in == 7'b1001011;
  assign _182_ = in == 7'b1001010;
  assign _183_ = in == 7'b1001001;
  assign _184_ = in == 7'b1001000;
  assign _185_ = in == 7'b1000111;
  assign _186_ = in == 7'b1000110;
  assign _187_ = in == 7'b1000101;
  assign _188_ = in == 7'b1000100;
  assign _189_ = in == 7'b1000011;
  assign _190_ = in == 7'b1000010;
  assign _191_ = in == 7'b1000001;
  assign _192_ = in == 7'b1000000;
  assign _193_ = in == 6'b111111;
  assign _194_ = in == 6'b111110;
  assign _195_ = in == 6'b111101;
  assign _196_ = in == 6'b111100;
  assign _197_ = in == 6'b111011;
  assign _198_ = in == 6'b111010;
  assign _199_ = in == 6'b111001;
  assign _200_ = in == 6'b111000;
  assign _201_ = in == 6'b110111;
  assign _202_ = in == 6'b110110;
  assign _203_ = in == 6'b110101;
  assign _204_ = in == 6'b110100;
  assign _205_ = in == 6'b110011;
  assign _206_ = in == 6'b110010;
  assign _207_ = in == 6'b110001;
  assign _208_ = in == 6'b110000;
  assign _209_ = in == 6'b101111;
  assign _210_ = in == 6'b101110;
  assign _211_ = in == 6'b101101;
  assign _212_ = in == 6'b101100;
  assign _213_ = in == 6'b101011;
  assign _214_ = in == 6'b101010;
  assign _215_ = in == 6'b101001;
  assign _216_ = in == 6'b101000;
  assign _217_ = in == 6'b100111;
  assign _218_ = in == 6'b100110;
  assign _219_ = in == 6'b100101;
  assign _220_ = in == 6'b100100;
  assign _221_ = in == 6'b100011;
  assign _222_ = in == 6'b100010;
  assign _223_ = in == 6'b100001;
  assign _224_ = in == 6'b100000;
  assign _225_ = in == 5'b11111;
  assign _226_ = in == 5'b11110;
  assign _227_ = in == 5'b11101;
  assign _228_ = in == 5'b11100;
  assign _229_ = in == 5'b11011;
  assign _230_ = in == 5'b11010;
  assign _231_ = in == 5'b11001;
  assign _232_ = in == 5'b11000;
  assign _233_ = in == 5'b10111;
  assign _234_ = in == 5'b10110;
  assign _235_ = in == 5'b10101;
  assign _236_ = in == 5'b10100;
  assign _237_ = in == 5'b10011;
  assign _238_ = in == 5'b10010;
  assign _239_ = in == 5'b10001;
  assign _240_ = in == 5'b10000;
  assign _241_ = in == 4'b1111;
  assign _242_ = in == 4'b1110;
  assign _243_ = in == 4'b1101;
  assign _244_ = in == 4'b1100;
  assign _245_ = in == 4'b1011;
  assign _246_ = in == 4'b1010;
  assign _247_ = in == 4'b1001;
  assign _248_ = in == 4'b1000;
  assign _249_ = in == 3'b111;
  assign _250_ = in == 3'b110;
  assign _251_ = in == 3'b101;
  assign _252_ = in == 3'b100;
  assign _253_ = in == 2'b11;
  assign _254_ = in == 2'b10;
  assign _255_ = in == 1'b1;
endmodule
