module SDP_Y_CORE_Y_alu_core(nvdla_core_clk, nvdla_core_rstn, chn_alu_in_rsc_z, chn_alu_in_rsc_vz, chn_alu_in_rsc_lz, chn_alu_op_rsc_z, chn_alu_op_rsc_vz, chn_alu_op_rsc_lz, cfg_alu_bypass_rsc_triosy_lz, cfg_alu_src_rsc_triosy_lz, cfg_alu_op_rsc_triosy_lz, cfg_alu_algo_rsc_triosy_lz, cfg_precision, chn_alu_out_rsc_z, chn_alu_out_rsc_vz, chn_alu_out_rsc_lz, chn_alu_in_rsci_oswt, chn_alu_in_rsci_oswt_unreg, chn_alu_op_rsci_oswt, chn_alu_op_rsci_oswt_unreg, cfg_alu_bypass_rsci_d, cfg_alu_src_rsci_d, cfg_alu_op_rsci_d, cfg_alu_algo_rsci_d, chn_alu_out_rsci_oswt, chn_alu_out_rsci_oswt_unreg, cfg_alu_bypass_rsc_triosy_obj_oswt, cfg_alu_src_rsc_triosy_obj_oswt, cfg_alu_op_rsc_triosy_obj_oswt, cfg_alu_algo_rsc_triosy_obj_oswt, cfg_alu_bypass_rsc_triosy_obj_oswt_unreg_pff);
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16440" *)
  wire _0000_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16440" *)
  wire _0001_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16440" *)
  wire _0002_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16440" *)
  wire _0003_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16440" *)
  wire _0004_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16440" *)
  wire _0005_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16440" *)
  wire _0006_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16440" *)
  wire _0007_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16440" *)
  wire _0008_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16440" *)
  wire _0009_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16440" *)
  wire _0010_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16440" *)
  wire _0011_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16440" *)
  wire _0012_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16440" *)
  wire _0013_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16440" *)
  wire _0014_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16440" *)
  wire _0015_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16440" *)
  wire _0016_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16525" *)
  wire [31:0] _0017_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16525" *)
  wire [31:0] _0018_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16525" *)
  wire [31:0] _0019_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16525" *)
  wire [31:0] _0020_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16525" *)
  wire [31:0] _0021_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16525" *)
  wire [31:0] _0022_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16525" *)
  wire [31:0] _0023_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16525" *)
  wire [31:0] _0024_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16542" *)
  wire [48:0] _0025_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16542" *)
  wire [48:0] _0026_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16542" *)
  wire [48:0] _0027_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16542" *)
  wire [48:0] _0028_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16576" *)
  wire [5:0] _0029_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16576" *)
  wire [5:0] _0030_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16576" *)
  wire [5:0] _0031_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16576" *)
  wire [5:0] _0032_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16593" *)
  wire [7:0] _0033_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16593" *)
  wire [7:0] _0034_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16593" *)
  wire [7:0] _0035_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16593" *)
  wire [7:0] _0036_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16593" *)
  wire [7:0] _0037_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16593" *)
  wire [7:0] _0038_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16593" *)
  wire [7:0] _0039_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16593" *)
  wire [7:0] _0040_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16695" *)
  wire [2:0] _0041_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16695" *)
  wire [2:0] _0042_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16695" *)
  wire [2:0] _0043_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16695" *)
  wire [2:0] _0044_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16701" *)
  wire [8:0] _0045_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16701" *)
  wire [8:0] _0046_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16701" *)
  wire [8:0] _0047_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16701" *)
  wire [8:0] _0048_;
  wire [22:0] _0049_;
  wire [22:0] _0050_;
  wire [22:0] _0051_;
  wire [22:0] _0052_;
  wire [22:0] _0053_;
  wire [22:0] _0054_;
  wire [22:0] _0055_;
  wire [22:0] _0056_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13741" *)
  wire [127:0] _0057_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13934" *)
  wire [127:0] _0058_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14064" *)
  wire [30:0] _0059_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14064" *)
  wire [30:0] _0060_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14064" *)
  wire [30:0] _0061_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14064" *)
  wire [30:0] _0062_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14885" *)
  wire _0063_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14532" *)
  wire _0064_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15240" *)
  wire _0065_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15240" *)
  wire _0066_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14885" *)
  wire _0067_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14532" *)
  wire _0068_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14554" *)
  wire _0069_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14885" *)
  wire _0070_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14564" *)
  wire _0071_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15232" *)
  wire _0072_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14341" *)
  wire [21:0] _0073_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14377" *)
  wire [7:0] _0074_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15028" *)
  wire _0075_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14512" *)
  wire _0076_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14732" *)
  wire [7:0] _0077_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13851" *)
  wire [7:0] _0078_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14732" *)
  wire [7:0] _0079_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13851" *)
  wire [7:0] _0080_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14732" *)
  wire [7:0] _0081_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13851" *)
  wire [7:0] _0082_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14732" *)
  wire [7:0] _0083_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13851" *)
  wire [7:0] _0084_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14212" *)
  wire _0085_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14212" *)
  wire _0086_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14212" *)
  wire _0087_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14212" *)
  wire _0088_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14732" *)
  wire [7:0] _0089_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13851" *)
  wire [7:0] _0090_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14732" *)
  wire [7:0] _0091_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13851" *)
  wire [7:0] _0092_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14732" *)
  wire [7:0] _0093_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13851" *)
  wire [7:0] _0094_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14732" *)
  wire [7:0] _0095_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13851" *)
  wire [7:0] _0096_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14668" *)
  wire [49:0] _0097_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13986" *)
  wire [49:0] _0098_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14668" *)
  wire [49:0] _0099_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13986" *)
  wire [49:0] _0100_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14668" *)
  wire [49:0] _0101_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13986" *)
  wire [49:0] _0102_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14668" *)
  wire [49:0] _0103_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13986" *)
  wire [49:0] _0104_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13821" *)
  wire _0105_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13821" *)
  wire _0106_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13821" *)
  wire _0107_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13821" *)
  wire _0108_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14416" *)
  wire _0109_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14398" *)
  wire _0110_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14359" *)
  wire _0111_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14478" *)
  wire _0112_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14093" *)
  wire [7:0] _0113_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14103" *)
  wire [7:0] _0114_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14113" *)
  wire [7:0] _0115_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14123" *)
  wire [7:0] _0116_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15158" *)
  wire [7:0] _0117_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14817" *)
  wire [7:0] _0118_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13964" *)
  wire [7:0] _0119_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15168" *)
  wire [7:0] _0120_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14828" *)
  wire [7:0] _0121_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13964" *)
  wire [7:0] _0122_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15178" *)
  wire [7:0] _0123_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14839" *)
  wire [7:0] _0124_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13964" *)
  wire [7:0] _0125_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15188" *)
  wire [7:0] _0126_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14850" *)
  wire [7:0] _0127_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13964" *)
  wire [7:0] _0128_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15140" *)
  wire _0129_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15140" *)
  wire _0130_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15140" *)
  wire _0131_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14900" *)
  wire _0132_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14313" *)
  wire _0133_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15140" *)
  wire _0134_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14900" *)
  wire _0135_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14313" *)
  wire _0136_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15140" *)
  wire _0137_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14900" *)
  wire _0138_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14313" *)
  wire _0139_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15274" *)
  wire _0140_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14900" *)
  wire _0141_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14313" *)
  wire _0142_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15282" *)
  wire _0143_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14962" *)
  wire _0144_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14496" *)
  wire _0145_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15406" *)
  wire _0146_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15406" *)
  wire _0147_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15140" *)
  wire _0148_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14900" *)
  wire _0149_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14313" *)
  wire _0150_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14450" *)
  wire _0151_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15224" *)
  wire _0152_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14875" *)
  wire _0153_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14442" *)
  wire _0154_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14468" *)
  wire [21:0] _0155_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14468" *)
  wire [7:0] _0156_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15469" *)
  wire _0157_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14952" *)
  wire [30:0] _0158_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14388" *)
  wire [30:0] _0159_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14952" *)
  wire [30:0] _0160_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14388" *)
  wire [30:0] _0161_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14944" *)
  wire [30:0] _0162_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14351" *)
  wire [30:0] _0163_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14936" *)
  wire [30:0] _0164_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14460" *)
  wire [30:0] _0165_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15262" *)
  wire [30:0] _0166_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14924" *)
  wire [30:0] _0167_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14329" *)
  wire [30:0] _0168_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15262" *)
  wire [30:0] _0169_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14924" *)
  wire [30:0] _0170_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14329" *)
  wire [30:0] _0171_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15262" *)
  wire [30:0] _0172_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14924" *)
  wire [30:0] _0173_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14329" *)
  wire [30:0] _0174_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15254" *)
  wire [30:0] _0175_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14916" *)
  wire [30:0] _0176_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14434" *)
  wire [30:0] _0177_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14682" *)
  wire _0178_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14026" *)
  wire _0179_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14690" *)
  wire _0180_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14036" *)
  wire _0181_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14698" *)
  wire _0182_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14046" *)
  wire _0183_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14660" *)
  wire _0184_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14016" *)
  wire _0185_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14981" *)
  wire [21:0] _0186_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15017" *)
  wire [7:0] _0187_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14981" *)
  wire [21:0] _0188_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14542" *)
  wire [21:0] _0189_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14995" *)
  wire [7:0] _0190_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14981" *)
  wire [21:0] _0191_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14542" *)
  wire [21:0] _0192_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15006" *)
  wire [7:0] _0193_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14981" *)
  wire [21:0] _0194_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14542" *)
  wire [21:0] _0195_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14970" *)
  wire [7:0] _0196_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13934" *)
  wire _0197_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14628" *)
  wire _0198_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14212" *)
  wire _0199_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13934" *)
  wire _0200_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14636" *)
  wire _0201_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14212" *)
  wire _0202_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13934" *)
  wire _0203_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14644" *)
  wire _0204_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14212" *)
  wire _0205_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13934" *)
  wire _0206_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14652" *)
  wire _0207_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14212" *)
  wire _0208_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15512" *)
  wire _0209_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15453" *)
  wire _0210_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15512" *)
  wire _0211_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15453" *)
  wire _0212_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15501" *)
  wire _0213_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15437" *)
  wire _0214_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15512" *)
  wire _0215_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15437" *)
  wire _0216_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15490" *)
  wire _0217_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15530" *)
  wire _0218_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15479" *)
  wire _0219_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14861" *)
  wire _0220_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14198" *)
  wire _0221_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13741" *)
  wire _0222_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15210" *)
  wire _0223_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13821" *)
  wire _0224_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13964" *)
  wire _0225_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14861" *)
  wire _0226_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14198" *)
  wire _0227_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13741" *)
  wire _0228_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15210" *)
  wire _0229_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13821" *)
  wire _0230_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13964" *)
  wire _0231_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14861" *)
  wire _0232_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14198" *)
  wire _0233_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13741" *)
  wire _0234_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15210" *)
  wire _0235_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13821" *)
  wire _0236_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13964" *)
  wire _0237_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14861" *)
  wire _0238_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14198" *)
  wire _0239_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13741" *)
  wire _0240_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15210" *)
  wire _0241_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13821" *)
  wire _0242_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13964" *)
  wire _0243_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14732" *)
  wire _0244_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13851" *)
  wire _0245_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13821" *)
  wire _0246_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14574" *)
  wire _0247_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14131" *)
  wire _0248_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14762" *)
  wire _0249_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14706" *)
  wire _0250_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13986" *)
  wire _0251_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14614" *)
  wire _0252_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14238" *)
  wire _0253_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15388" *)
  wire _0254_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14732" *)
  wire _0255_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13851" *)
  wire _0256_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15198" *)
  wire _0257_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13821" *)
  wire _0258_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14584" *)
  wire _0259_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14143" *)
  wire _0260_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14762" *)
  wire _0261_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14706" *)
  wire _0262_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13986" *)
  wire _0263_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14614" *)
  wire _0264_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14238" *)
  wire _0265_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15427" *)
  wire _0266_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15332" *)
  wire _0267_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14732" *)
  wire _0268_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13851" *)
  wire _0269_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15198" *)
  wire _0270_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14720" *)
  wire _0271_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13821" *)
  wire _0272_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14594" *)
  wire _0273_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14155" *)
  wire _0274_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14762" *)
  wire _0275_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14706" *)
  wire _0276_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13986" *)
  wire _0277_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14614" *)
  wire _0278_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14238" *)
  wire _0279_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15388" *)
  wire _0280_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14732" *)
  wire _0281_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13851" *)
  wire _0282_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15198" *)
  wire _0283_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14720" *)
  wire _0284_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13821" *)
  wire _0285_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14604" *)
  wire _0286_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14167" *)
  wire _0287_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14762" *)
  wire _0288_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14706" *)
  wire _0289_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13986" *)
  wire _0290_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14614" *)
  wire _0291_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14238" *)
  wire _0292_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15388" *)
  wire _0293_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13934" *)
  wire _0294_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14064" *)
  wire _0295_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14512" *)
  wire _0296_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14809" *)
  wire [1:0] _0297_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14792" *)
  wire [1:0] _0298_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14784" *)
  wire [1:0] _0299_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13775" *)
  wire [1:0] _0300_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13917" *)
  wire [1:0] _0301_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14056" *)
  wire [1:0] _0302_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14504" *)
  wire [1:0] _0303_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13759" *)
  wire [1:0] _0304_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13784" *)
  wire [31:0] _0305_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14800" *)
  wire _0306_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13794" *)
  wire _0307_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13620" *)
  wire _0308_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13634" *)
  wire _0309_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13620" *)
  wire _0310_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13724" *)
  wire _0311_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13642" *)
  wire _0312_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13669" *)
  wire [21:0] _0313_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13669" *)
  wire [7:0] _0314_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13669" *)
  wire _0315_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13657" *)
  wire [21:0] _0316_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13669" *)
  wire [7:0] _0317_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13669" *)
  wire _0318_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13642" *)
  wire _0319_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13657" *)
  wire [21:0] _0320_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13669" *)
  wire [7:0] _0321_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13669" *)
  wire _0322_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13697" *)
  wire _0323_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13706" *)
  wire [21:0] _0324_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13706" *)
  wire [7:0] _0325_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13669" *)
  wire _0326_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13642" *)
  wire _0327_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13620" *)
  wire _0328_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13917" *)
  wire [30:0] _0329_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13917" *)
  wire [30:0] _0330_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13917" *)
  wire [30:0] _0331_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13917" *)
  wire [30:0] _0332_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15090" *)
  wire [22:0] _0333_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15050" *)
  wire [22:0] _0334_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15126" *)
  wire [7:0] _0335_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14426" *)
  wire [7:0] _0336_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15099" *)
  wire [22:0] _0337_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15060" *)
  wire [22:0] _0338_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15126" *)
  wire [7:0] _0339_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14408" *)
  wire [7:0] _0340_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15108" *)
  wire [22:0] _0341_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15070" *)
  wire [22:0] _0342_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15126" *)
  wire [7:0] _0343_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14369" *)
  wire [7:0] _0344_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15117" *)
  wire [22:0] _0345_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15080" *)
  wire [22:0] _0346_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15126" *)
  wire [7:0] _0347_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14488" *)
  wire [7:0] _0348_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13741" *)
  wire _0349_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13934" *)
  wire _0350_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14064" *)
  wire _0351_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14512" *)
  wire _0352_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13804" *)
  wire _0353_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13934" *)
  wire _0354_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14064" *)
  wire _0355_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14512" *)
  wire _0356_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13733" *)
  wire _0357_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13813" *)
  wire _0358_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13956" *)
  wire _0359_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14084" *)
  wire _0360_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15028" *)
  wire _0361_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14512" *)
  wire _0362_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15028" *)
  wire _0363_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14512" *)
  wire _0364_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15028" *)
  wire _0365_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14512" *)
  wire _0366_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14188" *)
  wire [22:0] _0367_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14179" *)
  wire [7:0] _0368_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14303" *)
  wire [22:0] _0369_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14294" *)
  wire [7:0] _0370_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14284" *)
  wire [22:0] _0371_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14275" *)
  wire [7:0] _0372_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14265" *)
  wire [22:0] _0373_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14256" *)
  wire [7:0] _0374_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13851" *)
  wire _0375_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13851" *)
  wire _0376_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13851" *)
  wire _0377_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13851" *)
  wire _0378_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15301" *)
  wire [30:0] _0379_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15290" *)
  wire _0380_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15322" *)
  wire [30:0] _0381_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15311" *)
  wire _0382_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15355" *)
  wire [30:0] _0383_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15344" *)
  wire _0384_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15377" *)
  wire [30:0] _0385_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15366" *)
  wire _0386_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13767" *)
  wire [1:0] _0387_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13620" *)
  wire _0388_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13716" *)
  wire _0389_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13642" *)
  wire _0390_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13642" *)
  wire _0391_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13642" *)
  wire _0392_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13697" *)
  wire _0393_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13794" *)
  wire _0394_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13851" *)
  wire _0395_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13851" *)
  wire _0396_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13851" *)
  wire _0397_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13851" *)
  wire _0398_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13851" *)
  wire _0399_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13851" *)
  wire _0400_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13851" *)
  wire _0401_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13851" *)
  wire _0402_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13986" *)
  wire _0403_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13986" *)
  wire _0404_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13986" *)
  wire _0405_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13986" *)
  wire _0406_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14016" *)
  wire _0407_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14026" *)
  wire _0408_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14036" *)
  wire _0409_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14046" *)
  wire _0410_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14131" *)
  wire _0411_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14143" *)
  wire _0412_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14155" *)
  wire _0413_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14167" *)
  wire _0414_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14238" *)
  wire _0415_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14238" *)
  wire _0416_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14238" *)
  wire _0417_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14238" *)
  wire _0418_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14359" *)
  wire _0419_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14398" *)
  wire _0420_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14416" *)
  wire _0421_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14478" *)
  wire _0422_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14564" *)
  wire _0423_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14720" *)
  wire _0424_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14720" *)
  wire _0425_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14875" *)
  wire _0426_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14885" *)
  wire _0427_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14885" *)
  wire _0428_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14885" *)
  wire _0429_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15332" *)
  wire _0430_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15530" *)
  wire _0431_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14341" *)
  wire [21:0] _0432_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15050" *)
  wire [22:0] _0433_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15060" *)
  wire [22:0] _0434_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15070" *)
  wire [22:0] _0435_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15080" *)
  wire [22:0] _0436_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13775" *)
  wire [1:0] _0437_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13917" *)
  wire [30:0] _0438_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13784" *)
  wire [31:0] _0439_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13986" *)
  wire [49:0] _0440_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13986" *)
  wire [49:0] _0441_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13986" *)
  wire [49:0] _0442_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13986" *)
  wire [49:0] _0443_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13851" *)
  wire [7:0] _0444_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13851" *)
  wire [7:0] _0445_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13851" *)
  wire [7:0] _0446_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13851" *)
  wire [7:0] _0447_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13851" *)
  wire [7:0] _0448_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13851" *)
  wire [7:0] _0449_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13851" *)
  wire [7:0] _0450_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13851" *)
  wire [7:0] _0451_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14093" *)
  wire [7:0] _0452_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14103" *)
  wire [7:0] _0453_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14113" *)
  wire [7:0] _0454_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14377" *)
  wire [7:0] _0455_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15158" *)
  wire [7:0] _0456_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15168" *)
  wire [7:0] _0457_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15178" *)
  wire [7:0] _0458_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15188" *)
  wire [7:0] _0459_;
  wire [8:0] _0460_;
  wire [23:0] _0461_;
  wire [23:0] _0462_;
  wire [8:0] _0463_;
  wire [23:0] _0464_;
  wire [8:0] _0465_;
  wire [8:0] _0466_;
  wire [8:0] _0467_;
  wire [8:0] _0468_;
  wire [8:0] _0469_;
  wire [8:0] _0470_;
  wire [8:0] _0471_;
  wire [8:0] _0472_;
  wire [23:0] _0473_;
  wire [8:0] _0474_;
  wire [8:0] _0475_;
  wire [23:0] _0476_;
  wire [23:0] _0477_;
  wire [23:0] _0478_;
  wire [23:0] _0479_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12265" *)
  wire _0480_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12272" *)
  wire _0481_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12272" *)
  wire _0482_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12275" *)
  wire _0483_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12278" *)
  wire _0484_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12282" *)
  wire _0485_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12287" *)
  wire _0486_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12288" *)
  wire _0487_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12288" *)
  wire _0488_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12289" *)
  wire _0489_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12290" *)
  wire _0490_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12291" *)
  wire _0491_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12295" *)
  wire _0492_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12298" *)
  wire _0493_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12312" *)
  wire _0494_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12333" *)
  wire _0495_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12427" *)
  wire _0496_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12427" *)
  wire _0497_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12427" *)
  wire _0498_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12447" *)
  wire _0499_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12450" *)
  wire _0500_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12455" *)
  wire _0501_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12456" *)
  wire _0502_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12456" *)
  wire _0503_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12456" *)
  wire _0504_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12458" *)
  wire _0505_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12460" *)
  wire _0506_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12462" *)
  wire _0507_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12464" *)
  wire _0508_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12471" *)
  wire _0509_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12471" *)
  wire _0510_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12474" *)
  wire _0511_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12481" *)
  wire _0512_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12508" *)
  wire _0513_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12509" *)
  wire _0514_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12509" *)
  wire _0515_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12510" *)
  wire _0516_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12510" *)
  wire _0517_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12510" *)
  wire _0518_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12511" *)
  wire _0519_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12517" *)
  wire _0520_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12524" *)
  wire _0521_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12524" *)
  wire _0522_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12528" *)
  wire _0523_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12528" *)
  wire _0524_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12529" *)
  wire _0525_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12529" *)
  wire _0526_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12530" *)
  wire _0527_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12530" *)
  wire _0528_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12536" *)
  wire _0529_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12537" *)
  wire _0530_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12537" *)
  wire _0531_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12537" *)
  wire _0532_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12571" *)
  wire _0533_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12572" *)
  wire _0534_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12600" *)
  wire _0535_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12603" *)
  wire _0536_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12603" *)
  wire _0537_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12623" *)
  wire _0538_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12625" *)
  wire _0539_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12625" *)
  wire _0540_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12627" *)
  wire _0541_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12629" *)
  wire _0542_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12659" *)
  wire _0543_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12669" *)
  wire _0544_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12680" *)
  wire _0545_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12691" *)
  wire _0546_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12823" *)
  wire _0547_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12974" *)
  wire _0548_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12976" *)
  wire _0549_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12976" *)
  wire _0550_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12978" *)
  wire _0551_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12980" *)
  wire _0552_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13006" *)
  wire _0553_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13006" *)
  wire _0554_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13006" *)
  wire _0555_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13007" *)
  wire _0556_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13008" *)
  wire _0557_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13008" *)
  wire _0558_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13009" *)
  wire _0559_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13137" *)
  wire _0560_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13195" *)
  wire _0561_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13286" *)
  wire _0562_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13290" *)
  wire _0563_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13294" *)
  wire _0564_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13294" *)
  wire _0565_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13294" *)
  wire _0566_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13295" *)
  wire _0567_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13295" *)
  wire _0568_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13352" *)
  wire _0569_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13383" *)
  wire _0570_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13383" *)
  wire _0571_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13384" *)
  wire _0572_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13384" *)
  wire _0573_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13384" *)
  wire _0574_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13385" *)
  wire _0575_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13424" *)
  wire _0576_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13447" *)
  wire _0577_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13447" *)
  wire _0578_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13450" *)
  wire _0579_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13450" *)
  wire _0580_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13450" *)
  wire _0581_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13458" *)
  wire _0582_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13461" *)
  wire _0583_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13465" *)
  wire _0584_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13465" *)
  wire _0585_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13466" *)
  wire _0586_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13474" *)
  wire _0587_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13505" *)
  wire _0588_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13513" *)
  wire _0589_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13514" *)
  wire _0590_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13521" *)
  wire _0591_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13522" *)
  wire _0592_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13522" *)
  wire _0593_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13530" *)
  wire _0594_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13533" *)
  wire _0595_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13537" *)
  wire _0596_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13537" *)
  wire _0597_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13538" *)
  wire _0598_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13539" *)
  wire _0599_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13542" *)
  wire _0600_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13542" *)
  wire _0601_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13542" *)
  wire _0602_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13543" *)
  wire _0603_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13543" *)
  wire _0604_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13543" *)
  wire _0605_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13545" *)
  wire _0606_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13545" *)
  wire _0607_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13545" *)
  wire _0608_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13546" *)
  wire _0609_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13546" *)
  wire _0610_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13547" *)
  wire _0611_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13547" *)
  wire _0612_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13547" *)
  wire _0613_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13550" *)
  wire _0614_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13551" *)
  wire _0615_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13552" *)
  wire _0616_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13553" *)
  wire _0617_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13553" *)
  wire _0618_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13555" *)
  wire _0619_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13557" *)
  wire _0620_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13559" *)
  wire _0621_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13578" *)
  wire _0622_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13578" *)
  wire _0623_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13579" *)
  wire _0624_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13583" *)
  wire _0625_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13583" *)
  wire _0626_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13585" *)
  wire _0627_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13587" *)
  wire _0628_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13587" *)
  wire _0629_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13628" *)
  wire _0630_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13638" *)
  wire _0631_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13701" *)
  wire _0632_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13720" *)
  wire _0633_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13728" *)
  wire _0634_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13729" *)
  wire _0635_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13729" *)
  wire _0636_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13729" *)
  wire _0637_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13737" *)
  wire _0638_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13763" *)
  wire _0639_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13771" *)
  wire _0640_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13779" *)
  wire _0641_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13788" *)
  wire _0642_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13788" *)
  wire _0643_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13798" *)
  wire _0644_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13799" *)
  wire _0645_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13809" *)
  wire _0646_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13817" *)
  wire _0647_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13960" *)
  wire _0648_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14021" *)
  wire _0649_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14031" *)
  wire _0650_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14041" *)
  wire _0651_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14051" *)
  wire _0652_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14060" *)
  wire _0653_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14088" *)
  wire _0654_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14089" *)
  wire _0655_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14097" *)
  wire _0656_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14098" *)
  wire _0657_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14108" *)
  wire _0658_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14118" *)
  wire _0659_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14127" *)
  wire _0660_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14137" *)
  wire _0661_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14149" *)
  wire _0662_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14161" *)
  wire _0663_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14173" *)
  wire _0664_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14183" *)
  wire _0665_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14183" *)
  wire _0666_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14183" *)
  wire _0667_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14184" *)
  wire _0668_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14184" *)
  wire _0669_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14192" *)
  wire _0670_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14193" *)
  wire _0671_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14193" *)
  wire _0672_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14193" *)
  wire _0673_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14194" *)
  wire _0674_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14194" *)
  wire _0675_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14229" *)
  wire _0676_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14231" *)
  wire _0677_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14233" *)
  wire _0678_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14235" *)
  wire _0679_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14260" *)
  wire _0680_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14261" *)
  wire _0681_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14261" *)
  wire _0682_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14269" *)
  wire _0683_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14270" *)
  wire _0684_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14270" *)
  wire _0685_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14270" *)
  wire _0686_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14271" *)
  wire _0687_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14271" *)
  wire _0688_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14279" *)
  wire _0689_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14280" *)
  wire _0690_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14280" *)
  wire _0691_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14288" *)
  wire _0692_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14289" *)
  wire _0693_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14289" *)
  wire _0694_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14289" *)
  wire _0695_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14290" *)
  wire _0696_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14290" *)
  wire _0697_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14298" *)
  wire _0698_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14299" *)
  wire _0699_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14299" *)
  wire _0700_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14307" *)
  wire _0701_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14308" *)
  wire _0702_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14308" *)
  wire _0703_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14308" *)
  wire _0704_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14309" *)
  wire _0705_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14309" *)
  wire _0706_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14345" *)
  wire _0707_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14346" *)
  wire _0708_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14346" *)
  wire _0709_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14355" *)
  wire _0710_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14363" *)
  wire _0711_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14364" *)
  wire _0712_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14364" *)
  wire _0713_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14373" *)
  wire _0714_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14383" *)
  wire _0715_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14383" *)
  wire _0716_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14383" *)
  wire _0717_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14402" *)
  wire _0718_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14403" *)
  wire _0719_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14403" *)
  wire _0720_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14412" *)
  wire _0721_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14420" *)
  wire _0722_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14421" *)
  wire _0723_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14421" *)
  wire _0724_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14430" *)
  wire _0725_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14438" *)
  wire _0726_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14446" *)
  wire _0727_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14456" *)
  wire _0728_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14456" *)
  wire _0729_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14456" *)
  wire _0730_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14456" *)
  wire _0731_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14464" *)
  wire _0732_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14482" *)
  wire _0733_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14483" *)
  wire _0734_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14483" *)
  wire _0735_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14492" *)
  wire _0736_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14500" *)
  wire _0737_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14508" *)
  wire _0738_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14558" *)
  wire _0739_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14569" *)
  wire _0740_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14579" *)
  wire _0741_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14589" *)
  wire _0742_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14599" *)
  wire _0743_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14609" *)
  wire _0744_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14632" *)
  wire _0745_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14640" *)
  wire _0746_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14648" *)
  wire _0747_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14656" *)
  wire _0748_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14664" *)
  wire _0749_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14664" *)
  wire _0750_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14686" *)
  wire _0751_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14694" *)
  wire _0752_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14702" *)
  wire _0753_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14788" *)
  wire _0754_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14796" *)
  wire _0755_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14805" *)
  wire _0756_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14813" *)
  wire _0757_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14821" *)
  wire _0758_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14821" *)
  wire _0759_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14832" *)
  wire _0760_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14832" *)
  wire _0761_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14843" *)
  wire _0762_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14843" *)
  wire _0763_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14854" *)
  wire _0764_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14854" *)
  wire _0765_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14880" *)
  wire _0766_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14920" *)
  wire _0767_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14940" *)
  wire _0768_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14948" *)
  wire _0769_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14966" *)
  wire _0770_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14974" *)
  wire _0771_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14975" *)
  wire _0772_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15000" *)
  wire _0773_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15011" *)
  wire _0774_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15022" *)
  wire _0775_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15055" *)
  wire _0776_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15065" *)
  wire _0777_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15075" *)
  wire _0778_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15085" *)
  wire _0779_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15095" *)
  wire _0780_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15104" *)
  wire _0781_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15113" *)
  wire _0782_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15122" *)
  wire _0783_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15154" *)
  wire _0784_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15155" *)
  wire _0785_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15163" *)
  wire _0786_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15163" *)
  wire _0787_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15163" *)
  wire _0788_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15173" *)
  wire _0789_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15173" *)
  wire _0790_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15173" *)
  wire _0791_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15183" *)
  wire _0792_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15183" *)
  wire _0793_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15183" *)
  wire _0794_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15193" *)
  wire _0795_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15193" *)
  wire _0796_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15193" *)
  wire _0797_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15228" *)
  wire _0798_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15236" *)
  wire _0799_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15258" *)
  wire _0800_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15278" *)
  wire _0801_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15286" *)
  wire _0802_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15294" *)
  wire _0803_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15295" *)
  wire _0804_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15295" *)
  wire _0805_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15296" *)
  wire _0806_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15296" *)
  wire _0807_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15296" *)
  wire _0808_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15296" *)
  wire _0809_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15297" *)
  wire _0810_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15297" *)
  wire _0811_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15297" *)
  wire _0812_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15305" *)
  wire _0813_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15306" *)
  wire _0814_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15306" *)
  wire _0815_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15306" *)
  wire _0816_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15306" *)
  wire _0817_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15307" *)
  wire _0818_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15307" *)
  wire _0819_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15316" *)
  wire _0820_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15316" *)
  wire _0821_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15317" *)
  wire _0822_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15317" *)
  wire _0823_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15317" *)
  wire _0824_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15317" *)
  wire _0825_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15318" *)
  wire _0826_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15318" *)
  wire _0827_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15318" *)
  wire _0828_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15326" *)
  wire _0829_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15327" *)
  wire _0830_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15327" *)
  wire _0831_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15327" *)
  wire _0832_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15327" *)
  wire _0833_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15328" *)
  wire _0834_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15328" *)
  wire _0835_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15337" *)
  wire _0836_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15338" *)
  wire _0837_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15338" *)
  wire _0838_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15349" *)
  wire _0839_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15349" *)
  wire _0840_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15350" *)
  wire _0841_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15350" *)
  wire _0842_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15350" *)
  wire _0843_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15350" *)
  wire _0844_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15351" *)
  wire _0845_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15351" *)
  wire _0846_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15351" *)
  wire _0847_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15359" *)
  wire _0848_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15359" *)
  wire _0849_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15360" *)
  wire _0850_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15360" *)
  wire _0851_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15360" *)
  wire _0852_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15361" *)
  wire _0853_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15361" *)
  wire _0854_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15361" *)
  wire _0855_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15362" *)
  wire _0856_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15370" *)
  wire _0857_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15370" *)
  wire _0858_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15371" *)
  wire _0859_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15371" *)
  wire _0860_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15371" *)
  wire _0861_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15371" *)
  wire _0862_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15372" *)
  wire _0863_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15372" *)
  wire _0864_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15381" *)
  wire _0865_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15382" *)
  wire _0866_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15382" *)
  wire _0867_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15382" *)
  wire _0868_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15383" *)
  wire _0869_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15383" *)
  wire _0870_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15383" *)
  wire _0871_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15384" *)
  wire _0872_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15432" *)
  wire _0873_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15475" *)
  wire _0874_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15475" *)
  wire _0875_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15483" *)
  wire _0876_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15484" *)
  wire _0877_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15495" *)
  wire _0878_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15506" *)
  wire _0879_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15534" *)
  wire _0880_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15534" *)
  wire _0881_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15567" *)
  wire _0882_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15569" *)
  wire _0883_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15569" *)
  wire _0884_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15571" *)
  wire _0885_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15573" *)
  wire _0886_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15587" *)
  wire _0887_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15589" *)
  wire _0888_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15589" *)
  wire _0889_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15591" *)
  wire _0890_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15593" *)
  wire _0891_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15616" *)
  wire _0892_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15775" *)
  wire _0893_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15783" *)
  wire _0894_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15791" *)
  wire _0895_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15799" *)
  wire _0896_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15859" *)
  wire _0897_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15859" *)
  wire _0898_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15887" *)
  wire _0899_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15897" *)
  wire _0900_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15907" *)
  wire _0901_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15917" *)
  wire _0902_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15943" *)
  wire _0903_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15950" *)
  wire _0904_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15952" *)
  wire _0905_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15954" *)
  wire _0906_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16047" *)
  wire _0907_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16047" *)
  wire _0908_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16049" *)
  wire _0909_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16049" *)
  wire _0910_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16055" *)
  wire _0911_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16055" *)
  wire _0912_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16057" *)
  wire _0913_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16057" *)
  wire _0914_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16070" *)
  wire _0915_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16074" *)
  wire _0916_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16080" *)
  wire _0917_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16084" *)
  wire _0918_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16115" *)
  wire _0919_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16115" *)
  wire _0920_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16118" *)
  wire _0921_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16118" *)
  wire _0922_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16129" *)
  wire _0923_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16129" *)
  wire _0924_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16132" *)
  wire _0925_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16132" *)
  wire _0926_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16141" *)
  wire _0927_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16159" *)
  wire _0928_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16163" *)
  wire _0929_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16170" *)
  wire _0930_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16174" *)
  wire _0931_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16264" *)
  wire _0932_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16264" *)
  wire _0933_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16264" *)
  wire _0934_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16264" *)
  wire _0935_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16264" *)
  wire _0936_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16264" *)
  wire _0937_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16264" *)
  wire _0938_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16264" *)
  wire _0939_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16264" *)
  wire _0940_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16264" *)
  wire _0941_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16264" *)
  wire _0942_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16265" *)
  wire _0943_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16265" *)
  wire _0944_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16265" *)
  wire _0945_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16265" *)
  wire _0946_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16265" *)
  wire _0947_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16265" *)
  wire _0948_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16265" *)
  wire _0949_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16265" *)
  wire _0950_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16265" *)
  wire _0951_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16265" *)
  wire _0952_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16265" *)
  wire _0953_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16266" *)
  wire _0954_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16266" *)
  wire _0955_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16266" *)
  wire _0956_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16266" *)
  wire _0957_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16266" *)
  wire _0958_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16266" *)
  wire _0959_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16266" *)
  wire _0960_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16266" *)
  wire _0961_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16266" *)
  wire _0962_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16266" *)
  wire _0963_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16266" *)
  wire _0964_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16278" *)
  wire _0965_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16278" *)
  wire _0966_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16278" *)
  wire _0967_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16278" *)
  wire _0968_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16278" *)
  wire _0969_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16278" *)
  wire _0970_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16278" *)
  wire _0971_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16278" *)
  wire _0972_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16278" *)
  wire _0973_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16278" *)
  wire _0974_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16279" *)
  wire _0975_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16279" *)
  wire _0976_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16279" *)
  wire _0977_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16279" *)
  wire _0978_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16279" *)
  wire _0979_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16279" *)
  wire _0980_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16279" *)
  wire _0981_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16279" *)
  wire _0982_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16279" *)
  wire _0983_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16279" *)
  wire _0984_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16280" *)
  wire _0985_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16280" *)
  wire _0986_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16280" *)
  wire _0987_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16280" *)
  wire _0988_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16280" *)
  wire _0989_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16280" *)
  wire _0990_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16280" *)
  wire _0991_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16280" *)
  wire _0992_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16280" *)
  wire _0993_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16280" *)
  wire _0994_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16281" *)
  wire _0995_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16281" *)
  wire _0996_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16281" *)
  wire _0997_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16281" *)
  wire _0998_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16281" *)
  wire _0999_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16281" *)
  wire _1000_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16281" *)
  wire _1001_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16281" *)
  wire _1002_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16281" *)
  wire _1003_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16281" *)
  wire _1004_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16294" *)
  wire _1005_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16294" *)
  wire _1006_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16295" *)
  wire _1007_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16295" *)
  wire _1008_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16296" *)
  wire _1009_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16296" *)
  wire _1010_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16297" *)
  wire _1011_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16297" *)
  wire _1012_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16298" *)
  wire _1013_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16298" *)
  wire _1014_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16313" *)
  wire _1015_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16313" *)
  wire _1016_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16314" *)
  wire _1017_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16314" *)
  wire _1018_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16315" *)
  wire _1019_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16315" *)
  wire _1020_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16316" *)
  wire _1021_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16316" *)
  wire _1022_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16317" *)
  wire _1023_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16317" *)
  wire _1024_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16318" *)
  wire _1025_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16318" *)
  wire _1026_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16319" *)
  wire _1027_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16319" *)
  wire _1028_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16330" *)
  wire [21:0] _1029_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16330" *)
  wire [21:0] _1030_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16330" *)
  wire [21:0] _1031_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16330" *)
  wire [21:0] _1032_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16330" *)
  wire [21:0] _1033_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16331" *)
  wire [21:0] _1034_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16331" *)
  wire [21:0] _1035_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16331" *)
  wire [21:0] _1036_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16331" *)
  wire [21:0] _1037_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16331" *)
  wire [21:0] _1038_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16332" *)
  wire [21:0] _1039_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16332" *)
  wire [21:0] _1040_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16332" *)
  wire [21:0] _1041_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16332" *)
  wire [21:0] _1042_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16332" *)
  wire [21:0] _1043_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16344" *)
  wire [21:0] _1044_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16345" *)
  wire [21:0] _1045_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16346" *)
  wire [21:0] _1046_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16347" *)
  wire [21:0] _1047_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16358" *)
  wire [30:0] _1048_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16358" *)
  wire [30:0] _1049_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16358" *)
  wire [30:0] _1050_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16358" *)
  wire [30:0] _1051_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16359" *)
  wire [30:0] _1052_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16359" *)
  wire [30:0] _1053_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16359" *)
  wire [30:0] _1054_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16359" *)
  wire [30:0] _1055_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16360" *)
  wire [30:0] _1056_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16360" *)
  wire [30:0] _1057_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16360" *)
  wire [30:0] _1058_;
  wire [6:0] _1059_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16371" *)
  wire [7:0] _1060_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16371" *)
  wire [7:0] _1061_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16371" *)
  wire [7:0] _1062_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16371" *)
  wire [7:0] _1063_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16371" *)
  wire [7:0] _1064_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16371" *)
  wire [7:0] _1065_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16371" *)
  wire [7:0] _1066_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16371" *)
  wire [7:0] _1067_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16371" *)
  wire [7:0] _1068_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16371" *)
  wire [7:0] _1069_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16371" *)
  wire [7:0] _1070_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16371" *)
  wire [7:0] _1071_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16371" *)
  wire [7:0] _1072_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16371" *)
  wire [7:0] _1073_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16371" *)
  wire [7:0] _1074_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16371" *)
  wire [7:0] _1075_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16372" *)
  wire [7:0] _1076_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16372" *)
  wire [7:0] _1077_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16372" *)
  wire [7:0] _1078_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16372" *)
  wire [7:0] _1079_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16372" *)
  wire [7:0] _1080_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16372" *)
  wire [7:0] _1081_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16372" *)
  wire [7:0] _1082_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16372" *)
  wire [7:0] _1083_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16372" *)
  wire [7:0] _1084_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16372" *)
  wire [7:0] _1085_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16372" *)
  wire [7:0] _1086_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16372" *)
  wire [7:0] _1087_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16372" *)
  wire [7:0] _1088_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16372" *)
  wire [7:0] _1089_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16372" *)
  wire [7:0] _1090_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16372" *)
  wire [7:0] _1091_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16373" *)
  wire [7:0] _1092_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16373" *)
  wire [7:0] _1093_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16373" *)
  wire [7:0] _1094_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16373" *)
  wire [7:0] _1095_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16373" *)
  wire [7:0] _1096_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16373" *)
  wire [7:0] _1097_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16373" *)
  wire [7:0] _1098_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16373" *)
  wire [7:0] _1099_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16373" *)
  wire [7:0] _1100_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16373" *)
  wire [7:0] _1101_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16373" *)
  wire [7:0] _1102_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16373" *)
  wire [7:0] _1103_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16373" *)
  wire [7:0] _1104_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16373" *)
  wire [7:0] _1105_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16373" *)
  wire [7:0] _1106_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16373" *)
  wire [7:0] _1107_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16387" *)
  wire [7:0] _1108_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16387" *)
  wire [7:0] _1109_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16388" *)
  wire [7:0] _1110_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16388" *)
  wire [7:0] _1111_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16389" *)
  wire [7:0] _1112_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16389" *)
  wire [7:0] _1113_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16390" *)
  wire [7:0] _1114_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16390" *)
  wire [7:0] _1115_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16391" *)
  wire [7:0] _1116_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16391" *)
  wire [7:0] _1117_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16392" *)
  wire [7:0] _1118_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16392" *)
  wire [7:0] _1119_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16407" *)
  wire [7:0] _1120_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16408" *)
  wire [7:0] _1121_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16409" *)
  wire [7:0] _1122_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16410" *)
  wire [7:0] _1123_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16411" *)
  wire [7:0] _1124_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16412" *)
  wire [7:0] _1125_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16413" *)
  wire [7:0] _1126_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16429" *)
  wire [7:0] _1127_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16430" *)
  wire [7:0] _1128_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16431" *)
  wire [7:0] _1129_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16432" *)
  wire [7:0] _1130_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16433" *)
  wire [7:0] _1131_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16434" *)
  wire [7:0] _1132_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16435" *)
  wire [7:0] _1133_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16436" *)
  wire [7:0] _1134_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16360" *)
  wire [30:0] _1135_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13206" *)
  wire [7:0] _1136_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13221" *)
  wire [7:0] _1137_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12820" *)
  wire _1138_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12821" *)
  wire _1139_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12880" *)
  wire _1140_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12900" *)
  wire _1141_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12920" *)
  wire _1142_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12940" *)
  wire _1143_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13137" *)
  wire _1144_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13529" *)
  wire _1145_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13532" *)
  wire _1146_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12281" *)
  wire _1147_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12336" *)
  wire _1148_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12546" *)
  wire _1149_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12670" *)
  wire _1150_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12671" *)
  wire _1151_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12681" *)
  wire _1152_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12682" *)
  wire _1153_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12692" *)
  wire _1154_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12693" *)
  wire _1155_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12759" *)
  wire _1156_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12760" *)
  wire _1157_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12761" *)
  wire _1158_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12762" *)
  wire _1159_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12811" *)
  wire _1160_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12812" *)
  wire _1161_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12813" *)
  wire _1162_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12814" *)
  wire _1163_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12826" *)
  wire _1164_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12827" *)
  wire _1165_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13256" *)
  wire _1166_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13270" *)
  wire _1167_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13436" *)
  wire _1168_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13534" *)
  wire _1169_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13535" *)
  wire _1170_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13536" *)
  wire _1171_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15246" *)
  wire _1172_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15249" *)
  wire _1173_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11932" *)
  wire [6:0] _1174_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11943" *)
  wire [6:0] _1175_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11954" *)
  wire [6:0] _1176_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11965" *)
  wire [6:0] _1177_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11976" *)
  wire [6:0] _1178_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11987" *)
  wire [6:0] _1179_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11998" *)
  wire [6:0] _1180_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12009" *)
  wire [6:0] _1181_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12267" *)
  wire _1182_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12269" *)
  wire _1183_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12273" *)
  wire _1184_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12275" *)
  wire _1185_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12275" *)
  wire _1186_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12278" *)
  wire _1187_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12280" *)
  wire _1188_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12285" *)
  wire _1189_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12289" *)
  wire _1190_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12291" *)
  wire _1191_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12296" *)
  wire _1192_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12298" *)
  wire _1193_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12299" *)
  wire _1194_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12311" *)
  wire _1195_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12312" *)
  wire _1196_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12314" *)
  wire _1197_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12315" *)
  wire _1198_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12316" *)
  wire _1199_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12324" *)
  wire _1200_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12333" *)
  wire _1201_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12336" *)
  wire _1202_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12337" *)
  wire _1203_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12342" *)
  wire _1204_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12343" *)
  wire _1205_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12345" *)
  wire _1206_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12349" *)
  wire _1207_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12356" *)
  wire _1208_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12364" *)
  wire _1209_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12380" *)
  wire _1210_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12396" *)
  wire _1211_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12408" *)
  wire _1212_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12409" *)
  wire _1213_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12416" *)
  wire _1214_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12417" *)
  wire _1215_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12418" *)
  wire _1216_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12421" *)
  wire _1217_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12422" *)
  wire _1218_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12423" *)
  wire _1219_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12429" *)
  wire _1220_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12432" *)
  wire _1221_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12434" *)
  wire _1222_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12435" *)
  wire _1223_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12439" *)
  wire _1224_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12441" *)
  wire _1225_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12442" *)
  wire _1226_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12447" *)
  wire _1227_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12450" *)
  wire _1228_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12451" *)
  wire _1229_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12456" *)
  wire _1230_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12458" *)
  wire _1231_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12460" *)
  wire _1232_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12462" *)
  wire _1233_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12464" *)
  wire _1234_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12465" *)
  wire _1235_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12471" *)
  wire _1236_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12474" *)
  wire _1237_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12481" *)
  wire _1238_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12482" *)
  wire _1239_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12485" *)
  wire _1240_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12489" *)
  wire _1241_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12492" *)
  wire _1242_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12494" *)
  wire _1243_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12496" *)
  wire _1244_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12504" *)
  wire _1245_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12517" *)
  wire _1246_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12517" *)
  wire _1247_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12519" *)
  wire _1248_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12519" *)
  wire _1249_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12520" *)
  wire _1250_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12520" *)
  wire _1251_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12524" *)
  wire _1252_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12533" *)
  wire _1253_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12539" *)
  wire _1254_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12548" *)
  wire _1255_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12570" *)
  wire _1256_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12573" *)
  wire _1257_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12588" *)
  wire _1258_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12600" *)
  wire _1259_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12622" *)
  wire _1260_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12624" *)
  wire _1261_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12628" *)
  wire _1262_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12658" *)
  wire _1263_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12668" *)
  wire _1264_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12679" *)
  wire _1265_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12690" *)
  wire _1266_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12703" *)
  wire _1267_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12715" *)
  wire _1268_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12727" *)
  wire _1269_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12739" *)
  wire _1270_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12751" *)
  wire _1271_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12752" *)
  wire _1272_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12753" *)
  wire _1273_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12754" *)
  wire _1274_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12811" *)
  wire _1275_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12813" *)
  wire _1276_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12823" *)
  wire _1277_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12973" *)
  wire _1278_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12975" *)
  wire _1279_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12979" *)
  wire _1280_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13000" *)
  wire _1281_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13002" *)
  wire _1282_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13006" *)
  wire _1283_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13077" *)
  wire _1284_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13084" *)
  wire _1285_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13091" *)
  wire _1286_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13098" *)
  wire _1287_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13125" *)
  wire _1288_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13125" *)
  wire _1289_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13126" *)
  wire _1290_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13132" *)
  wire _1291_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13132" *)
  wire _1292_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13137" *)
  wire _1293_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13146" *)
  wire _1294_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13147" *)
  wire _1295_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13148" *)
  wire _1296_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13160" *)
  wire _1297_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13161" *)
  wire _1298_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13162" *)
  wire _1299_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13178" *)
  wire _1300_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13185" *)
  wire _1301_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13188" *)
  wire _1302_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13195" *)
  wire _1303_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13198" *)
  wire _1304_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13199" *)
  wire _1305_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13200" *)
  wire _1306_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13201" *)
  wire _1307_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13202" *)
  wire _1308_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13203" *)
  wire _1309_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13204" *)
  wire _1310_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13205" *)
  wire _1311_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13211" *)
  wire [7:0] _1312_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13216" *)
  wire [7:0] _1313_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13226" *)
  wire _1314_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13274" *)
  wire _1315_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13280" *)
  wire _1316_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13286" *)
  wire _1317_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13295" *)
  wire _1318_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13323" *)
  wire _1319_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13329" *)
  wire _1320_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13332" *)
  wire _1321_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13334" *)
  wire _1322_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13352" *)
  wire _1323_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13412" *)
  wire _1324_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13427" *)
  wire _1325_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13447" *)
  wire _1326_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13450" *)
  wire _1327_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13450" *)
  wire _1328_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13451" *)
  wire _1329_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13452" *)
  wire _1330_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13462" *)
  wire _1331_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13493" *)
  wire _1332_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13495" *)
  wire _1333_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13497" *)
  wire _1334_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13499" *)
  wire _1335_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13501" *)
  wire _1336_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13505" *)
  wire _1337_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13508" *)
  wire _1338_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13509" *)
  wire _1339_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13521" *)
  wire _1340_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13525" *)
  wire _1341_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13543" *)
  wire _1342_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13596" *)
  wire _1343_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13596" *)
  wire _1344_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13598" *)
  wire _1345_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13598" *)
  wire _1346_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13600" *)
  wire _1347_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13600" *)
  wire _1348_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13602" *)
  wire _1349_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13602" *)
  wire _1350_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13628" *)
  wire _1351_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13628" *)
  wire _1352_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13721" *)
  wire _1353_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13730" *)
  wire _1354_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13738" *)
  wire _1355_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13763" *)
  wire _1356_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13771" *)
  wire _1357_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13779" *)
  wire _1358_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13809" *)
  wire _1359_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13818" *)
  wire _1360_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13948" *)
  wire _1361_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13961" *)
  wire _1362_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14090" *)
  wire _1363_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14192" *)
  wire _1364_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14193" *)
  wire _1365_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14355" *)
  wire _1366_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14438" *)
  wire _1367_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14446" *)
  wire _1368_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14455" *)
  wire _1369_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14455" *)
  wire _1370_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14464" *)
  wire _1371_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14500" *)
  wire _1372_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14508" *)
  wire _1373_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14788" *)
  wire _1374_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14796" *)
  wire _1375_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14804" *)
  wire _1376_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14879" *)
  wire _1377_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14920" *)
  wire _1378_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14940" *)
  wire _1379_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14948" *)
  wire _1380_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14966" *)
  wire _1381_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15095" *)
  wire _1382_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15104" *)
  wire _1383_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15113" *)
  wire _1384_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15122" *)
  wire _1385_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15154" *)
  wire _1386_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15294" *)
  wire _1387_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15305" *)
  wire _1388_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15315" *)
  wire _1389_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15326" *)
  wire _1390_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15348" *)
  wire _1391_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15359" *)
  wire _1392_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15372" *)
  wire _1393_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15381" *)
  wire _1394_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15432" *)
  wire _1395_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15475" *)
  wire _1396_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15475" *)
  wire _1397_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15483" *)
  wire _1398_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15494" *)
  wire _1399_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15506" *)
  wire _1400_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15534" *)
  wire _1401_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15566" *)
  wire _1402_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15568" *)
  wire _1403_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15572" *)
  wire _1404_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15586" *)
  wire _1405_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15588" *)
  wire _1406_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15592" *)
  wire _1407_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15616" *)
  wire _1408_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15625" *)
  wire _1409_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15677" *)
  wire _1410_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15678" *)
  wire _1411_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15679" *)
  wire _1412_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15682" *)
  wire _1413_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15685" *)
  wire _1414_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15704" *)
  wire _1415_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15705" *)
  wire _1416_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15706" *)
  wire _1417_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15709" *)
  wire _1418_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15712" *)
  wire _1419_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15731" *)
  wire _1420_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15732" *)
  wire _1421_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15733" *)
  wire _1422_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15736" *)
  wire _1423_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15739" *)
  wire _1424_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15760" *)
  wire _1425_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15761" *)
  wire _1426_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15771" *)
  wire _1427_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15775" *)
  wire _1428_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15779" *)
  wire _1429_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15783" *)
  wire _1430_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15787" *)
  wire _1431_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15791" *)
  wire _1432_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15795" *)
  wire _1433_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15799" *)
  wire _1434_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15803" *)
  wire _1435_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15814" *)
  wire _1436_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15821" *)
  wire _1437_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15828" *)
  wire _1438_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15845" *)
  wire _1439_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15854" *)
  wire _1440_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15858" *)
  wire _1441_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15868" *)
  wire _1442_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15921" *)
  wire _1443_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15926" *)
  wire _1444_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15931" *)
  wire _1445_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15936" *)
  wire _1446_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15943" *)
  wire _1447_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15946" *)
  wire _1448_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15950" *)
  wire _1449_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15952" *)
  wire _1450_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15954" *)
  wire _1451_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15966" *)
  wire _1452_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15967" *)
  wire _1453_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15977" *)
  wire _1454_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15982" *)
  wire _1455_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15982" *)
  wire _1456_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15985" *)
  wire _1457_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15990" *)
  wire _1458_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15990" *)
  wire _1459_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15993" *)
  wire _1460_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15998" *)
  wire _1461_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15998" *)
  wire _1462_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16001" *)
  wire _1463_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16006" *)
  wire _1464_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16006" *)
  wire _1465_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16046" *)
  wire _1466_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16054" *)
  wire _1467_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16114" *)
  wire _1468_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16128" *)
  wire _1469_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16141" *)
  wire _1470_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16145" *)
  wire _1471_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16163" *)
  wire _1472_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16174" *)
  wire _1473_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16216" *)
  wire _1474_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16225" *)
  wire _1475_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16234" *)
  wire _1476_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16243" *)
  wire _1477_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12268" *)
  wire _1478_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12270" *)
  wire _1479_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12271" *)
  wire _1480_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12271" *)
  wire _1481_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12271" *)
  wire _1482_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12275" *)
  wire _1483_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12275" *)
  wire _1484_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12297" *)
  wire _1485_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12298" *)
  wire _1486_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12299" *)
  wire _1487_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12311" *)
  wire _1488_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12314" *)
  wire _1489_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12315" *)
  wire _1490_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12316" *)
  wire _1491_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12328" *)
  wire _1492_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12328" *)
  wire _1493_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12334" *)
  wire _1494_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12337" *)
  wire _1495_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12337" *)
  wire _1496_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12337" *)
  wire _1497_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12338" *)
  wire _1498_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12338" *)
  wire _1499_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12340" *)
  wire _1500_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12340" *)
  wire _1501_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12342" *)
  wire _1502_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12346" *)
  wire _1503_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12346" *)
  wire _1504_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12346" *)
  wire _1505_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12350" *)
  wire _1506_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12351" *)
  wire _1507_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12368" *)
  wire _1508_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12368" *)
  wire _1509_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12384" *)
  wire _1510_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12384" *)
  wire _1511_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12400" *)
  wire _1512_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12400" *)
  wire _1513_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12406" *)
  wire _1514_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12409" *)
  wire _1515_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12410" *)
  wire _1516_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12413" *)
  wire _1517_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12413" *)
  wire _1518_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12414" *)
  wire _1519_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12418" *)
  wire _1520_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12419" *)
  wire _1521_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12437" *)
  wire _1522_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12437" *)
  wire _1523_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12439" *)
  wire _1524_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12453" *)
  wire _1525_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12454" *)
  wire _1526_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12454" *)
  wire _1527_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12466" *)
  wire _1528_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12466" *)
  wire _1529_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12466" *)
  wire _1530_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12467" *)
  wire _1531_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12467" *)
  wire _1532_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12471" *)
  wire _1533_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12471" *)
  wire _1534_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12486" *)
  wire _1535_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12486" *)
  wire _1536_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12486" *)
  wire _1537_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12487" *)
  wire _1538_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12492" *)
  wire _1539_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12492" *)
  wire _1540_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12493" *)
  wire _1541_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12494" *)
  wire _1542_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12499" *)
  wire _1543_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12502" *)
  wire _1544_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12502" *)
  wire _1545_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12508" *)
  wire _1546_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12508" *)
  wire _1547_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12518" *)
  wire _1548_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12519" *)
  wire _1549_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12519" *)
  wire _1550_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12520" *)
  wire _1551_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12520" *)
  wire _1552_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12521" *)
  wire _1553_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12521" *)
  wire _1554_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12521" *)
  wire _1555_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12521" *)
  wire _1556_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12524" *)
  wire _1557_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12524" *)
  wire _1558_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12532" *)
  wire _1559_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12533" *)
  wire _1560_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12534" *)
  wire _1561_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12539" *)
  wire _1562_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12539" *)
  wire _1563_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12543" *)
  wire _1564_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12544" *)
  wire _1565_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12544" *)
  wire _1566_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12545" *)
  wire _1567_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12545" *)
  wire _1568_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12546" *)
  wire _1569_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12546" *)
  wire _1570_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12546" *)
  wire _1571_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12546" *)
  wire _1572_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12548" *)
  wire _1573_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12548" *)
  wire _1574_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12576" *)
  wire _1575_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12577" *)
  wire _1576_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12590" *)
  wire _1577_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12591" *)
  wire _1578_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12592" *)
  wire _1579_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12596" *)
  wire _1580_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12622" *)
  wire _1581_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12639" *)
  wire _1582_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12711" *)
  wire _1583_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12723" *)
  wire _1584_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12735" *)
  wire _1585_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12747" *)
  wire _1586_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12767" *)
  wire _1587_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12767" *)
  wire _1588_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12810" *)
  wire _1589_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12812" *)
  wire _1590_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12814" *)
  wire _1591_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12816" *)
  wire _1592_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12818" *)
  wire _1593_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12818" *)
  wire _1594_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12883" *)
  wire _1595_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12883" *)
  wire _1596_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12884" *)
  wire _1597_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12884" *)
  wire _1598_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12885" *)
  wire _1599_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12885" *)
  wire _1600_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12886" *)
  wire _1601_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12886" *)
  wire _1602_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12887" *)
  wire _1603_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12887" *)
  wire _1604_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12888" *)
  wire _1605_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12888" *)
  wire _1606_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12889" *)
  wire _1607_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12889" *)
  wire _1608_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12890" *)
  wire _1609_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12890" *)
  wire _1610_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12891" *)
  wire _1611_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12891" *)
  wire _1612_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12892" *)
  wire _1613_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12892" *)
  wire _1614_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12893" *)
  wire _1615_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12893" *)
  wire _1616_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12894" *)
  wire _1617_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12894" *)
  wire _1618_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12903" *)
  wire _1619_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12903" *)
  wire _1620_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12904" *)
  wire _1621_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12904" *)
  wire _1622_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12905" *)
  wire _1623_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12905" *)
  wire _1624_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12906" *)
  wire _1625_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12906" *)
  wire _1626_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12907" *)
  wire _1627_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12907" *)
  wire _1628_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12908" *)
  wire _1629_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12908" *)
  wire _1630_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12909" *)
  wire _1631_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12909" *)
  wire _1632_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12910" *)
  wire _1633_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12910" *)
  wire _1634_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12911" *)
  wire _1635_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12911" *)
  wire _1636_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12912" *)
  wire _1637_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12912" *)
  wire _1638_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12913" *)
  wire _1639_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12913" *)
  wire _1640_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12914" *)
  wire _1641_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12914" *)
  wire _1642_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12923" *)
  wire _1643_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12923" *)
  wire _1644_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12924" *)
  wire _1645_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12924" *)
  wire _1646_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12925" *)
  wire _1647_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12925" *)
  wire _1648_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12926" *)
  wire _1649_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12926" *)
  wire _1650_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12927" *)
  wire _1651_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12927" *)
  wire _1652_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12928" *)
  wire _1653_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12928" *)
  wire _1654_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12929" *)
  wire _1655_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12929" *)
  wire _1656_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12930" *)
  wire _1657_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12930" *)
  wire _1658_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12931" *)
  wire _1659_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12931" *)
  wire _1660_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12932" *)
  wire _1661_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12932" *)
  wire _1662_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12933" *)
  wire _1663_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12933" *)
  wire _1664_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12934" *)
  wire _1665_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12934" *)
  wire _1666_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12943" *)
  wire _1667_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12943" *)
  wire _1668_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12944" *)
  wire _1669_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12944" *)
  wire _1670_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12945" *)
  wire _1671_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12945" *)
  wire _1672_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12946" *)
  wire _1673_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12946" *)
  wire _1674_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12947" *)
  wire _1675_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12947" *)
  wire _1676_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12948" *)
  wire _1677_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12948" *)
  wire _1678_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12949" *)
  wire _1679_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12949" *)
  wire _1680_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12950" *)
  wire _1681_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12950" *)
  wire _1682_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12951" *)
  wire _1683_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12951" *)
  wire _1684_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12952" *)
  wire _1685_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12952" *)
  wire _1686_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12953" *)
  wire _1687_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12953" *)
  wire _1688_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12954" *)
  wire _1689_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12954" *)
  wire _1690_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12973" *)
  wire _1691_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12995" *)
  wire _1692_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12997" *)
  wire _1693_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12999" *)
  wire _1694_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13006" *)
  wire _1695_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13007" *)
  wire _1696_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13007" *)
  wire _1697_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13008" *)
  wire _1698_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13009" *)
  wire _1699_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13075" *)
  wire _1700_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13082" *)
  wire _1701_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13089" *)
  wire _1702_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13096" *)
  wire _1703_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13125" *)
  wire _1704_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13126" *)
  wire _1705_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13129" *)
  wire _1706_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13132" *)
  wire _1707_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13137" *)
  wire _1708_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13137" *)
  wire _1709_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13147" *)
  wire _1710_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13148" *)
  wire _1711_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13151" *)
  wire _1712_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13161" *)
  wire _1713_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13162" *)
  wire _1714_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13165" *)
  wire _1715_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13169" *)
  wire _1716_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13175" *)
  wire _1717_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13178" *)
  wire _1718_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13182" *)
  wire _1719_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13185" *)
  wire _1720_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13194" *)
  wire _1721_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13271" *)
  wire _1722_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13271" *)
  wire _1723_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13274" *)
  wire _1724_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13291" *)
  wire _1725_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13293" *)
  wire _1726_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13295" *)
  wire _1727_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13297" *)
  wire _1728_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13300" *)
  wire _1729_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13302" *)
  wire _1730_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13304" *)
  wire _1731_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13304" *)
  wire _1732_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13305" *)
  wire _1733_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13312" *)
  wire _1734_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13312" *)
  wire _1735_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13313" *)
  wire _1736_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13314" *)
  wire _1737_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13314" *)
  wire _1738_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13314" *)
  wire _1739_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13316" *)
  wire _1740_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13317" *)
  wire _1741_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13317" *)
  wire _1742_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13322" *)
  wire _1743_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13324" *)
  wire _1744_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13324" *)
  wire _1745_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13324" *)
  wire _1746_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13325" *)
  wire _1747_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13326" *)
  wire _1748_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13328" *)
  wire _1749_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13330" *)
  wire _1750_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13330" *)
  wire _1751_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13330" *)
  wire _1752_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13331" *)
  wire _1753_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13331" *)
  wire _1754_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13333" *)
  wire _1755_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13335" *)
  wire _1756_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13341" *)
  wire _1757_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13344" *)
  wire _1758_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13347" *)
  wire _1759_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13354" *)
  wire _1760_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13365" *)
  wire _1761_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13371" *)
  wire _1762_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13371" *)
  wire _1763_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13377" *)
  wire _1764_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13380" *)
  wire _1765_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13388" *)
  wire _1766_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13391" *)
  wire _1767_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13394" *)
  wire _1768_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13396" *)
  wire _1769_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13403" *)
  wire _1770_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13414" *)
  wire _1771_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13425" *)
  wire _1772_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13427" *)
  wire _1773_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13429" *)
  wire _1774_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13436" *)
  wire _1775_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13436" *)
  wire _1776_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13436" *)
  wire _1777_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13439" *)
  wire _1778_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13449" *)
  wire _1779_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13456" *)
  wire _1780_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13484" *)
  wire _1781_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13485" *)
  wire _1782_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13485" *)
  wire _1783_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13487" *)
  wire _1784_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13488" *)
  wire _1785_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13490" *)
  wire _1786_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13490" *)
  wire _1787_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13491" *)
  wire _1788_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13491" *)
  wire _1789_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13491" *)
  wire _1790_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13492" *)
  wire _1791_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13493" *)
  wire _1792_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13493" *)
  wire _1793_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13494" *)
  wire _1794_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13512" *)
  wire _1795_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13512" *)
  wire _1796_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13516" *)
  wire _1797_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13543" *)
  wire _1798_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13548" *)
  wire _1799_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13596" *)
  wire _1800_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13598" *)
  wire _1801_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13600" *)
  wire _1802_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13602" *)
  wire _1803_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13720" *)
  wire _1804_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13729" *)
  wire _1805_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13729" *)
  wire _1806_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13737" *)
  wire _1807_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13788" *)
  wire _1808_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13799" *)
  wire _1809_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13799" *)
  wire _1810_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13809" *)
  wire _1811_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13809" *)
  wire _1812_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13817" *)
  wire _1813_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13960" *)
  wire _1814_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14088" *)
  wire _1815_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14184" *)
  wire _1816_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14192" *)
  wire _1817_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14194" *)
  wire _1818_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14261" *)
  wire _1819_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14269" *)
  wire _1820_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14271" *)
  wire _1821_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14280" *)
  wire _1822_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14288" *)
  wire _1823_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14290" *)
  wire _1824_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14299" *)
  wire _1825_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14307" *)
  wire _1826_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14309" *)
  wire _1827_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14345" *)
  wire _1828_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14346" *)
  wire _1829_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14364" *)
  wire _1830_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14383" *)
  wire _1831_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14403" *)
  wire _1832_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14421" *)
  wire _1833_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14454" *)
  wire _1834_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14455" *)
  wire _1835_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14455" *)
  wire _1836_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14455" *)
  wire _1837_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14483" *)
  wire _1838_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14796" *)
  wire _1839_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14804" *)
  wire _1840_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14804" *)
  wire _1841_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14821" *)
  wire _1842_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14821" *)
  wire _1843_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14832" *)
  wire _1844_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14832" *)
  wire _1845_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14843" *)
  wire _1846_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14843" *)
  wire _1847_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14854" *)
  wire _1848_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14854" *)
  wire _1849_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15094" *)
  wire _1850_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15095" *)
  wire _1851_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15095" *)
  wire _1852_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15104" *)
  wire _1853_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15113" *)
  wire _1854_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15122" *)
  wire _1855_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15163" *)
  wire _1856_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15173" *)
  wire _1857_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15183" *)
  wire _1858_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15193" *)
  wire _1859_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15305" *)
  wire _1860_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15326" *)
  wire _1861_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15338" *)
  wire _1862_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15372" *)
  wire _1863_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15381" *)
  wire _1864_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15473" *)
  wire _1865_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15474" *)
  wire _1866_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15474" *)
  wire _1867_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15474" *)
  wire _1868_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15475" *)
  wire _1869_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15475" *)
  wire _1870_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15534" *)
  wire _1871_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15566" *)
  wire _1872_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15582" *)
  wire _1873_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15586" *)
  wire _1874_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15602" *)
  wire _1875_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15625" *)
  wire _1876_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15626" *)
  wire _1877_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15627" *)
  wire _1878_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15628" *)
  wire _1879_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15628" *)
  wire _1880_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15630" *)
  wire _1881_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15630" *)
  wire _1882_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15630" *)
  wire _1883_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15633" *)
  wire _1884_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15633" *)
  wire _1885_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15635" *)
  wire _1886_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15636" *)
  wire _1887_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15636" *)
  wire _1888_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15638" *)
  wire _1889_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15638" *)
  wire _1890_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15638" *)
  wire _1891_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15641" *)
  wire _1892_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15643" *)
  wire _1893_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15644" *)
  wire _1894_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15644" *)
  wire _1895_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15646" *)
  wire _1896_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15646" *)
  wire _1897_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15646" *)
  wire _1898_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15649" *)
  wire _1899_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15651" *)
  wire _1900_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15652" *)
  wire _1901_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15652" *)
  wire _1902_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15654" *)
  wire _1903_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15654" *)
  wire _1904_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15654" *)
  wire _1905_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15657" *)
  wire _1906_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15660" *)
  wire _1907_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15660" *)
  wire _1908_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15663" *)
  wire _1909_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15664" *)
  wire _1910_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15664" *)
  wire _1911_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15664" *)
  wire _1912_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15665" *)
  wire _1913_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15665" *)
  wire _1914_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15667" *)
  wire _1915_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15667" *)
  wire _1916_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15667" *)
  wire _1917_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15668" *)
  wire _1918_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15668" *)
  wire _1919_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15668" *)
  wire _1920_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15670" *)
  wire _1921_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15673" *)
  wire _1922_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15673" *)
  wire _1923_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15674" *)
  wire _1924_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15674" *)
  wire _1925_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15677" *)
  wire _1926_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15677" *)
  wire _1927_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15680" *)
  wire _1928_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15680" *)
  wire _1929_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15680" *)
  wire _1930_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15681" *)
  wire _1931_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15681" *)
  wire _1932_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15681" *)
  wire _1933_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15682" *)
  wire _1934_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15682" *)
  wire _1935_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15682" *)
  wire _1936_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15684" *)
  wire _1937_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15684" *)
  wire _1938_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15684" *)
  wire _1939_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15685" *)
  wire _1940_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15685" *)
  wire _1941_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15685" *)
  wire _1942_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15686" *)
  wire _1943_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15688" *)
  wire _1944_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15690" *)
  wire _1945_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15691" *)
  wire _1946_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15691" *)
  wire _1947_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15691" *)
  wire _1948_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15692" *)
  wire _1949_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15692" *)
  wire _1950_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15694" *)
  wire _1951_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15694" *)
  wire _1952_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15694" *)
  wire _1953_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15695" *)
  wire _1954_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15695" *)
  wire _1955_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15695" *)
  wire _1956_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15697" *)
  wire _1957_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15701" *)
  wire _1958_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15701" *)
  wire _1959_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15704" *)
  wire _1960_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15704" *)
  wire _1961_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15707" *)
  wire _1962_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15707" *)
  wire _1963_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15707" *)
  wire _1964_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15708" *)
  wire _1965_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15708" *)
  wire _1966_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15708" *)
  wire _1967_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15709" *)
  wire _1968_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15709" *)
  wire _1969_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15709" *)
  wire _1970_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15711" *)
  wire _1971_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15711" *)
  wire _1972_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15711" *)
  wire _1973_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15712" *)
  wire _1974_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15712" *)
  wire _1975_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15712" *)
  wire _1976_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15713" *)
  wire _1977_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15715" *)
  wire _1978_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15717" *)
  wire _1979_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15718" *)
  wire _1980_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15718" *)
  wire _1981_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15718" *)
  wire _1982_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15719" *)
  wire _1983_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15719" *)
  wire _1984_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15721" *)
  wire _1985_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15721" *)
  wire _1986_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15721" *)
  wire _1987_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15722" *)
  wire _1988_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15722" *)
  wire _1989_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15722" *)
  wire _1990_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15724" *)
  wire _1991_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15728" *)
  wire _1992_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15728" *)
  wire _1993_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15731" *)
  wire _1994_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15731" *)
  wire _1995_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15734" *)
  wire _1996_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15734" *)
  wire _1997_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15734" *)
  wire _1998_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15735" *)
  wire _1999_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15735" *)
  wire _2000_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15735" *)
  wire _2001_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15736" *)
  wire _2002_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15736" *)
  wire _2003_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15736" *)
  wire _2004_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15738" *)
  wire _2005_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15738" *)
  wire _2006_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15738" *)
  wire _2007_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15739" *)
  wire _2008_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15739" *)
  wire _2009_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15739" *)
  wire _2010_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15740" *)
  wire _2011_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15742" *)
  wire _2012_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15744" *)
  wire _2013_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15745" *)
  wire _2014_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15745" *)
  wire _2015_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15745" *)
  wire _2016_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15746" *)
  wire _2017_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15746" *)
  wire _2018_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15746" *)
  wire _2019_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15747" *)
  wire _2020_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15747" *)
  wire _2021_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15749" *)
  wire _2022_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15749" *)
  wire _2023_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15749" *)
  wire _2024_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15750" *)
  wire _2025_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15750" *)
  wire _2026_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15751" *)
  wire _2027_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15751" *)
  wire _2028_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15751" *)
  wire _2029_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15751" *)
  wire _2030_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15753" *)
  wire _2031_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15756" *)
  wire _2032_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15757" *)
  wire _2033_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15757" *)
  wire _2034_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15757" *)
  wire _2035_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15758" *)
  wire _2036_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15758" *)
  wire _2037_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15762" *)
  wire _2038_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15762" *)
  wire _2039_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15762" *)
  wire _2040_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15766" *)
  wire _2041_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15766" *)
  wire _2042_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15767" *)
  wire _2043_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15767" *)
  wire _2044_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15767" *)
  wire _2045_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15770" *)
  wire _2046_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15770" *)
  wire _2047_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15770" *)
  wire _2048_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15772" *)
  wire _2049_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15772" *)
  wire _2050_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15772" *)
  wire _2051_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15775" *)
  wire _2052_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15775" *)
  wire _2053_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15778" *)
  wire _2054_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15778" *)
  wire _2055_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15778" *)
  wire _2056_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15780" *)
  wire _2057_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15780" *)
  wire _2058_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15780" *)
  wire _2059_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15783" *)
  wire _2060_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15786" *)
  wire _2061_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15786" *)
  wire _2062_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15786" *)
  wire _2063_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15788" *)
  wire _2064_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15788" *)
  wire _2065_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15788" *)
  wire _2066_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15791" *)
  wire _2067_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15794" *)
  wire _2068_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15794" *)
  wire _2069_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15794" *)
  wire _2070_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15796" *)
  wire _2071_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15796" *)
  wire _2072_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15796" *)
  wire _2073_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15799" *)
  wire _2074_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15802" *)
  wire _2075_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15803" *)
  wire _2076_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15804" *)
  wire _2077_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15807" *)
  wire _2078_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15807" *)
  wire _2079_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15807" *)
  wire _2080_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15811" *)
  wire _2081_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15811" *)
  wire _2082_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15811" *)
  wire _2083_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15811" *)
  wire _2084_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15814" *)
  wire _2085_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15814" *)
  wire _2086_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15818" *)
  wire _2087_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15818" *)
  wire _2088_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15821" *)
  wire _2089_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15821" *)
  wire _2090_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15825" *)
  wire _2091_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15825" *)
  wire _2092_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15828" *)
  wire _2093_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15828" *)
  wire _2094_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15831" *)
  wire _2095_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15831" *)
  wire _2096_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15831" *)
  wire _2097_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15834" *)
  wire _2098_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15835" *)
  wire _2099_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15835" *)
  wire _2100_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15837" *)
  wire _2101_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15838" *)
  wire _2102_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15838" *)
  wire _2103_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15841" *)
  wire _2104_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15842" *)
  wire _2105_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15842" *)
  wire _2106_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15842" *)
  wire _2107_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15846" *)
  wire _2108_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15846" *)
  wire _2109_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15846" *)
  wire _2110_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15847" *)
  wire _2111_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15847" *)
  wire _2112_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15851" *)
  wire _2113_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15851" *)
  wire _2114_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15854" *)
  wire _2115_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15854" *)
  wire _2116_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15861" *)
  wire _2117_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15862" *)
  wire _2118_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15862" *)
  wire _2119_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15862" *)
  wire _2120_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15880" *)
  wire _2121_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15880" *)
  wire _2122_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15880" *)
  wire _2123_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15881" *)
  wire _2124_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15881" *)
  wire _2125_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15881" *)
  wire _2126_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15882" *)
  wire _2127_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15886" *)
  wire _2128_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15887" *)
  wire _2129_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15887" *)
  wire _2130_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15887" *)
  wire _2131_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15890" *)
  wire _2132_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15890" *)
  wire _2133_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15890" *)
  wire _2134_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15891" *)
  wire _2135_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15891" *)
  wire _2136_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15891" *)
  wire _2137_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15892" *)
  wire _2138_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15896" *)
  wire _2139_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15897" *)
  wire _2140_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15897" *)
  wire _2141_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15897" *)
  wire _2142_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15900" *)
  wire _2143_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15900" *)
  wire _2144_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15900" *)
  wire _2145_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15901" *)
  wire _2146_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15901" *)
  wire _2147_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15901" *)
  wire _2148_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15902" *)
  wire _2149_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15906" *)
  wire _2150_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15907" *)
  wire _2151_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15907" *)
  wire _2152_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15907" *)
  wire _2153_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15910" *)
  wire _2154_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15910" *)
  wire _2155_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15910" *)
  wire _2156_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15911" *)
  wire _2157_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15911" *)
  wire _2158_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15911" *)
  wire _2159_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15912" *)
  wire _2160_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15916" *)
  wire _2161_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15917" *)
  wire _2162_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15917" *)
  wire _2163_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15917" *)
  wire _2164_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15919" *)
  wire _2165_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15920" *)
  wire _2166_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15920" *)
  wire _2167_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15921" *)
  wire _2168_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15922" *)
  wire _2169_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15924" *)
  wire _2170_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15925" *)
  wire _2171_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15925" *)
  wire _2172_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15926" *)
  wire _2173_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15927" *)
  wire _2174_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15929" *)
  wire _2175_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15930" *)
  wire _2176_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15930" *)
  wire _2177_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15931" *)
  wire _2178_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15932" *)
  wire _2179_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15934" *)
  wire _2180_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15935" *)
  wire _2181_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15935" *)
  wire _2182_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15936" *)
  wire _2183_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15937" *)
  wire _2184_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15959" *)
  wire _2185_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15962" *)
  wire _2186_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15962" *)
  wire _2187_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15963" *)
  wire _2188_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15963" *)
  wire _2189_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15963" *)
  wire _2190_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15964" *)
  wire _2191_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15966" *)
  wire _2192_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15967" *)
  wire _2193_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15967" *)
  wire _2194_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15971" *)
  wire _2195_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15971" *)
  wire _2196_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15972" *)
  wire _2197_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15972" *)
  wire _2198_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15974" *)
  wire _2199_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15974" *)
  wire _2200_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15977" *)
  wire _2201_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15977" *)
  wire _2202_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15977" *)
  wire _2203_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15978" *)
  wire _2204_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15978" *)
  wire _2205_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15978" *)
  wire _2206_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15981" *)
  wire _2207_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15982" *)
  wire _2208_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15982" *)
  wire _2209_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15982" *)
  wire _2210_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15982" *)
  wire _2211_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15982" *)
  wire _2212_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15985" *)
  wire _2213_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15986" *)
  wire _2214_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15986" *)
  wire _2215_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15986" *)
  wire _2216_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15990" *)
  wire _2217_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15990" *)
  wire _2218_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15990" *)
  wire _2219_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15990" *)
  wire _2220_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15993" *)
  wire _2221_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15994" *)
  wire _2222_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15994" *)
  wire _2223_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15994" *)
  wire _2224_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15998" *)
  wire _2225_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15998" *)
  wire _2226_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15998" *)
  wire _2227_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15998" *)
  wire _2228_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16001" *)
  wire _2229_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16002" *)
  wire _2230_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16002" *)
  wire _2231_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16002" *)
  wire _2232_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16006" *)
  wire _2233_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16006" *)
  wire _2234_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16006" *)
  wire _2235_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16006" *)
  wire _2236_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16011" *)
  wire _2237_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16012" *)
  wire _2238_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16012" *)
  wire _2239_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16013" *)
  wire _2240_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16013" *)
  wire _2241_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16013" *)
  wire _2242_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16015" *)
  wire _2243_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16016" *)
  wire _2244_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16016" *)
  wire _2245_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16017" *)
  wire _2246_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16017" *)
  wire _2247_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16017" *)
  wire _2248_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16020" *)
  wire _2249_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16021" *)
  wire _2250_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16021" *)
  wire _2251_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16022" *)
  wire _2252_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16022" *)
  wire _2253_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16022" *)
  wire _2254_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16024" *)
  wire _2255_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16025" *)
  wire _2256_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16025" *)
  wire _2257_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16026" *)
  wire _2258_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16026" *)
  wire _2259_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16026" *)
  wire _2260_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16029" *)
  wire _2261_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16030" *)
  wire _2262_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16030" *)
  wire _2263_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16031" *)
  wire _2264_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16031" *)
  wire _2265_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16031" *)
  wire _2266_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16033" *)
  wire _2267_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16034" *)
  wire _2268_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16034" *)
  wire _2269_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16035" *)
  wire _2270_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16035" *)
  wire _2271_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16035" *)
  wire _2272_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16038" *)
  wire _2273_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16039" *)
  wire _2274_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16039" *)
  wire _2275_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16039" *)
  wire _2276_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16040" *)
  wire _2277_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16040" *)
  wire _2278_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16042" *)
  wire _2279_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16043" *)
  wire _2280_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16043" *)
  wire _2281_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16043" *)
  wire _2282_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16044" *)
  wire _2283_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16044" *)
  wire _2284_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16063" *)
  wire _2285_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16066" *)
  wire _2286_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16089" *)
  wire _2287_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16092" *)
  wire _2288_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16093" *)
  wire _2289_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16094" *)
  wire _2290_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16094" *)
  wire _2291_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16095" *)
  wire _2292_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16095" *)
  wire _2293_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16099" *)
  wire _2294_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16100" *)
  wire _2295_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16100" *)
  wire _2296_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16101" *)
  wire _2297_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16101" *)
  wire _2298_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16101" *)
  wire _2299_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16115" *)
  wire _2300_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16118" *)
  wire _2301_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16129" *)
  wire _2302_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16132" *)
  wire _2303_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16145" *)
  wire _2304_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16145" *)
  wire _2305_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16146" *)
  wire _2306_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16157" *)
  wire _2307_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16168" *)
  wire _2308_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16265" *)
  wire _2309_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16265" *)
  wire _2310_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16265" *)
  wire _2311_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16265" *)
  wire _2312_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16265" *)
  wire _2313_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16265" *)
  wire _2314_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16265" *)
  wire _2315_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16265" *)
  wire _2316_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16265" *)
  wire _2317_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16265" *)
  wire _2318_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16265" *)
  wire _2319_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16266" *)
  wire _2320_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16266" *)
  wire _2321_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16266" *)
  wire _2322_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16266" *)
  wire _2323_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16266" *)
  wire _2324_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16266" *)
  wire _2325_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16266" *)
  wire _2326_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16266" *)
  wire _2327_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16266" *)
  wire _2328_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16266" *)
  wire _2329_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16266" *)
  wire _2330_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16279" *)
  wire _2331_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16279" *)
  wire _2332_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16279" *)
  wire _2333_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16279" *)
  wire _2334_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16279" *)
  wire _2335_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16279" *)
  wire _2336_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16279" *)
  wire _2337_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16279" *)
  wire _2338_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16279" *)
  wire _2339_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16279" *)
  wire _2340_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16280" *)
  wire _2341_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16280" *)
  wire _2342_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16280" *)
  wire _2343_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16280" *)
  wire _2344_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16280" *)
  wire _2345_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16280" *)
  wire _2346_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16280" *)
  wire _2347_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16280" *)
  wire _2348_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16280" *)
  wire _2349_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16280" *)
  wire _2350_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16281" *)
  wire _2351_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16281" *)
  wire _2352_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16281" *)
  wire _2353_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16281" *)
  wire _2354_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16281" *)
  wire _2355_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16281" *)
  wire _2356_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16295" *)
  wire _2357_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16295" *)
  wire _2358_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16296" *)
  wire _2359_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16296" *)
  wire _2360_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16297" *)
  wire _2361_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16297" *)
  wire _2362_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16314" *)
  wire _2363_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16314" *)
  wire _2364_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16315" *)
  wire _2365_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16315" *)
  wire _2366_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16316" *)
  wire _2367_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16316" *)
  wire _2368_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16317" *)
  wire _2369_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16317" *)
  wire _2370_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16318" *)
  wire _2371_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16318" *)
  wire _2372_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16319" *)
  wire _2373_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16319" *)
  wire _2374_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16331" *)
  wire [21:0] _2375_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16331" *)
  wire [21:0] _2376_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16331" *)
  wire [21:0] _2377_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16331" *)
  wire [21:0] _2378_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16331" *)
  wire [21:0] _2379_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16332" *)
  wire [21:0] _2380_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16332" *)
  wire [21:0] _2381_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16332" *)
  wire [21:0] _2382_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16345" *)
  wire [21:0] _2383_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16346" *)
  wire [21:0] _2384_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16359" *)
  wire [30:0] _2385_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16359" *)
  wire [30:0] _2386_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16359" *)
  wire [30:0] _2387_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16359" *)
  wire [30:0] _2388_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16372" *)
  wire [7:0] _2389_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16372" *)
  wire [7:0] _2390_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16372" *)
  wire [7:0] _2391_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16372" *)
  wire [7:0] _2392_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16372" *)
  wire [7:0] _2393_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16372" *)
  wire [7:0] _2394_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16372" *)
  wire [7:0] _2395_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16372" *)
  wire [7:0] _2396_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16372" *)
  wire [7:0] _2397_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16372" *)
  wire [7:0] _2398_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16372" *)
  wire [7:0] _2399_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16372" *)
  wire [7:0] _2400_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16372" *)
  wire [7:0] _2401_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16372" *)
  wire [7:0] _2402_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16372" *)
  wire [7:0] _2403_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16372" *)
  wire [7:0] _2404_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16373" *)
  wire [7:0] _2405_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16373" *)
  wire [7:0] _2406_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16373" *)
  wire [7:0] _2407_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16373" *)
  wire [7:0] _2408_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16373" *)
  wire [7:0] _2409_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16373" *)
  wire [7:0] _2410_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16373" *)
  wire [7:0] _2411_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16373" *)
  wire [7:0] _2412_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16373" *)
  wire [7:0] _2413_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16373" *)
  wire [7:0] _2414_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16373" *)
  wire [7:0] _2415_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16388" *)
  wire [7:0] _2416_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16388" *)
  wire [7:0] _2417_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16389" *)
  wire [7:0] _2418_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16389" *)
  wire [7:0] _2419_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16390" *)
  wire [7:0] _2420_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16390" *)
  wire [7:0] _2421_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16391" *)
  wire [7:0] _2422_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16391" *)
  wire [7:0] _2423_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16408" *)
  wire [7:0] _2424_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16409" *)
  wire [7:0] _2425_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16410" *)
  wire [7:0] _2426_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16411" *)
  wire [7:0] _2427_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16412" *)
  wire [7:0] _2428_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16430" *)
  wire [7:0] _2429_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16431" *)
  wire [7:0] _2430_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16432" *)
  wire [7:0] _2431_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16433" *)
  wire [7:0] _2432_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16434" *)
  wire [7:0] _2433_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16435" *)
  wire [7:0] _2434_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12657" *)
  wire _2435_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12667" *)
  wire _2436_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12678" *)
  wire _2437_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12689" *)
  wire _2438_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11074" *)
  wire AluIn_data_and_1_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11108" *)
  wire AluIn_data_and_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10890" *)
  wire [30:0] AluIn_data_mux1h_11_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10893" *)
  wire [30:0] AluIn_data_mux1h_13_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10884" *)
  wire [30:0] AluIn_data_mux1h_7_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10887" *)
  wire [30:0] AluIn_data_mux1h_9_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10593" *)
  reg [127:0] AluIn_data_sva_127;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10594" *)
  reg [127:0] AluIn_data_sva_128;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10768" *)
  reg [30:0] AluIn_data_sva_3_126_96_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10771" *)
  reg [30:0] AluIn_data_sva_3_30_0_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10770" *)
  reg [30:0] AluIn_data_sva_3_62_32_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10769" *)
  reg [30:0] AluIn_data_sva_3_94_64_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10589" *)
  reg AluOut_data_0_0_sva_10;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10590" *)
  reg AluOut_data_0_0_sva_11;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10588" *)
  reg AluOut_data_0_0_sva_9;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10585" *)
  reg AluOut_data_1_0_sva_10;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10586" *)
  reg AluOut_data_1_0_sva_11;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10587" *)
  reg AluOut_data_1_0_sva_12;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10507" *)
  reg AluOut_data_2_0_lpi_1_dfm_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10583" *)
  reg AluOut_data_2_0_sva_10;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10584" *)
  reg AluOut_data_2_0_sva_11;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10983" *)
  wire AluOut_data_2_0_sva_3_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10582" *)
  reg AluOut_data_2_0_sva_9;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10506" *)
  reg [21:0] AluOut_data_2_22_1_lpi_1_dfm_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10938" *)
  wire [21:0] AluOut_data_2_22_1_lpi_1_dfm_3_mx1w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10505" *)
  reg [7:0] AluOut_data_2_30_23_lpi_1_dfm_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10939" *)
  wire [7:0] AluOut_data_2_30_23_lpi_1_dfm_3_mx1w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10621" *)
  reg AluOut_data_2_31_lpi_1_dfm_6;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10622" *)
  reg AluOut_data_2_31_lpi_1_dfm_7;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11119" *)
  wire AluOut_data_and_12_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11098" *)
  wire AluOut_data_and_15_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11101" *)
  wire AluOut_data_and_17_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11560" *)
  wire AluOut_data_and_3_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10825" *)
  wire AluOut_data_and_5_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11554" *)
  wire AluOut_data_and_7_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11087" *)
  wire AluOut_data_and_8_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11550" *)
  wire AluOut_data_or_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11552" *)
  wire AluOut_data_or_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11558" *)
  wire AluOut_data_or_3_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11556" *)
  wire AluOut_data_or_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10782" *)
  wire FpAdd_8U_23U_FpAdd_8U_23U_nor_11_m1c;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10781" *)
  wire FpAdd_8U_23U_FpAdd_8U_23U_nor_5_m1c;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10780" *)
  wire FpAdd_8U_23U_FpAdd_8U_23U_nor_7_m1c;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10779" *)
  wire FpAdd_8U_23U_FpAdd_8U_23U_nor_9_m1c;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11321" *)
  wire [22:0] FpAdd_8U_23U_FpAdd_8U_23U_or_4_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11342" *)
  wire [22:0] FpAdd_8U_23U_FpAdd_8U_23U_or_5_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11351" *)
  wire [22:0] FpAdd_8U_23U_FpAdd_8U_23U_or_6_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11360" *)
  wire [22:0] FpAdd_8U_23U_FpAdd_8U_23U_or_7_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11010" *)
  wire [48:0] FpAdd_8U_23U_a_int_mant_p1_1_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11009" *)
  wire [48:0] FpAdd_8U_23U_a_int_mant_p1_2_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11008" *)
  wire [48:0] FpAdd_8U_23U_a_int_mant_p1_3_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11007" *)
  wire [48:0] FpAdd_8U_23U_a_int_mant_p1_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10920" *)
  wire FpAdd_8U_23U_a_right_shift_qelse_and_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10922" *)
  wire FpAdd_8U_23U_a_right_shift_qelse_and_tmp_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10924" *)
  wire FpAdd_8U_23U_a_right_shift_qelse_and_tmp_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10926" *)
  wire FpAdd_8U_23U_a_right_shift_qelse_and_tmp_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10485" *)
  reg [7:0] FpAdd_8U_23U_a_right_shift_qr_1_lpi_1_dfm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10601" *)
  reg [7:0] FpAdd_8U_23U_a_right_shift_qr_1_lpi_1_dfm_5;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10960" *)
  wire [7:0] FpAdd_8U_23U_a_right_shift_qr_1_lpi_1_dfm_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10489" *)
  reg [7:0] FpAdd_8U_23U_a_right_shift_qr_2_lpi_1_dfm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10606" *)
  reg [7:0] FpAdd_8U_23U_a_right_shift_qr_2_lpi_1_dfm_5;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10956" *)
  wire [7:0] FpAdd_8U_23U_a_right_shift_qr_2_lpi_1_dfm_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10493" *)
  reg [7:0] FpAdd_8U_23U_a_right_shift_qr_3_lpi_1_dfm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10611" *)
  reg [7:0] FpAdd_8U_23U_a_right_shift_qr_3_lpi_1_dfm_5;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10952" *)
  wire [7:0] FpAdd_8U_23U_a_right_shift_qr_3_lpi_1_dfm_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10497" *)
  reg [7:0] FpAdd_8U_23U_a_right_shift_qr_lpi_1_dfm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10616" *)
  reg [7:0] FpAdd_8U_23U_a_right_shift_qr_lpi_1_dfm_5;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10948" *)
  wire [7:0] FpAdd_8U_23U_a_right_shift_qr_lpi_1_dfm_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10998" *)
  wire [48:0] FpAdd_8U_23U_addend_larger_asn_13_mx0w1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10995" *)
  wire [48:0] FpAdd_8U_23U_addend_larger_asn_19_mx0w1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11004" *)
  wire [48:0] FpAdd_8U_23U_addend_larger_asn_1_mx0w1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11001" *)
  wire [48:0] FpAdd_8U_23U_addend_larger_asn_7_mx0w1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10996" *)
  wire [48:0] FpAdd_8U_23U_addend_larger_qr_1_lpi_1_dfm_mx0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10999" *)
  wire [48:0] FpAdd_8U_23U_addend_larger_qr_2_lpi_1_dfm_mx0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11002" *)
  wire [48:0] FpAdd_8U_23U_addend_larger_qr_3_lpi_1_dfm_mx0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11005" *)
  wire [48:0] FpAdd_8U_23U_addend_larger_qr_lpi_1_dfm_mx0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10997" *)
  wire [48:0] FpAdd_8U_23U_addend_smaller_qr_1_lpi_1_dfm_mx0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11000" *)
  wire [48:0] FpAdd_8U_23U_addend_smaller_qr_2_lpi_1_dfm_mx0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11003" *)
  wire [48:0] FpAdd_8U_23U_addend_smaller_qr_3_lpi_1_dfm_mx0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11006" *)
  wire [48:0] FpAdd_8U_23U_addend_smaller_qr_lpi_1_dfm_mx0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11132" *)
  wire FpAdd_8U_23U_and_10_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11196" *)
  wire FpAdd_8U_23U_and_13_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11198" *)
  wire FpAdd_8U_23U_and_15_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11133" *)
  wire FpAdd_8U_23U_and_16_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11659" *)
  wire FpAdd_8U_23U_and_19_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10516" *)
  reg FpAdd_8U_23U_and_1_tmp_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11661" *)
  wire FpAdd_8U_23U_and_21_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11134" *)
  wire FpAdd_8U_23U_and_22_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11719" *)
  wire FpAdd_8U_23U_and_25_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11721" *)
  wire FpAdd_8U_23U_and_27_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11182" *)
  wire FpAdd_8U_23U_and_28_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11195" *)
  wire FpAdd_8U_23U_and_29_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10513" *)
  reg FpAdd_8U_23U_and_2_tmp_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11197" *)
  wire FpAdd_8U_23U_and_30_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11658" *)
  wire FpAdd_8U_23U_and_31_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11660" *)
  wire FpAdd_8U_23U_and_32_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11718" *)
  wire FpAdd_8U_23U_and_33_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11720" *)
  wire FpAdd_8U_23U_and_34_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11075" *)
  wire FpAdd_8U_23U_and_39_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10522" *)
  reg FpAdd_8U_23U_and_3_tmp_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11131" *)
  wire FpAdd_8U_23U_and_4_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11181" *)
  wire FpAdd_8U_23U_and_6_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11183" *)
  wire FpAdd_8U_23U_and_9_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11180" *)
  wire FpAdd_8U_23U_and_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10519" *)
  reg FpAdd_8U_23U_and_tmp_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11895" *)
  wire [7:0] FpAdd_8U_23U_b_right_shift_qif_mux_15_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11896" *)
  wire [7:0] FpAdd_8U_23U_b_right_shift_qif_mux_16_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11899" *)
  wire [7:0] FpAdd_8U_23U_b_right_shift_qif_mux_17_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11900" *)
  wire [7:0] FpAdd_8U_23U_b_right_shift_qif_mux_18_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11903" *)
  wire [7:0] FpAdd_8U_23U_b_right_shift_qif_mux_19_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11904" *)
  wire [7:0] FpAdd_8U_23U_b_right_shift_qif_mux_20_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11907" *)
  wire [7:0] FpAdd_8U_23U_b_right_shift_qif_mux_21_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11908" *)
  wire [7:0] FpAdd_8U_23U_b_right_shift_qif_mux_22_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10486" *)
  reg [7:0] FpAdd_8U_23U_b_right_shift_qr_1_lpi_1_dfm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10602" *)
  reg [7:0] FpAdd_8U_23U_b_right_shift_qr_1_lpi_1_dfm_5;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10959" *)
  wire [7:0] FpAdd_8U_23U_b_right_shift_qr_1_lpi_1_dfm_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10490" *)
  reg [7:0] FpAdd_8U_23U_b_right_shift_qr_2_lpi_1_dfm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10607" *)
  reg [7:0] FpAdd_8U_23U_b_right_shift_qr_2_lpi_1_dfm_5;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10955" *)
  wire [7:0] FpAdd_8U_23U_b_right_shift_qr_2_lpi_1_dfm_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10494" *)
  reg [7:0] FpAdd_8U_23U_b_right_shift_qr_3_lpi_1_dfm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10612" *)
  reg [7:0] FpAdd_8U_23U_b_right_shift_qr_3_lpi_1_dfm_5;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10951" *)
  wire [7:0] FpAdd_8U_23U_b_right_shift_qr_3_lpi_1_dfm_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10498" *)
  reg [7:0] FpAdd_8U_23U_b_right_shift_qr_lpi_1_dfm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10617" *)
  reg [7:0] FpAdd_8U_23U_b_right_shift_qr_lpi_1_dfm_5;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10947" *)
  wire [7:0] FpAdd_8U_23U_b_right_shift_qr_lpi_1_dfm_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11915" *)
  wire [48:0] FpAdd_8U_23U_else_2_mux_10_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11916" *)
  wire [48:0] FpAdd_8U_23U_else_2_mux_11_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11919" *)
  wire [48:0] FpAdd_8U_23U_else_2_mux_12_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11920" *)
  wire [48:0] FpAdd_8U_23U_else_2_mux_13_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11923" *)
  wire [48:0] FpAdd_8U_23U_else_2_mux_14_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11924" *)
  wire [48:0] FpAdd_8U_23U_else_2_mux_15_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11911" *)
  wire [48:0] FpAdd_8U_23U_else_2_mux_8_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11912" *)
  wire [48:0] FpAdd_8U_23U_else_2_mux_9_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10928" *)
  wire FpAdd_8U_23U_if_2_and_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10930" *)
  wire FpAdd_8U_23U_if_2_and_tmp_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10932" *)
  wire FpAdd_8U_23U_if_2_and_tmp_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10934" *)
  wire FpAdd_8U_23U_if_2_and_tmp_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10818" *)
  wire FpAdd_8U_23U_if_3_and_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10916" *)
  wire FpAdd_8U_23U_if_3_if_and_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10917" *)
  wire FpAdd_8U_23U_if_3_if_and_tmp_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10918" *)
  wire FpAdd_8U_23U_if_3_if_and_tmp_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10919" *)
  wire FpAdd_8U_23U_if_3_if_and_tmp_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11012" *)
  wire [48:0] FpAdd_8U_23U_int_mant_1_lpi_1_dfm_2_mx0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11018" *)
  wire [48:0] FpAdd_8U_23U_int_mant_2_lpi_1_dfm_2_mx0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11016" *)
  wire [48:0] FpAdd_8U_23U_int_mant_3_lpi_1_dfm_2_mx0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11014" *)
  wire [48:0] FpAdd_8U_23U_int_mant_4_lpi_1_dfm_2_mx0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10487" *)
  reg [49:0] FpAdd_8U_23U_int_mant_p1_1_lpi_1_dfm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10603" *)
  reg [49:0] FpAdd_8U_23U_int_mant_p1_1_lpi_1_dfm_5;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10491" *)
  reg [49:0] FpAdd_8U_23U_int_mant_p1_2_lpi_1_dfm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10608" *)
  reg [49:0] FpAdd_8U_23U_int_mant_p1_2_lpi_1_dfm_5;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10495" *)
  reg [49:0] FpAdd_8U_23U_int_mant_p1_3_lpi_1_dfm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10613" *)
  reg [49:0] FpAdd_8U_23U_int_mant_p1_3_lpi_1_dfm_5;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11089" *)
  wire FpAdd_8U_23U_int_mant_p1_and_12_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11116" *)
  wire FpAdd_8U_23U_int_mant_p1_and_4_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10817" *)
  wire FpAdd_8U_23U_int_mant_p1_and_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10499" *)
  reg [49:0] FpAdd_8U_23U_int_mant_p1_lpi_1_dfm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10618" *)
  reg [49:0] FpAdd_8U_23U_int_mant_p1_lpi_1_dfm_5;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11076" *)
  wire FpAdd_8U_23U_int_mant_p1_or_3_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10847" *)
  wire FpAdd_8U_23U_is_a_greater_lor_1_lpi_1_dfm_1_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10525" *)
  reg FpAdd_8U_23U_is_a_greater_lor_1_lpi_1_dfm_6;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10848" *)
  wire FpAdd_8U_23U_is_a_greater_lor_2_lpi_1_dfm_1_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10524" *)
  reg FpAdd_8U_23U_is_a_greater_lor_2_lpi_1_dfm_6;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10849" *)
  wire FpAdd_8U_23U_is_a_greater_lor_3_lpi_1_dfm_1_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10526" *)
  reg FpAdd_8U_23U_is_a_greater_lor_3_lpi_1_dfm_6;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10850" *)
  wire FpAdd_8U_23U_is_a_greater_lor_lpi_1_dfm_1_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10527" *)
  reg FpAdd_8U_23U_is_a_greater_lor_lpi_1_dfm_6;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11162" *)
  wire FpAdd_8U_23U_is_a_greater_oif_aelse_acc_1_itm_23_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11887" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22" *)
  wire [23:0] FpAdd_8U_23U_is_a_greater_oif_aelse_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11163" *)
  wire FpAdd_8U_23U_is_a_greater_oif_aelse_acc_2_itm_23_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11889" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22" *)
  wire [23:0] FpAdd_8U_23U_is_a_greater_oif_aelse_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11164" *)
  wire FpAdd_8U_23U_is_a_greater_oif_aelse_acc_3_itm_23_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11891" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22" *)
  wire [23:0] FpAdd_8U_23U_is_a_greater_oif_aelse_acc_3_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11161" *)
  wire FpAdd_8U_23U_is_a_greater_oif_aelse_acc_itm_23_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11885" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22" *)
  wire [23:0] FpAdd_8U_23U_is_a_greater_oif_aelse_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11071" *)
  wire FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_or_7_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11115" *)
  wire FpAdd_8U_23U_is_addition_and_8_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10819" *)
  wire FpAdd_8U_23U_is_addition_and_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10973" *)
  wire FpAdd_8U_23U_is_inf_1_lpi_1_dfm_2_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10518" *)
  reg FpAdd_8U_23U_is_inf_1_lpi_1_dfm_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10972" *)
  wire FpAdd_8U_23U_is_inf_2_lpi_1_dfm_2_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10515" *)
  reg FpAdd_8U_23U_is_inf_2_lpi_1_dfm_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10971" *)
  wire FpAdd_8U_23U_is_inf_3_lpi_1_dfm_2_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10512" *)
  reg FpAdd_8U_23U_is_inf_3_lpi_1_dfm_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10974" *)
  wire FpAdd_8U_23U_is_inf_lpi_1_dfm_2_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10521" *)
  reg FpAdd_8U_23U_is_inf_lpi_1_dfm_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11354" *)
  wire FpAdd_8U_23U_is_inf_mux_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11345" *)
  wire FpAdd_8U_23U_is_inf_mux_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11324" *)
  wire FpAdd_8U_23U_is_inf_mux_3_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11363" *)
  wire FpAdd_8U_23U_is_inf_mux_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10520" *)
  reg [7:0] FpAdd_8U_23U_o_expo_1_lpi_1_dfm_13;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10967" *)
  wire [7:0] FpAdd_8U_23U_o_expo_1_lpi_1_dfm_2_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10517" *)
  reg [7:0] FpAdd_8U_23U_o_expo_2_lpi_1_dfm_13;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10968" *)
  wire [7:0] FpAdd_8U_23U_o_expo_2_lpi_1_dfm_2_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10514" *)
  reg [7:0] FpAdd_8U_23U_o_expo_3_lpi_1_dfm_13;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10969" *)
  wire [7:0] FpAdd_8U_23U_o_expo_3_lpi_1_dfm_2_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11077" *)
  wire FpAdd_8U_23U_o_expo_FpAdd_8U_23U_o_expo_or_2_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10523" *)
  reg [7:0] FpAdd_8U_23U_o_expo_lpi_1_dfm_13;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10970" *)
  wire [7:0] FpAdd_8U_23U_o_expo_lpi_1_dfm_2_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10484" *)
  reg [7:0] FpAdd_8U_23U_qr_2_lpi_1_dfm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10599" *)
  reg [7:0] FpAdd_8U_23U_qr_2_lpi_1_dfm_6;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10600" *)
  reg [7:0] FpAdd_8U_23U_qr_2_lpi_1_dfm_7;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10977" *)
  wire FpAdd_8U_23U_qr_2_lpi_1_dfm_mx0c1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10488" *)
  reg [7:0] FpAdd_8U_23U_qr_3_lpi_1_dfm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10604" *)
  reg [7:0] FpAdd_8U_23U_qr_3_lpi_1_dfm_6;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10605" *)
  reg [7:0] FpAdd_8U_23U_qr_3_lpi_1_dfm_7;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10978" *)
  wire FpAdd_8U_23U_qr_3_lpi_1_dfm_mx0c1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10492" *)
  reg [7:0] FpAdd_8U_23U_qr_4_lpi_1_dfm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10609" *)
  reg [7:0] FpAdd_8U_23U_qr_4_lpi_1_dfm_6;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10610" *)
  reg [7:0] FpAdd_8U_23U_qr_4_lpi_1_dfm_7;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10979" *)
  wire FpAdd_8U_23U_qr_4_lpi_1_dfm_mx0c1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10496" *)
  reg [7:0] FpAdd_8U_23U_qr_lpi_1_dfm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10614" *)
  reg [7:0] FpAdd_8U_23U_qr_lpi_1_dfm_6;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10615" *)
  reg [7:0] FpAdd_8U_23U_qr_lpi_1_dfm_7;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10980" *)
  wire FpAdd_8U_23U_qr_lpi_1_dfm_mx0c1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11189" *)
  wire [21:0] FpAlu_8U_23U_FpAlu_8U_23U_mux_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11174" *)
  wire [21:0] FpAlu_8U_23U_FpAlu_8U_23U_mux_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11107" *)
  wire FpAlu_8U_23U_and_102_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11654" *)
  wire [7:0] FpAlu_8U_23U_and_10_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11651" *)
  wire [21:0] FpAlu_8U_23U_and_11_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10783" *)
  wire FpAlu_8U_23U_and_12_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10795" *)
  wire FpAlu_8U_23U_and_24_m1c;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11022" *)
  wire FpAlu_8U_23U_and_30_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11023" *)
  wire FpAlu_8U_23U_and_31_m1c;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10793" *)
  wire FpAlu_8U_23U_and_34_m1c;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10791" *)
  wire FpAlu_8U_23U_and_36_m1c;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10788" *)
  wire FpAlu_8U_23U_and_38_m1c;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10710" *)
  reg FpAlu_8U_23U_and_3_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11053" *)
  wire FpAlu_8U_23U_and_40_m1c;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11024" *)
  wire FpAlu_8U_23U_and_44_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11025" *)
  wire FpAlu_8U_23U_and_45_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11050" *)
  wire FpAlu_8U_23U_and_48_m1c;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11176" *)
  wire [7:0] FpAlu_8U_23U_and_4_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11051" *)
  wire FpAlu_8U_23U_and_52_m1c;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11052" *)
  wire FpAlu_8U_23U_and_56_m1c;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11173" *)
  wire [21:0] FpAlu_8U_23U_and_5_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11803" *)
  wire FpAlu_8U_23U_and_61_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11722" *)
  wire FpAlu_8U_23U_and_62_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11595" *)
  wire FpAlu_8U_23U_and_66_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11596" *)
  wire FpAlu_8U_23U_and_67_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11597" *)
  wire FpAlu_8U_23U_and_68_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11598" *)
  wire FpAlu_8U_23U_and_69_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10704" *)
  reg FpAlu_8U_23U_and_6_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11599" *)
  wire FpAlu_8U_23U_and_72_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11600" *)
  wire FpAlu_8U_23U_and_73_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11587" *)
  wire FpAlu_8U_23U_and_74_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11588" *)
  wire FpAlu_8U_23U_and_75_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11589" *)
  wire FpAlu_8U_23U_and_76_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11590" *)
  wire FpAlu_8U_23U_and_77_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11191" *)
  wire [7:0] FpAlu_8U_23U_and_7_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11591" *)
  wire FpAlu_8U_23U_and_80_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11593" *)
  wire FpAlu_8U_23U_and_81_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11083" *)
  wire FpAlu_8U_23U_and_82_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11094" *)
  wire FpAlu_8U_23U_and_88_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11188" *)
  wire [21:0] FpAlu_8U_23U_and_8_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11103" *)
  wire FpAlu_8U_23U_and_94_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11518" *)
  wire FpAlu_8U_23U_and_9_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11519" *)
  wire FpAlu_8U_23U_and_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10785" *)
  wire FpAlu_8U_23U_equal_tmp_1_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10558" *)
  reg FpAlu_8U_23U_equal_tmp_21;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10559" *)
  reg FpAlu_8U_23U_equal_tmp_22;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10560" *)
  reg FpAlu_8U_23U_equal_tmp_23;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10561" *)
  reg FpAlu_8U_23U_equal_tmp_24;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10562" *)
  reg FpAlu_8U_23U_equal_tmp_25;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10563" *)
  reg FpAlu_8U_23U_equal_tmp_26;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10567" *)
  reg FpAlu_8U_23U_equal_tmp_27;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10568" *)
  reg FpAlu_8U_23U_equal_tmp_28;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10569" *)
  reg FpAlu_8U_23U_equal_tmp_29;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10784" *)
  wire FpAlu_8U_23U_equal_tmp_2_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10570" *)
  reg FpAlu_8U_23U_equal_tmp_30;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10571" *)
  reg FpAlu_8U_23U_equal_tmp_31;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10572" *)
  reg FpAlu_8U_23U_equal_tmp_32;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10573" *)
  reg FpAlu_8U_23U_equal_tmp_33;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10574" *)
  reg FpAlu_8U_23U_equal_tmp_34;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10575" *)
  reg FpAlu_8U_23U_equal_tmp_35;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10796" *)
  wire FpAlu_8U_23U_equal_tmp_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11576" *)
  wire FpAlu_8U_23U_mux1h_144_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11177" *)
  wire [7:0] FpAlu_8U_23U_mux1h_145_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11172" *)
  wire FpAlu_8U_23U_mux1h_147_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11579" *)
  wire FpAlu_8U_23U_mux1h_148_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11192" *)
  wire [7:0] FpAlu_8U_23U_mux1h_149_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11187" *)
  wire FpAlu_8U_23U_mux1h_151_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10695" *)
  reg FpAlu_8U_23U_mux1h_152_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11655" *)
  wire [7:0] FpAlu_8U_23U_mux1h_153_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11652" *)
  wire [21:0] FpAlu_8U_23U_mux1h_154_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11650" *)
  wire FpAlu_8U_23U_mux1h_155_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10686" *)
  reg FpAlu_8U_23U_mux1h_33_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11715" *)
  wire [7:0] FpAlu_8U_23U_mux1h_34_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11713" *)
  wire [21:0] FpAlu_8U_23U_mux1h_35_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11559" *)
  wire FpAlu_8U_23U_mux_20_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11557" *)
  wire FpAlu_8U_23U_mux_21_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10564" *)
  reg FpAlu_8U_23U_nor_dfs_4;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10565" *)
  reg FpAlu_8U_23U_nor_dfs_5;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10566" *)
  reg FpAlu_8U_23U_nor_dfs_6;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10789" *)
  wire FpAlu_8U_23U_nor_dfs_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11019" *)
  wire FpAlu_8U_23U_o_0_lpi_1_dfm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10504" *)
  reg FpAlu_8U_23U_o_0_lpi_1_dfm_4;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10982" *)
  wire FpAlu_8U_23U_o_0_sva_2_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10579" *)
  reg FpAlu_8U_23U_o_0_sva_7;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10580" *)
  reg FpAlu_8U_23U_o_0_sva_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10581" *)
  reg FpAlu_8U_23U_o_0_sva_9;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11020" *)
  wire [21:0] FpAlu_8U_23U_o_22_1_lpi_1_dfm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10503" *)
  reg [21:0] FpAlu_8U_23U_o_22_1_lpi_1_dfm_4;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11021" *)
  wire [7:0] FpAlu_8U_23U_o_30_23_lpi_1_dfm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10502" *)
  reg [7:0] FpAlu_8U_23U_o_30_23_lpi_1_dfm_4;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11092" *)
  wire FpAlu_8U_23U_o_FpAlu_8U_23U_o_or_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11577" *)
  wire FpAlu_8U_23U_or_145_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11578" *)
  wire FpAlu_8U_23U_or_146_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11580" *)
  wire FpAlu_8U_23U_or_147_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11581" *)
  wire FpAlu_8U_23U_or_148_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11120" *)
  wire FpAlu_8U_23U_or_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11805" *)
  wire FpCmp_8U_23U_false_else_1_FpCmp_8U_23U_false_else_1_and_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11785" *)
  (* unused_bits = "0 1 2 3 4 5 6 7" *)
  wire [8:0] FpCmp_8U_23U_false_else_if_acc_10_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11764" *)
  (* unused_bits = "0 1 2 3 4 5 6 7" *)
  wire [8:0] FpCmp_8U_23U_false_else_if_acc_4_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11157" *)
  wire FpCmp_8U_23U_false_else_if_acc_6_itm_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11819" *)
  (* unused_bits = "0 1 2 3 4 5 6 7" *)
  wire [8:0] FpCmp_8U_23U_false_else_if_acc_6_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11777" *)
  (* unused_bits = "0 1 2 3 4 5 6 7" *)
  wire [8:0] FpCmp_8U_23U_false_else_if_acc_8_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11806" *)
  wire FpCmp_8U_23U_false_if_1_FpCmp_8U_23U_false_if_1_or_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10797" *)
  wire FpCmp_8U_23U_false_is_abs_a_greater_2_lpi_1_dfm_1_mx0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10993" *)
  wire FpCmp_8U_23U_false_is_abs_a_greater_2_lpi_1_dfm_1_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10500" *)
  reg FpCmp_8U_23U_false_is_abs_a_greater_2_lpi_1_dfm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11804" *)
  wire FpCmp_8U_23U_false_mux_4_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11046" *)
  wire [31:0] FpCmp_8U_23U_false_o_1_lpi_1_dfm_1_mx0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10754" *)
  reg [30:0] FpCmp_8U_23U_false_o_1_lpi_1_dfm_6_30_0_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10755" *)
  reg [30:0] FpCmp_8U_23U_false_o_1_lpi_1_dfm_7_30_0_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11049" *)
  wire [31:0] FpCmp_8U_23U_false_o_2_lpi_1_dfm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10752" *)
  reg [30:0] FpCmp_8U_23U_false_o_2_lpi_1_dfm_7_30_0_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10753" *)
  reg [30:0] FpCmp_8U_23U_false_o_2_lpi_1_dfm_8_30_0_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11047" *)
  wire [31:0] FpCmp_8U_23U_false_o_3_lpi_1_dfm_1_mx0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10750" *)
  reg [30:0] FpCmp_8U_23U_false_o_3_lpi_1_dfm_7_30_0_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10751" *)
  reg [30:0] FpCmp_8U_23U_false_o_3_lpi_1_dfm_8_30_0_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11085" *)
  wire FpCmp_8U_23U_false_o_and_1_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11095" *)
  wire FpCmp_8U_23U_false_o_and_6_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11048" *)
  wire [31:0] FpCmp_8U_23U_false_o_lpi_1_dfm_1_mx0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10748" *)
  reg [30:0] FpCmp_8U_23U_false_o_lpi_1_dfm_8_30_0_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10749" *)
  reg [30:0] FpCmp_8U_23U_false_o_lpi_1_dfm_9_30_0_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11158" *)
  wire FpCmp_8U_23U_true_else_else_if_acc_4_itm_23;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11821" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22" *)
  wire [23:0] FpCmp_8U_23U_true_else_else_if_acc_4_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11783" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22" *)
  wire [23:0] FpCmp_8U_23U_true_else_else_if_acc_6_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11775" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22" *)
  wire [23:0] FpCmp_8U_23U_true_else_else_if_acc_7_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11766" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22" *)
  wire [23:0] FpCmp_8U_23U_true_else_else_if_acc_8_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11160" *)
  wire FpCmp_8U_23U_true_if_acc_10_itm_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11826" *)
  (* unused_bits = "0 1 2 3 4 5 6 7" *)
  wire [8:0] FpCmp_8U_23U_true_if_acc_10_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11155" *)
  wire FpCmp_8U_23U_true_if_acc_4_itm_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11815" *)
  (* unused_bits = "0 1 2 3 4 5 6 7" *)
  wire [8:0] FpCmp_8U_23U_true_if_acc_4_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11156" *)
  wire FpCmp_8U_23U_true_if_acc_6_itm_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11817" *)
  (* unused_bits = "0 1 2 3 4 5 6 7" *)
  wire [8:0] FpCmp_8U_23U_true_if_acc_6_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11159" *)
  wire FpCmp_8U_23U_true_if_acc_8_itm_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11824" *)
  (* unused_bits = "0 1 2 3 4 5 6 7" *)
  wire [8:0] FpCmp_8U_23U_true_if_acc_8_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11042" *)
  wire [31:0] FpCmp_8U_23U_true_o_1_lpi_1_dfm_1_mx0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10765" *)
  reg [30:0] FpCmp_8U_23U_true_o_1_lpi_1_dfm_5_30_0_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10766" *)
  reg [30:0] FpCmp_8U_23U_true_o_1_lpi_1_dfm_6_30_0_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10767" *)
  reg [30:0] FpCmp_8U_23U_true_o_1_lpi_1_dfm_7_30_0_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11043" *)
  wire [31:0] FpCmp_8U_23U_true_o_2_lpi_1_dfm_1_mx0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10762" *)
  reg [30:0] FpCmp_8U_23U_true_o_2_lpi_1_dfm_5_30_0_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10763" *)
  reg [30:0] FpCmp_8U_23U_true_o_2_lpi_1_dfm_6_30_0_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10764" *)
  reg [30:0] FpCmp_8U_23U_true_o_2_lpi_1_dfm_7_30_0_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11044" *)
  wire [31:0] FpCmp_8U_23U_true_o_3_lpi_1_dfm_1_mx0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10759" *)
  reg [30:0] FpCmp_8U_23U_true_o_3_lpi_1_dfm_5_30_0_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10760" *)
  reg [30:0] FpCmp_8U_23U_true_o_3_lpi_1_dfm_6_30_0_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10761" *)
  reg [30:0] FpCmp_8U_23U_true_o_3_lpi_1_dfm_7_30_0_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11093" *)
  wire FpCmp_8U_23U_true_o_and_5_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11102" *)
  wire FpCmp_8U_23U_true_o_and_9_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11084" *)
  wire FpCmp_8U_23U_true_o_and_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11045" *)
  wire [31:0] FpCmp_8U_23U_true_o_lpi_1_dfm_1_mx0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10756" *)
  reg [30:0] FpCmp_8U_23U_true_o_lpi_1_dfm_5_30_0_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10757" *)
  reg [30:0] FpCmp_8U_23U_true_o_lpi_1_dfm_6_30_0_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10758" *)
  reg [30:0] FpCmp_8U_23U_true_o_lpi_1_dfm_7_30_0_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11117" *)
  wire FpMantRNE_49U_24U_else_and_4_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10815" *)
  wire FpMantRNE_49U_24U_else_and_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11017" *)
  wire FpMantRNE_49U_24U_else_carry_1_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11015" *)
  wire FpMantRNE_49U_24U_else_carry_2_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11013" *)
  wire FpMantRNE_49U_24U_else_carry_3_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11011" *)
  wire FpMantRNE_49U_24U_else_carry_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11712" *)
  wire [48:0] FpNormalize_8U_49U_FpNormalize_8U_49U_and_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11711" *)
  wire [48:0] FpNormalize_8U_49U_FpNormalize_8U_49U_and_3_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11710" *)
  wire [48:0] FpNormalize_8U_49U_FpNormalize_8U_49U_and_5_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11709" *)
  wire [48:0] FpNormalize_8U_49U_FpNormalize_8U_49U_and_7_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11671" *)
  wire [5:0] FpNormalize_8U_49U_else_mux_4_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11675" *)
  wire [5:0] FpNormalize_8U_49U_else_mux_5_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11679" *)
  wire [5:0] FpNormalize_8U_49U_else_mux_6_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11683" *)
  wire [5:0] FpNormalize_8U_49U_else_mux_7_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10642" *)
  reg FpNormalize_8U_49U_if_or_1_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10643" *)
  reg FpNormalize_8U_49U_if_or_1_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10963" *)
  wire FpNormalize_8U_49U_if_or_1_itm_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10655" *)
  reg FpNormalize_8U_49U_if_or_2_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10656" *)
  reg FpNormalize_8U_49U_if_or_2_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10964" *)
  wire FpNormalize_8U_49U_if_or_2_itm_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10668" *)
  reg FpNormalize_8U_49U_if_or_3_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10669" *)
  reg FpNormalize_8U_49U_if_or_3_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10965" *)
  wire FpNormalize_8U_49U_if_or_3_itm_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10630" *)
  reg FpNormalize_8U_49U_if_or_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10631" *)
  reg FpNormalize_8U_49U_if_or_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10962" *)
  wire FpNormalize_8U_49U_if_or_itm_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11055" *)
  wire FpNormalize_8U_49U_oelse_not_11;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11056" *)
  wire FpNormalize_8U_49U_oelse_not_13;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11057" *)
  wire FpNormalize_8U_49U_oelse_not_15;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11054" *)
  wire FpNormalize_8U_49U_oelse_not_9;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11748" *)
  wire IntSaturation_33U_32U_IntSaturation_33U_32U_nor_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11752" *)
  wire IntSaturation_33U_32U_IntSaturation_33U_32U_nor_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11750" *)
  wire IntSaturation_33U_32U_IntSaturation_33U_32U_nor_3_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11754" *)
  wire IntSaturation_33U_32U_IntSaturation_33U_32U_nor_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11478" *)
  wire IntSaturation_33U_32U_IntSaturation_33U_32U_or_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11477" *)
  wire IntSaturation_33U_32U_IntSaturation_33U_32U_or_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11476" *)
  wire IntSaturation_33U_32U_IntSaturation_33U_32U_or_3_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11096" *)
  wire IntSaturation_33U_32U_IntSaturation_33U_32U_or_7_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11468" *)
  wire IntSaturation_33U_32U_IntSaturation_33U_32U_or_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11097" *)
  wire IntSaturation_33U_32U_and_11_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11755" *)
  wire IntSaturation_33U_32U_and_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11749" *)
  wire IntSaturation_33U_32U_and_3_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11753" *)
  wire IntSaturation_33U_32U_and_5_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11751" *)
  wire IntSaturation_33U_32U_and_7_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11088" *)
  wire IntSaturation_33U_32U_and_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11106" *)
  wire IntSaturation_33U_32U_if_and_9_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11041" *)
  wire [30:0] IntSaturation_33U_32U_o_31_1_1_lpi_1_dfm_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11038" *)
  wire [30:0] IntSaturation_33U_32U_o_31_1_2_lpi_1_dfm_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11040" *)
  wire [30:0] IntSaturation_33U_32U_o_31_1_3_lpi_1_dfm_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11039" *)
  wire [30:0] IntSaturation_33U_32U_o_31_1_lpi_1_dfm_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10714" *)
  reg [21:0] IntSaturation_33U_32U_slc_IntSaturation_33U_32U_o_31_1_1_21_0_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10713" *)
  reg [7:0] IntSaturation_33U_32U_slc_IntSaturation_33U_32U_o_31_1_1_29_22_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10702" *)
  reg [21:0] IntSaturation_33U_32U_slc_IntSaturation_33U_32U_o_31_1_21_0_itm_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10703" *)
  reg [21:0] IntSaturation_33U_32U_slc_IntSaturation_33U_32U_o_31_1_21_0_itm_4;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10701" *)
  reg [7:0] IntSaturation_33U_32U_slc_IntSaturation_33U_32U_o_31_1_29_22_itm_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10708" *)
  reg [21:0] IntSaturation_33U_32U_slc_IntSaturation_33U_32U_o_31_1_2_21_0_itm_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10709" *)
  reg [21:0] IntSaturation_33U_32U_slc_IntSaturation_33U_32U_o_31_1_2_21_0_itm_4;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10707" *)
  reg [7:0] IntSaturation_33U_32U_slc_IntSaturation_33U_32U_o_31_1_2_29_22_itm_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10697" *)
  reg [21:0] IntSaturation_33U_32U_slc_IntSaturation_33U_32U_o_31_1_3_21_0_itm_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10698" *)
  reg [21:0] IntSaturation_33U_32U_slc_IntSaturation_33U_32U_o_31_1_3_21_0_itm_4;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10696" *)
  reg [7:0] IntSaturation_33U_32U_slc_IntSaturation_33U_32U_o_31_1_3_29_22_itm_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11082" *)
  wire IsNaN_8U_23U_1_aelse_and_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10553" *)
  reg IsNaN_8U_23U_1_land_1_lpi_1_dfm_7;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10554" *)
  reg IsNaN_8U_23U_1_land_1_lpi_1_dfm_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10555" *)
  reg IsNaN_8U_23U_1_land_1_lpi_1_dfm_9;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10790" *)
  wire IsNaN_8U_23U_1_land_1_lpi_1_dfm_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10550" *)
  reg IsNaN_8U_23U_1_land_2_lpi_1_dfm_7;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10551" *)
  reg IsNaN_8U_23U_1_land_2_lpi_1_dfm_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10552" *)
  reg IsNaN_8U_23U_1_land_2_lpi_1_dfm_9;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10787" *)
  wire IsNaN_8U_23U_1_land_2_lpi_1_dfm_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10547" *)
  reg IsNaN_8U_23U_1_land_3_lpi_1_dfm_7;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10548" *)
  reg IsNaN_8U_23U_1_land_3_lpi_1_dfm_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10549" *)
  reg IsNaN_8U_23U_1_land_3_lpi_1_dfm_9;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10792" *)
  wire IsNaN_8U_23U_1_land_3_lpi_1_dfm_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10544" *)
  reg IsNaN_8U_23U_1_land_lpi_1_dfm_7;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10545" *)
  reg IsNaN_8U_23U_1_land_lpi_1_dfm_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10546" *)
  reg IsNaN_8U_23U_1_land_lpi_1_dfm_9;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10794" *)
  wire IsNaN_8U_23U_1_land_lpi_1_dfm_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10676" *)
  reg IsNaN_8U_23U_2_IsNaN_8U_23U_2_nor_1_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10677" *)
  reg IsNaN_8U_23U_2_IsNaN_8U_23U_2_nor_1_itm_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10990" *)
  wire IsNaN_8U_23U_2_IsNaN_8U_23U_2_nor_1_itm_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10678" *)
  reg IsNaN_8U_23U_2_IsNaN_8U_23U_2_nor_2_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10679" *)
  reg IsNaN_8U_23U_2_IsNaN_8U_23U_2_nor_2_itm_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10988" *)
  wire IsNaN_8U_23U_2_IsNaN_8U_23U_2_nor_2_itm_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10680" *)
  reg IsNaN_8U_23U_2_IsNaN_8U_23U_2_nor_3_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10681" *)
  reg IsNaN_8U_23U_2_IsNaN_8U_23U_2_nor_3_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10991" *)
  wire IsNaN_8U_23U_2_IsNaN_8U_23U_2_nor_3_itm_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10674" *)
  reg IsNaN_8U_23U_2_IsNaN_8U_23U_2_nor_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10675" *)
  reg IsNaN_8U_23U_2_IsNaN_8U_23U_2_nor_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10989" *)
  wire IsNaN_8U_23U_2_IsNaN_8U_23U_2_nor_itm_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11111" *)
  wire IsNaN_8U_23U_2_IsNaN_8U_23U_2_or_3_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11109" *)
  wire IsNaN_8U_23U_2_IsNaN_8U_23U_2_or_5_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11110" *)
  wire IsNaN_8U_23U_2_IsNaN_8U_23U_4_or_2_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11121" *)
  wire IsNaN_8U_23U_2_and_6_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11166" *)
  wire IsNaN_8U_23U_2_and_9_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10828" *)
  wire IsNaN_8U_23U_2_and_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10800" *)
  wire IsNaN_8U_23U_2_nor_2_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10798" *)
  wire IsNaN_8U_23U_2_nor_3_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10346" *)
  wire IsNaN_8U_23U_3_nor_10_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10349" *)
  wire IsNaN_8U_23U_3_nor_4_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10348" *)
  wire IsNaN_8U_23U_3_nor_6_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10347" *)
  wire IsNaN_8U_23U_3_nor_8_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10801" *)
  wire IsNaN_8U_23U_4_IsNaN_8U_23U_4_nand_2_itm_mx0w2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10799" *)
  wire IsNaN_8U_23U_4_IsNaN_8U_23U_4_nand_3_itm_mx0w2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10683" *)
  reg IsNaN_8U_23U_4_nor_2_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10684" *)
  reg IsNaN_8U_23U_4_nor_3_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10685" *)
  reg IsNaN_8U_23U_4_nor_3_itm_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11091" *)
  wire IsNaN_8U_23U_aelse_and_12_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11100" *)
  wire IsNaN_8U_23U_aelse_and_16_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11081" *)
  wire IsNaN_8U_23U_aelse_and_8_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11072" *)
  wire IsNaN_8U_23U_aelse_and_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10534" *)
  reg IsNaN_8U_23U_land_1_lpi_1_dfm_10;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10535" *)
  reg IsNaN_8U_23U_land_1_lpi_1_dfm_11;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10532" *)
  reg IsNaN_8U_23U_land_1_lpi_1_dfm_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10533" *)
  reg IsNaN_8U_23U_land_1_lpi_1_dfm_9;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10727" *)
  reg IsNaN_8U_23U_land_1_lpi_1_dfm_st_4;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10728" *)
  reg IsNaN_8U_23U_land_1_lpi_1_dfm_st_5;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10530" *)
  reg IsNaN_8U_23U_land_2_lpi_1_dfm_10;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10531" *)
  reg IsNaN_8U_23U_land_2_lpi_1_dfm_11;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10528" *)
  reg IsNaN_8U_23U_land_2_lpi_1_dfm_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10529" *)
  reg IsNaN_8U_23U_land_2_lpi_1_dfm_9;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10732" *)
  reg IsNaN_8U_23U_land_2_lpi_1_dfm_st_4;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10733" *)
  reg IsNaN_8U_23U_land_2_lpi_1_dfm_st_5;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10538" *)
  reg IsNaN_8U_23U_land_3_lpi_1_dfm_10;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10539" *)
  reg IsNaN_8U_23U_land_3_lpi_1_dfm_11;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10536" *)
  reg IsNaN_8U_23U_land_3_lpi_1_dfm_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10537" *)
  reg IsNaN_8U_23U_land_3_lpi_1_dfm_9;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10737" *)
  reg IsNaN_8U_23U_land_3_lpi_1_dfm_st_4;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10738" *)
  reg IsNaN_8U_23U_land_3_lpi_1_dfm_st_5;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10542" *)
  reg IsNaN_8U_23U_land_lpi_1_dfm_10;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10543" *)
  reg IsNaN_8U_23U_land_lpi_1_dfm_11;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10540" *)
  reg IsNaN_8U_23U_land_lpi_1_dfm_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10541" *)
  reg IsNaN_8U_23U_land_lpi_1_dfm_9;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10742" *)
  reg IsNaN_8U_23U_land_lpi_1_dfm_st_4;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10743" *)
  reg IsNaN_8U_23U_land_lpi_1_dfm_st_5;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10859" *)
  wire IsZero_8U_23U_1_and_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11118" *)
  wire IsZero_8U_23U_and_4_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11099" *)
  wire IsZero_8U_23U_and_6_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11728" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31 32" *)
  wire [33:0] acc_10_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11732" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31 32" *)
  wire [33:0] acc_11_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11909" *)
  (* unused_bits = "0" *)
  wire [50:0] acc_12_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11913" *)
  (* unused_bits = "0" *)
  wire [50:0] acc_13_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11917" *)
  (* unused_bits = "0" *)
  wire [50:0] acc_14_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11921" *)
  (* unused_bits = "0" *)
  wire [50:0] acc_15_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11673" *)
  (* unused_bits = "0" *)
  wire [8:0] acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11677" *)
  (* unused_bits = "0" *)
  wire [8:0] acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11681" *)
  (* unused_bits = "0" *)
  wire [8:0] acc_3_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11893" *)
  (* unused_bits = "0" *)
  wire [8:0] acc_4_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11897" *)
  (* unused_bits = "0" *)
  wire [8:0] acc_5_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11901" *)
  (* unused_bits = "0" *)
  wire [8:0] acc_6_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11905" *)
  (* unused_bits = "0" *)
  wire [8:0] acc_7_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11724" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31 32" *)
  wire [33:0] acc_8_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11736" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31 32" *)
  wire [33:0] acc_9_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11669" *)
  (* unused_bits = "0" *)
  wire [8:0] acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10822" *)
  wire alu_loop_bypass_if_and_6_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10823" *)
  wire alu_loop_bypass_if_and_7_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10626" *)
  reg alu_loop_op_1_FpAdd_8U_23U_IsZero_8U_23U_1_or_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10627" *)
  reg alu_loop_op_1_FpAdd_8U_23U_IsZero_8U_23U_1_or_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10958" *)
  wire alu_loop_op_1_FpAdd_8U_23U_IsZero_8U_23U_1_or_itm_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10625" *)
  reg alu_loop_op_1_FpAdd_8U_23U_IsZero_8U_23U_or_itm_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10994" *)
  wire alu_loop_op_1_FpAdd_8U_23U_IsZero_8U_23U_or_itm_mx0w2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12006" *)
  wire [7:0] alu_loop_op_1_FpAdd_8U_23U_a_left_shift_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11929" *)
  wire [7:0] alu_loop_op_1_FpAdd_8U_23U_b_left_shift_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11143" *)
  wire alu_loop_op_1_FpAdd_8U_23U_if_3_if_acc_1_itm_7_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11701" *)
  (* unused_bits = "0 1 2 3 4 5 6" *)
  wire [7:0] alu_loop_op_1_FpAdd_8U_23U_if_3_if_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11147" *)
  wire alu_loop_op_1_FpAdd_8U_23U_if_4_if_acc_1_itm_7_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11740" *)
  (* unused_bits = "0 1 2 3 4 5 6" *)
  wire [7:0] alu_loop_op_1_FpAdd_8U_23U_if_4_if_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11178" *)
  wire [7:0] alu_loop_op_1_FpAdd_8U_23U_if_4_if_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10633" *)
  reg alu_loop_op_1_FpAdd_8U_23U_if_4_if_slc_FpAdd_8U_23U_if_4_if_acc_1_7_svs_st_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10726" *)
  reg alu_loop_op_1_FpAdd_8U_23U_if_4_if_slc_FpAdd_8U_23U_if_4_if_acc_1_7_svs_st_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10341" *)
  wire alu_loop_op_1_FpAdd_8U_23U_is_a_greater_oif_equal_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10957" *)
  wire alu_loop_op_1_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10628" *)
  reg alu_loop_op_1_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_st;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10629" *)
  reg alu_loop_op_1_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10722" *)
  reg alu_loop_op_1_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11361" *)
  wire [22:0] alu_loop_op_1_FpMantRNE_49U_24U_else_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10632" *)
  reg alu_loop_op_1_FpMantRNE_49U_24U_else_and_svs_st;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10725" *)
  reg alu_loop_op_1_FpMantRNE_49U_24U_else_and_svs_st_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10345" *)
  wire alu_loop_op_1_FpMantRNE_49U_24U_else_and_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11807" *)
  (* unused_bits = "0 1 2 3 4 5 6 7" *)
  wire [8:0] alu_loop_op_1_FpNormalize_8U_49U_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10911" *)
  wire [48:0] alu_loop_op_1_FpNormalize_8U_49U_else_lshift_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11151" *)
  wire alu_loop_op_1_IntSaturation_33U_32U_else_if_acc_itm_2_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11756" *)
  (* unused_bits = "0 1" *)
  wire [2:0] alu_loop_op_1_IntSaturation_33U_32U_else_if_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11142" *)
  wire alu_loop_op_1_IntSaturation_33U_32U_if_acc_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11699" *)
  (* unused_bits = "0 1" *)
  wire [2:0] alu_loop_op_1_IntSaturation_33U_32U_if_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10557" *)
  reg alu_loop_op_1_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_svs_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10638" *)
  reg alu_loop_op_2_FpAdd_8U_23U_IsZero_8U_23U_1_or_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10639" *)
  reg alu_loop_op_2_FpAdd_8U_23U_IsZero_8U_23U_1_or_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10954" *)
  wire alu_loop_op_2_FpAdd_8U_23U_IsZero_8U_23U_1_or_itm_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10636" *)
  reg alu_loop_op_2_FpAdd_8U_23U_IsZero_8U_23U_or_itm_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10637" *)
  reg alu_loop_op_2_FpAdd_8U_23U_IsZero_8U_23U_or_itm_4;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10981" *)
  wire alu_loop_op_2_FpAdd_8U_23U_IsZero_8U_23U_or_itm_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11995" *)
  wire [7:0] alu_loop_op_2_FpAdd_8U_23U_a_left_shift_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11940" *)
  wire [7:0] alu_loop_op_2_FpAdd_8U_23U_b_left_shift_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11144" *)
  wire alu_loop_op_2_FpAdd_8U_23U_if_3_if_acc_4_itm_7_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11703" *)
  (* unused_bits = "0 1 2 3 4 5 6" *)
  wire [7:0] alu_loop_op_2_FpAdd_8U_23U_if_3_if_acc_4_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11148" *)
  wire alu_loop_op_2_FpAdd_8U_23U_if_4_if_acc_4_itm_7_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11742" *)
  (* unused_bits = "0 1 2 3 4 5 6" *)
  wire [7:0] alu_loop_op_2_FpAdd_8U_23U_if_4_if_acc_4_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11193" *)
  wire [7:0] alu_loop_op_2_FpAdd_8U_23U_if_4_if_acc_5_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10645" *)
  reg alu_loop_op_2_FpAdd_8U_23U_if_4_if_slc_FpAdd_8U_23U_if_4_if_acc_1_7_2_svs_st_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10731" *)
  reg alu_loop_op_2_FpAdd_8U_23U_if_4_if_slc_FpAdd_8U_23U_if_4_if_acc_1_7_2_svs_st_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10340" *)
  wire alu_loop_op_2_FpAdd_8U_23U_is_a_greater_oif_equal_2_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10953" *)
  wire alu_loop_op_2_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_2_svs_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10640" *)
  reg alu_loop_op_2_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_2_svs_st;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10641" *)
  reg alu_loop_op_2_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_2_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10729" *)
  reg alu_loop_op_2_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_2_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11352" *)
  wire [22:0] alu_loop_op_2_FpMantRNE_49U_24U_else_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10644" *)
  reg alu_loop_op_2_FpMantRNE_49U_24U_else_and_2_svs_st;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10730" *)
  reg alu_loop_op_2_FpMantRNE_49U_24U_else_and_2_svs_st_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10344" *)
  wire alu_loop_op_2_FpMantRNE_49U_24U_else_and_2_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11809" *)
  (* unused_bits = "0 1 2 3 4 5 6 7" *)
  wire [8:0] alu_loop_op_2_FpNormalize_8U_49U_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10910" *)
  wire [48:0] alu_loop_op_2_FpNormalize_8U_49U_else_lshift_2_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11152" *)
  wire alu_loop_op_2_IntSaturation_33U_32U_else_if_acc_1_itm_2_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11758" *)
  (* unused_bits = "0 1" *)
  wire [2:0] alu_loop_op_2_IntSaturation_33U_32U_else_if_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11139" *)
  wire alu_loop_op_2_IntSaturation_33U_32U_if_acc_1_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11689" *)
  (* unused_bits = "0 1" *)
  wire [2:0] alu_loop_op_2_IntSaturation_33U_32U_if_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10501" *)
  reg alu_loop_op_2_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_1_svs_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10619" *)
  reg alu_loop_op_2_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_1_svs_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10651" *)
  reg alu_loop_op_3_FpAdd_8U_23U_IsZero_8U_23U_1_or_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10652" *)
  reg alu_loop_op_3_FpAdd_8U_23U_IsZero_8U_23U_1_or_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10950" *)
  wire alu_loop_op_3_FpAdd_8U_23U_IsZero_8U_23U_1_or_itm_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10648" *)
  reg alu_loop_op_3_FpAdd_8U_23U_IsZero_8U_23U_or_itm_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10649" *)
  reg alu_loop_op_3_FpAdd_8U_23U_IsZero_8U_23U_or_itm_4;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10650" *)
  reg alu_loop_op_3_FpAdd_8U_23U_IsZero_8U_23U_or_itm_5;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10976" *)
  wire alu_loop_op_3_FpAdd_8U_23U_IsZero_8U_23U_or_itm_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11984" *)
  wire [7:0] alu_loop_op_3_FpAdd_8U_23U_a_left_shift_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11951" *)
  wire [7:0] alu_loop_op_3_FpAdd_8U_23U_b_left_shift_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11145" *)
  wire alu_loop_op_3_FpAdd_8U_23U_if_3_if_acc_2_itm_7_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11705" *)
  (* unused_bits = "0 1 2 3 4 5 6" *)
  wire [7:0] alu_loop_op_3_FpAdd_8U_23U_if_3_if_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11149" *)
  wire alu_loop_op_3_FpAdd_8U_23U_if_4_if_acc_2_itm_7_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11744" *)
  (* unused_bits = "0 1 2 3 4 5 6" *)
  wire [7:0] alu_loop_op_3_FpAdd_8U_23U_if_4_if_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11656" *)
  wire [7:0] alu_loop_op_3_FpAdd_8U_23U_if_4_if_acc_3_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10658" *)
  reg alu_loop_op_3_FpAdd_8U_23U_if_4_if_slc_FpAdd_8U_23U_if_4_if_acc_1_7_1_svs_st_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10736" *)
  reg alu_loop_op_3_FpAdd_8U_23U_if_4_if_slc_FpAdd_8U_23U_if_4_if_acc_1_7_1_svs_st_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10339" *)
  wire alu_loop_op_3_FpAdd_8U_23U_is_a_greater_oif_equal_1_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10949" *)
  wire alu_loop_op_3_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_1_svs_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10653" *)
  reg alu_loop_op_3_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_1_svs_st;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10654" *)
  reg alu_loop_op_3_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_1_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10734" *)
  reg alu_loop_op_3_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_1_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11343" *)
  wire [22:0] alu_loop_op_3_FpMantRNE_49U_24U_else_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10657" *)
  reg alu_loop_op_3_FpMantRNE_49U_24U_else_and_1_svs_st;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10735" *)
  reg alu_loop_op_3_FpMantRNE_49U_24U_else_and_1_svs_st_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10343" *)
  wire alu_loop_op_3_FpMantRNE_49U_24U_else_and_1_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11811" *)
  (* unused_bits = "0 1 2 3 4 5 6 7" *)
  wire [8:0] alu_loop_op_3_FpNormalize_8U_49U_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10909" *)
  wire [48:0] alu_loop_op_3_FpNormalize_8U_49U_else_lshift_1_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11153" *)
  wire alu_loop_op_3_IntSaturation_33U_32U_else_if_acc_itm_2_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11760" *)
  (* unused_bits = "0 1" *)
  wire [2:0] alu_loop_op_3_IntSaturation_33U_32U_else_if_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11141" *)
  wire alu_loop_op_3_IntSaturation_33U_32U_if_acc_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11697" *)
  (* unused_bits = "0 1" *)
  wire [2:0] alu_loop_op_3_IntSaturation_33U_32U_if_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10556" *)
  reg alu_loop_op_3_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_svs_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10664" *)
  reg alu_loop_op_4_FpAdd_8U_23U_IsZero_8U_23U_1_or_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10665" *)
  reg alu_loop_op_4_FpAdd_8U_23U_IsZero_8U_23U_1_or_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10946" *)
  wire alu_loop_op_4_FpAdd_8U_23U_IsZero_8U_23U_1_or_itm_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10661" *)
  reg alu_loop_op_4_FpAdd_8U_23U_IsZero_8U_23U_or_itm_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10662" *)
  reg alu_loop_op_4_FpAdd_8U_23U_IsZero_8U_23U_or_itm_4;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10663" *)
  reg alu_loop_op_4_FpAdd_8U_23U_IsZero_8U_23U_or_itm_5;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10975" *)
  wire alu_loop_op_4_FpAdd_8U_23U_IsZero_8U_23U_or_itm_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11973" *)
  wire [7:0] alu_loop_op_4_FpAdd_8U_23U_a_left_shift_acc_3_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11962" *)
  wire [7:0] alu_loop_op_4_FpAdd_8U_23U_b_left_shift_acc_3_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11146" *)
  wire alu_loop_op_4_FpAdd_8U_23U_if_3_if_acc_6_itm_7_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11707" *)
  (* unused_bits = "0 1 2 3 4 5 6" *)
  wire [7:0] alu_loop_op_4_FpAdd_8U_23U_if_3_if_acc_6_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11150" *)
  wire alu_loop_op_4_FpAdd_8U_23U_if_4_if_acc_6_itm_7_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11746" *)
  (* unused_bits = "0 1 2 3 4 5 6" *)
  wire [7:0] alu_loop_op_4_FpAdd_8U_23U_if_4_if_acc_6_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11716" *)
  wire [7:0] alu_loop_op_4_FpAdd_8U_23U_if_4_if_acc_7_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10671" *)
  reg alu_loop_op_4_FpAdd_8U_23U_if_4_if_slc_FpAdd_8U_23U_if_4_if_acc_1_7_3_svs_st_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10741" *)
  reg alu_loop_op_4_FpAdd_8U_23U_if_4_if_slc_FpAdd_8U_23U_if_4_if_acc_1_7_3_svs_st_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10338" *)
  wire alu_loop_op_4_FpAdd_8U_23U_is_a_greater_oif_equal_3_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10945" *)
  wire alu_loop_op_4_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_3_svs_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10666" *)
  reg alu_loop_op_4_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_3_svs_st;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10667" *)
  reg alu_loop_op_4_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_3_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10739" *)
  reg alu_loop_op_4_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_3_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11322" *)
  wire [22:0] alu_loop_op_4_FpMantRNE_49U_24U_else_acc_3_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10670" *)
  reg alu_loop_op_4_FpMantRNE_49U_24U_else_and_3_svs_st;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10740" *)
  reg alu_loop_op_4_FpMantRNE_49U_24U_else_and_3_svs_st_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10342" *)
  wire alu_loop_op_4_FpMantRNE_49U_24U_else_and_3_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11813" *)
  (* unused_bits = "0 1 2 3 4 5 6 7" *)
  wire [8:0] alu_loop_op_4_FpNormalize_8U_49U_acc_3_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10908" *)
  wire [48:0] alu_loop_op_4_FpNormalize_8U_49U_else_lshift_3_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11154" *)
  wire alu_loop_op_4_IntSaturation_33U_32U_else_if_acc_1_itm_2_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11762" *)
  (* unused_bits = "0 1" *)
  wire [2:0] alu_loop_op_4_IntSaturation_33U_32U_else_if_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11140" *)
  wire alu_loop_op_4_IntSaturation_33U_32U_if_acc_1_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11695" *)
  (* unused_bits = "0 1" *)
  wire [2:0] alu_loop_op_4_IntSaturation_33U_32U_if_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10620" *)
  reg alu_loop_op_4_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_1_svs_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11691" *)
  wire [31:0] alu_loop_op_else_alu_loop_op_else_mux_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11687" *)
  wire [31:0] alu_loop_op_else_alu_loop_op_else_mux_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11685" *)
  wire [31:0] alu_loop_op_else_alu_loop_op_else_mux_3_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11693" *)
  wire [31:0] alu_loop_op_else_alu_loop_op_else_mux_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11027" *)
  wire [32:0] alu_loop_op_else_else_else_else_ac_int_cctor_1_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11030" *)
  wire [32:0] alu_loop_op_else_else_else_else_ac_int_cctor_2_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11033" *)
  wire [32:0] alu_loop_op_else_else_else_else_ac_int_cctor_3_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11036" *)
  wire [32:0] alu_loop_op_else_else_else_else_ac_int_cctor_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11113" *)
  wire alu_loop_op_else_else_if_and_1_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11112" *)
  wire alu_loop_op_else_else_if_and_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10786" *)
  wire alu_loop_op_else_equal_tmp_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11738" *)
  wire [31:0] alu_loop_op_else_if_mux_10_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11739" *)
  wire [31:0] alu_loop_op_else_if_mux_11_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11730" *)
  wire [31:0] alu_loop_op_else_if_mux_12_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11731" *)
  wire [31:0] alu_loop_op_else_if_mux_13_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11734" *)
  wire [31:0] alu_loop_op_else_if_mux_14_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11735" *)
  wire [31:0] alu_loop_op_else_if_mux_15_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11726" *)
  wire [31:0] alu_loop_op_else_if_mux_8_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11727" *)
  wire [31:0] alu_loop_op_else_if_mux_9_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11026" *)
  wire [31:0] alu_loop_op_else_if_qr_31_0_1_lpi_1_dfm_mx0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11029" *)
  wire [31:0] alu_loop_op_else_if_qr_31_0_2_lpi_1_dfm_mx0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11032" *)
  wire [31:0] alu_loop_op_else_if_qr_31_0_3_lpi_1_dfm_mx0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11035" *)
  wire [31:0] alu_loop_op_else_if_qr_31_0_lpi_1_dfm_mx0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11551" *)
  wire alu_loop_op_else_mux_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11553" *)
  wire alu_loop_op_else_mux_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11561" *)
  wire alu_loop_op_else_mux_3_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11594" *)
  wire alu_loop_op_else_mux_4_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11592" *)
  wire alu_loop_op_else_mux_5_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11555" *)
  wire alu_loop_op_else_mux_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10992" *)
  wire alu_loop_op_else_nor_dfs;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10984" *)
  wire [31:0] alu_loop_op_else_o_32_1_1_lpi_1_dfm_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10985" *)
  wire [31:0] alu_loop_op_else_o_32_1_2_lpi_1_dfm_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10986" *)
  wire [31:0] alu_loop_op_else_o_32_1_3_lpi_1_dfm_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10987" *)
  wire [31:0] alu_loop_op_else_o_32_1_lpi_1_dfm_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10896" *)
  wire [31:0] alu_loop_op_else_o_mux1h_1_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10899" *)
  wire [31:0] alu_loop_op_else_o_mux1h_3_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10902" *)
  wire [31:0] alu_loop_op_else_o_mux1h_5_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10905" *)
  wire [31:0] alu_loop_op_else_o_mux1h_7_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10937" *)
  wire alu_loop_op_mux_204_mx1w1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11171" *)
  wire alu_loop_op_mux_209_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11186" *)
  wire alu_loop_op_mux_210_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11201" *)
  wire alu_loop_op_mux_212_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10576" *)
  reg alu_loop_op_unequal_tmp_6;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10577" *)
  reg alu_loop_op_unequal_tmp_7;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10578" *)
  reg alu_loop_op_unequal_tmp_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10867" *)
  wire and_167_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11325" *)
  wire and_192_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11346" *)
  wire and_196_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11355" *)
  wire and_200_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11364" *)
  wire and_204_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10869" *)
  wire and_211_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10870" *)
  wire and_213_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10871" *)
  wire and_215_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10872" *)
  wire and_217_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11407" *)
  wire and_218_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11408" *)
  wire and_220_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10873" *)
  wire and_231_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10874" *)
  wire and_233_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10875" *)
  wire and_235_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10876" *)
  wire and_237_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10877" *)
  wire and_239_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10878" *)
  wire and_241_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10879" *)
  wire and_243_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10880" *)
  wire and_245_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10882" *)
  wire and_293_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10808" *)
  wire and_297_m1c;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10883" *)
  wire and_328_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11793" *)
  wire and_336_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11797" *)
  wire and_338_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11801" *)
  wire and_340_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10777" *)
  wire and_357_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10855" *)
  wire and_37_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11790" *)
  wire and_443_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11782" *)
  wire and_444_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11771" *)
  wire and_446_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10831" *)
  wire and_451_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11860" *)
  wire and_474_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11545" *)
  wire and_478_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10851" *)
  wire and_481_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10842" *)
  wire and_484_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11534" *)
  wire and_485_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10829" *)
  wire and_486_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10860" *)
  wire and_489_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11426" *)
  wire and_493_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11423" *)
  wire and_494_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11420" *)
  wire and_495_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11417" *)
  wire and_496_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11291" *)
  wire and_497_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11280" *)
  wire and_498_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11268" *)
  wire and_499_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11256" *)
  wire and_500_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10852" *)
  wire and_501_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11204" *)
  wire and_502_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10861" *)
  wire and_524_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11090" *)
  wire and_550_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11080" *)
  wire and_564_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11414" *)
  wire and_729_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11136" *)
  wire and_734_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11604" *)
  wire and_74_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11086" *)
  wire and_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10868" *)
  wire and_dcpl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10439" *)
  wire and_dcpl_108;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10443" *)
  wire and_dcpl_127;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10454" *)
  wire and_dcpl_165;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10455" *)
  wire and_dcpl_167;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10456" *)
  wire and_dcpl_168;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10457" *)
  wire and_dcpl_169;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10458" *)
  wire and_dcpl_170;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10459" *)
  wire and_dcpl_171;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10462" *)
  wire and_dcpl_175;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10463" *)
  wire and_dcpl_179;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10350" *)
  wire and_dcpl_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10464" *)
  wire and_dcpl_207;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10465" *)
  wire and_dcpl_208;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10467" *)
  wire and_dcpl_214;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10468" *)
  wire and_dcpl_217;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10469" *)
  wire and_dcpl_219;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10470" *)
  wire and_dcpl_222;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10471" *)
  wire and_dcpl_225;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10473" *)
  wire and_dcpl_227;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10474" *)
  wire and_dcpl_229;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10475" *)
  wire and_dcpl_231;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10476" *)
  wire and_dcpl_234;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10477" *)
  wire and_dcpl_236;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10478" *)
  wire and_dcpl_239;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10479" *)
  wire and_dcpl_243;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10862" *)
  wire and_dcpl_269;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10413" *)
  wire and_dcpl_28;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10351" *)
  wire and_dcpl_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10414" *)
  wire and_dcpl_30;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10415" *)
  wire and_dcpl_32;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10416" *)
  wire and_dcpl_33;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10417" *)
  wire and_dcpl_34;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10881" *)
  wire and_dcpl_349;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10419" *)
  wire and_dcpl_35;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10420" *)
  wire and_dcpl_37;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10352" *)
  wire and_dcpl_4;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10421" *)
  wire and_dcpl_40;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10423" *)
  wire and_dcpl_43;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10424" *)
  wire and_dcpl_45;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10425" *)
  wire and_dcpl_46;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10426" *)
  wire and_dcpl_53;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10427" *)
  wire and_dcpl_64;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10428" *)
  wire and_dcpl_70;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10431" *)
  wire and_dcpl_77;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10432" *)
  wire and_dcpl_78;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10433" *)
  wire and_dcpl_80;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10434" *)
  wire and_dcpl_81;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10435" *)
  wire and_dcpl_83;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10436" *)
  wire and_dcpl_89;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10437" *)
  wire and_dcpl_96;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10438" *)
  wire and_dcpl_99;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10353" *)
  wire and_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10410" *)
  wire and_tmp_35;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10863" *)
  wire asn_267;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10592" *)
  reg [1:0] cfg_alu_algo_1_sva_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10624" *)
  reg [1:0] cfg_alu_algo_1_sva_st;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10682" *)
  reg [1:0] cfg_alu_algo_1_sva_st_20;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10717" *)
  reg [1:0] cfg_alu_algo_1_sva_st_22;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10719" *)
  reg [1:0] cfg_alu_algo_1_sva_st_23;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10721" *)
  reg [1:0] cfg_alu_algo_1_sva_st_24;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10724" *)
  reg [1:0] cfg_alu_algo_1_sva_st_25;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10744" *)
  reg [1:0] cfg_alu_algo_1_sva_st_28;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11138" *)
  wire [1:0] cfg_alu_algo_cfg_alu_algo_mux_3_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11069" *)
  wire cfg_alu_algo_cfg_alu_algo_or_3_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10281" *)
  output cfg_alu_algo_rsc_triosy_lz;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10320" *)
  wire cfg_alu_algo_rsc_triosy_obj_bawt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10299" *)
  input cfg_alu_algo_rsc_triosy_obj_oswt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10293" *)
  input [1:0] cfg_alu_algo_rsci_d;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10278" *)
  output cfg_alu_bypass_rsc_triosy_lz;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10317" *)
  wire cfg_alu_bypass_rsc_triosy_obj_bawt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10296" *)
  input cfg_alu_bypass_rsc_triosy_obj_oswt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10300" *)
  output cfg_alu_bypass_rsc_triosy_obj_oswt_unreg_pff;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10290" *)
  input cfg_alu_bypass_rsci_d;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10591" *)
  reg [31:0] cfg_alu_op_1_sva_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10280" *)
  output cfg_alu_op_rsc_triosy_lz;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10319" *)
  wire cfg_alu_op_rsc_triosy_obj_bawt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10298" *)
  input cfg_alu_op_rsc_triosy_obj_oswt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10292" *)
  input [31:0] cfg_alu_op_rsci_d;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10623" *)
  reg cfg_alu_src_1_sva_st;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10716" *)
  reg cfg_alu_src_1_sva_st_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10943" *)
  wire cfg_alu_src_1_sva_st_1_mx0c1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10279" *)
  output cfg_alu_src_rsc_triosy_lz;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10318" *)
  wire cfg_alu_src_rsc_triosy_obj_bawt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10297" *)
  input cfg_alu_src_rsc_triosy_obj_oswt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10291" *)
  input cfg_alu_src_rsci_d;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10282" *)
  input [1:0] cfg_precision;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10274" *)
  output chn_alu_in_rsc_lz;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10273" *)
  input chn_alu_in_rsc_vz;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10272" *)
  input [127:0] chn_alu_in_rsc_z;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10304" *)
  wire chn_alu_in_rsci_bawt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10307" *)
  wire [127:0] chn_alu_in_rsci_d_mxwt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10303" *)
  reg chn_alu_in_rsci_iswt0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10306" *)
  reg chn_alu_in_rsci_ld_core_psct;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10936" *)
  wire chn_alu_in_rsci_ld_core_psct_mx0c0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10286" *)
  input chn_alu_in_rsci_oswt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10287" *)
  output chn_alu_in_rsci_oswt_unreg;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10305" *)
  wire chn_alu_in_rsci_wen_comp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10277" *)
  output chn_alu_op_rsc_lz;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10276" *)
  input chn_alu_op_rsc_vz;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10275" *)
  input [127:0] chn_alu_op_rsc_z;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10310" *)
  wire chn_alu_op_rsci_bawt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10313" *)
  wire [127:0] chn_alu_op_rsci_d_mxwt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10309" *)
  reg chn_alu_op_rsci_iswt0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10312" *)
  reg chn_alu_op_rsci_ld_core_psct;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10940" *)
  wire chn_alu_op_rsci_ld_core_psct_mx0c1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10288" *)
  input chn_alu_op_rsci_oswt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10289" *)
  output chn_alu_op_rsci_oswt_unreg;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10311" *)
  wire chn_alu_op_rsci_wen_comp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11068" *)
  wire chn_alu_out_and_18_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10809" *)
  wire chn_alu_out_and_1_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10811" *)
  wire chn_alu_out_and_8_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10810" *)
  wire chn_alu_out_and_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11067" *)
  wire chn_alu_out_or_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10285" *)
  output chn_alu_out_rsc_lz;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10284" *)
  input chn_alu_out_rsc_vz;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10283" *)
  output [127:0] chn_alu_out_rsc_z;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10315" *)
  wire chn_alu_out_rsci_bawt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10336" *)
  reg chn_alu_out_rsci_d_0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10323" *)
  reg [21:0] chn_alu_out_rsci_d_118_97;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10322" *)
  reg [7:0] chn_alu_out_rsci_d_126_119;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10321" *)
  reg chn_alu_out_rsci_d_127;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10335" *)
  reg [21:0] chn_alu_out_rsci_d_22_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10334" *)
  reg [7:0] chn_alu_out_rsci_d_30_23;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10333" *)
  reg chn_alu_out_rsci_d_31;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10332" *)
  reg chn_alu_out_rsci_d_32;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10331" *)
  reg [21:0] chn_alu_out_rsci_d_54_33;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10330" *)
  reg [7:0] chn_alu_out_rsci_d_62_55;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10329" *)
  reg chn_alu_out_rsci_d_63;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10328" *)
  reg chn_alu_out_rsci_d_64;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10327" *)
  reg [21:0] chn_alu_out_rsci_d_86_65;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10326" *)
  reg [7:0] chn_alu_out_rsci_d_94_87;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10325" *)
  reg chn_alu_out_rsci_d_95;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10324" *)
  reg chn_alu_out_rsci_d_96;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10314" *)
  reg chn_alu_out_rsci_iswt0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10294" *)
  input chn_alu_out_rsci_oswt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10295" *)
  output chn_alu_out_rsci_oswt_unreg;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10316" *)
  wire chn_alu_out_rsci_wen_comp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10302" *)
  wire core_wen;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10308" *)
  wire core_wten;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10745" *)
  reg [30:0] else_AluOp_data_0_lpi_1_dfm_2_30_0_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10805" *)
  wire [31:0] else_AluOp_data_0_lpi_1_dfm_mx0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11059" *)
  wire [7:0] else_AluOp_data_0_lpi_1_dfm_mx1_tmp_30_23;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10807" *)
  wire [30:0] else_AluOp_data_0_lpi_1_dfm_mx3_30_0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10747" *)
  reg [30:0] else_AluOp_data_1_lpi_1_dfm_2_30_0_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10804" *)
  wire [31:0] else_AluOp_data_1_lpi_1_dfm_mx0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11060" *)
  wire [7:0] else_AluOp_data_1_lpi_1_dfm_mx1_tmp_30_23;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11061" *)
  wire [30:0] else_AluOp_data_1_lpi_1_dfm_mx2_30_0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10746" *)
  reg [30:0] else_AluOp_data_2_lpi_1_dfm_2_30_0_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10803" *)
  wire [31:0] else_AluOp_data_2_lpi_1_dfm_mx0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11062" *)
  wire [7:0] else_AluOp_data_2_lpi_1_dfm_mx1_tmp_30_23;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10806" *)
  wire [30:0] else_AluOp_data_2_lpi_1_dfm_mx3_30_0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10772" *)
  reg [30:0] else_AluOp_data_3_lpi_1_dfm_2_30_0_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10802" *)
  wire [31:0] else_AluOp_data_3_lpi_1_dfm_mx0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11058" *)
  wire [7:0] else_AluOp_data_3_lpi_1_dfm_mx1_tmp_30_23;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11073" *)
  wire else_AluOp_data_and_10_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11359" *)
  wire [22:0] else_AluOp_data_else_AluOp_data_mux_4_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11350" *)
  wire [22:0] else_AluOp_data_else_AluOp_data_mux_5_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11341" *)
  wire [22:0] else_AluOp_data_else_AluOp_data_mux_6_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11320" *)
  wire [22:0] else_AluOp_data_else_AluOp_data_mux_7_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10634" *)
  reg [22:0] else_AluOp_data_slc_else_AluOp_data_0_22_0_2_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10635" *)
  reg [22:0] else_AluOp_data_slc_else_AluOp_data_0_22_0_2_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10689" *)
  reg [7:0] else_AluOp_data_slc_else_AluOp_data_0_30_23_7_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10690" *)
  reg [7:0] else_AluOp_data_slc_else_AluOp_data_0_30_23_7_itm_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10646" *)
  reg [22:0] else_AluOp_data_slc_else_AluOp_data_1_22_0_7_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10647" *)
  reg [22:0] else_AluOp_data_slc_else_AluOp_data_1_22_0_7_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10691" *)
  reg [7:0] else_AluOp_data_slc_else_AluOp_data_1_30_23_21_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10692" *)
  reg [7:0] else_AluOp_data_slc_else_AluOp_data_1_30_23_21_itm_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10659" *)
  reg [22:0] else_AluOp_data_slc_else_AluOp_data_2_22_0_7_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10660" *)
  reg [22:0] else_AluOp_data_slc_else_AluOp_data_2_22_0_7_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10693" *)
  reg [7:0] else_AluOp_data_slc_else_AluOp_data_2_30_23_21_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10694" *)
  reg [7:0] else_AluOp_data_slc_else_AluOp_data_2_30_23_21_itm_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10672" *)
  reg [22:0] else_AluOp_data_slc_else_AluOp_data_3_22_0_12_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10673" *)
  reg [22:0] else_AluOp_data_slc_else_AluOp_data_3_22_0_12_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10687" *)
  reg [7:0] else_AluOp_data_slc_else_AluOp_data_3_30_23_35_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10688" *)
  reg [7:0] else_AluOp_data_slc_else_AluOp_data_3_30_23_35_itm_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11823" *)
  wire [22:0] else_else_mux_13_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10775" *)
  wire [8:0] else_mux_1_tmp_31_23;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10774" *)
  wire [8:0] else_mux_2_tmp_31_23;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10773" *)
  wire [8:0] else_mux_3_tmp_31_23;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10776" *)
  wire [8:0] else_mux_tmp_31_23;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10337" *)
  wire [1:0] fsm_output;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10595" *)
  reg io_read_cfg_alu_bypass_rsc_svs_5;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10596" *)
  reg io_read_cfg_alu_bypass_rsc_svs_6;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10597" *)
  reg io_read_cfg_alu_bypass_rsc_svs_7;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10598" *)
  reg io_read_cfg_alu_bypass_rsc_svs_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10715" *)
  reg io_read_cfg_alu_bypass_rsc_svs_st_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10718" *)
  reg io_read_cfg_alu_bypass_rsc_svs_st_5;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10720" *)
  reg io_read_cfg_alu_bypass_rsc_svs_st_6;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10723" *)
  reg io_read_cfg_alu_bypass_rsc_svs_st_7;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11063" *)
  wire [5:0] libraries_leading_sign_49_0_78e877fc94067377fcee479dbb0ed8e083a3_4;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11064" *)
  wire [5:0] libraries_leading_sign_49_0_78e877fc94067377fcee479dbb0ed8e083a3_5;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11065" *)
  wire [5:0] libraries_leading_sign_49_0_78e877fc94067377fcee479dbb0ed8e083a3_6;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11066" *)
  wire [5:0] libraries_leading_sign_49_0_78e877fc94067377fcee479dbb0ed8e083a3_7;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10778" *)
  wire main_stage_en_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10508" *)
  reg main_stage_v_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10942" *)
  wire main_stage_v_1_mx0c1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10509" *)
  reg main_stage_v_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10944" *)
  wire main_stage_v_2_mx0c1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10510" *)
  reg main_stage_v_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10961" *)
  wire main_stage_v_3_mx0c1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10511" *)
  reg main_stage_v_4;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10966" *)
  wire main_stage_v_4_mx0c1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11315" *)
  wire mux_100_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11330" *)
  wire mux_105_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11334" *)
  wire mux_106_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11329" *)
  wire mux_107_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11841" *)
  wire mux_108_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10913" *)
  wire mux_109_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11339" *)
  wire mux_110_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11337" *)
  wire mux_111_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11368" *)
  wire mux_124_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11371" *)
  wire mux_125_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11370" *)
  wire mux_126_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11377" *)
  wire mux_127_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11379" *)
  wire mux_128_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11382" *)
  wire mux_129_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11384" *)
  wire mux_130_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11387" *)
  wire mux_131_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11391" *)
  wire mux_132_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11390" *)
  wire mux_133_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11395" *)
  wire mux_134_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11394" *)
  wire mux_135_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11398" *)
  wire mux_136_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11400" *)
  wire mux_137_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11403" *)
  wire mux_138_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11404" *)
  wire mux_139_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11405" *)
  wire mux_140_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11843" *)
  wire mux_141_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11845" *)
  wire mux_142_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10914" *)
  wire mux_143_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11406" *)
  wire mux_144_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11415" *)
  wire mux_145_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11418" *)
  wire mux_146_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11421" *)
  wire mux_147_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11424" *)
  wire mux_148_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11428" *)
  wire mux_149_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11427" *)
  wire mux_150_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11432" *)
  wire mux_151_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11431" *)
  wire mux_152_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11436" *)
  wire mux_153_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11435" *)
  wire mux_154_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11440" *)
  wire mux_155_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11439" *)
  wire mux_156_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11443" *)
  wire mux_157_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11446" *)
  wire mux_158_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11449" *)
  wire mux_159_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11202" *)
  wire mux_15_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11452" *)
  wire mux_160_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11848" *)
  wire mux_162_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11850" *)
  wire mux_163_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11458" *)
  wire mux_164_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11459" *)
  wire mux_165_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11457" *)
  wire mux_166_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11456" *)
  wire mux_167_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11455" *)
  wire mux_168_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11828" *)
  wire mux_16_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11462" *)
  wire mux_171_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11461" *)
  wire mux_172_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11603" *)
  wire mux_173_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11602" *)
  wire mux_174_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11601" *)
  wire mux_175_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11465" *)
  wire mux_176_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10711" *)
  reg mux_177_itm_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10712" *)
  reg mux_177_itm_4;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11464" *)
  wire mux_177_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11852" *)
  wire mux_178_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10705" *)
  reg mux_181_itm_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10706" *)
  reg mux_181_itm_4;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11470" *)
  wire mux_181_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11469" *)
  wire mux_182_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11474" *)
  wire mux_183_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11473" *)
  wire mux_184_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11856" *)
  wire mux_185_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11858" *)
  wire mux_187_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10699" *)
  reg mux_189_itm_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10700" *)
  reg mux_189_itm_4;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11480" *)
  wire mux_189_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11208" *)
  wire mux_18_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11479" *)
  wire mux_190_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11484" *)
  wire mux_191_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11483" *)
  wire mux_192_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11489" *)
  wire mux_193_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11487" *)
  wire mux_194_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11492" *)
  wire mux_195_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11491" *)
  wire mux_196_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11496" *)
  wire mux_197_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11495" *)
  wire mux_198_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11500" *)
  wire mux_199_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11207" *)
  wire mux_19_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11499" *)
  wire mux_200_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11504" *)
  wire mux_201_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11503" *)
  wire mux_202_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11507" *)
  wire mux_203_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11506" *)
  wire mux_204_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11511" *)
  wire mux_205_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11510" *)
  wire mux_206_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11515" *)
  wire mux_207_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11514" *)
  wire mux_208_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11520" *)
  wire mux_209_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11210" *)
  wire mux_20_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11523" *)
  wire mux_210_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11526" *)
  wire mux_211_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11529" *)
  wire mux_212_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11533" *)
  wire mux_213_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11532" *)
  wire mux_214_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11536" *)
  wire mux_215_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11535" *)
  wire mux_216_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11537" *)
  wire mux_217_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11540" *)
  wire mux_218_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11542" *)
  wire mux_219_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11209" *)
  wire mux_21_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11546" *)
  wire mux_221_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11544" *)
  wire mux_222_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11562" *)
  wire mux_223_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11564" *)
  wire mux_224_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11566" *)
  wire mux_225_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11568" *)
  wire mux_226_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11206" *)
  wire mux_22_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11859" *)
  wire mux_233_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11205" *)
  wire mux_23_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11584" *)
  wire mux_243_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11586" *)
  wire mux_244_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11585" *)
  wire mux_245_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11583" *)
  wire mux_246_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11582" *)
  wire mux_247_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11865" *)
  wire mux_248_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11870" *)
  wire mux_249_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11830" *)
  wire mux_24_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11868" *)
  wire mux_250_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11863" *)
  wire mux_251_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11867" *)
  wire mux_253_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11864" *)
  wire mux_254_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11872" *)
  wire mux_255_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11877" *)
  wire mux_256_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11876" *)
  wire mux_257_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11875" *)
  wire mux_258_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11874" *)
  wire mux_259_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11871" *)
  wire mux_260_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11608" *)
  wire mux_262_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11610" *)
  wire mux_263_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11613" *)
  wire mux_264_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11614" *)
  wire mux_265_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11612" *)
  wire mux_266_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11611" *)
  wire mux_267_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11609" *)
  wire mux_268_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11607" *)
  wire mux_269_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11214" *)
  wire mux_26_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11606" *)
  wire mux_270_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11617" *)
  wire mux_271_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11619" *)
  wire mux_272_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11621" *)
  wire mux_273_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11620" *)
  wire mux_274_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11618" *)
  wire mux_275_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11616" *)
  wire mux_276_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11615" *)
  wire mux_277_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11879" *)
  wire mux_279_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11213" *)
  wire mux_27_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11165" *)
  wire mux_281_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10844" *)
  wire mux_282_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11628" *)
  wire mux_284_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11627" *)
  wire mux_285_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11626" *)
  wire mux_286_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11630" *)
  wire mux_287_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11625" *)
  wire mux_288_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11633" *)
  wire mux_289_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11216" *)
  wire mux_28_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11624" *)
  wire mux_290_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11638" *)
  wire mux_297_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11637" *)
  wire mux_298_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11636" *)
  wire mux_299_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11215" *)
  wire mux_29_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11640" *)
  wire mux_300_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11635" *)
  wire mux_301_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11643" *)
  wire mux_302_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11634" *)
  wire mux_303_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11645" *)
  wire mux_304_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11644" *)
  wire mux_305_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11647" *)
  wire mux_306_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11646" *)
  wire mux_307_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11212" *)
  wire mux_30_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11883" *)
  wire mux_310_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10843" *)
  wire mux_312_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11649" *)
  wire mux_313_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11648" *)
  wire mux_314_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11211" *)
  wire mux_31_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11328" *)
  wire mux_327_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11326" *)
  wire mux_328_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11349" *)
  wire mux_329_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11833" *)
  wire mux_32_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11347" *)
  wire mux_330_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11358" *)
  wire mux_331_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11356" *)
  wire mux_332_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11367" *)
  wire mux_333_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11365" *)
  wire mux_334_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10915" *)
  wire mux_337_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11769" *)
  wire mux_339_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11832" *)
  wire mux_33_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11773" *)
  wire mux_340_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11780" *)
  wire mux_341_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11788" *)
  wire mux_342_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11792" *)
  wire mux_343_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11796" *)
  wire mux_344_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11800" *)
  wire mux_345_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10912" *)
  wire mux_34_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11221" *)
  wire mux_35_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11410" *)
  wire mux_361_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11409" *)
  wire mux_362_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11570" *)
  wire mux_363_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11571" *)
  wire mux_364_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11572" *)
  wire mux_365_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11574" *)
  wire mux_366_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11220" *)
  wire mux_36_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11218" *)
  wire mux_37_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11374" *)
  wire mux_383_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11217" *)
  wire mux_38_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11223" *)
  wire mux_43_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11229" *)
  wire mux_44_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11228" *)
  wire mux_45_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11227" *)
  wire mux_46_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11838" *)
  wire mux_56_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11231" *)
  wire mux_58_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11230" *)
  wire mux_59_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11236" *)
  wire mux_60_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11235" *)
  wire mux_61_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11241" *)
  wire mux_62_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11240" *)
  wire mux_63_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11246" *)
  wire mux_64_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11245" *)
  wire mux_65_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11252" *)
  wire mux_66_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11250" *)
  wire mux_67_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11257" *)
  wire mux_69_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11255" *)
  wire mux_70_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11262" *)
  wire mux_73_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11253" *)
  wire mux_74_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11269" *)
  wire mux_75_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11267" *)
  wire mux_76_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11274" *)
  wire mux_79_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11265" *)
  wire mux_80_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11281" *)
  wire mux_81_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11279" *)
  wire mux_82_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11286" *)
  wire mux_85_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11277" *)
  wire mux_86_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11292" *)
  wire mux_87_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11290" *)
  wire mux_88_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11297" *)
  wire mux_91_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11289" *)
  wire mux_92_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11301" *)
  wire mux_93_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11300" *)
  wire mux_94_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11306" *)
  wire mux_95_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11305" *)
  wire mux_96_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11311" *)
  wire mux_97_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11310" *)
  wire mux_98_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11316" *)
  wire mux_99_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11412" *)
  wire mux_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11126" *)
  wire mux_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10357" *)
  wire mux_tmp_10;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10380" *)
  wire mux_tmp_146;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10387" *)
  wire mux_tmp_164;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10388" *)
  wire mux_tmp_165;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10390" *)
  wire mux_tmp_171;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10392" *)
  wire mux_tmp_173;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10355" *)
  wire mux_tmp_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10396" *)
  wire mux_tmp_227;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10399" *)
  wire mux_tmp_237;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10401" *)
  wire mux_tmp_246;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10406" *)
  wire mux_tmp_265;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10407" *)
  wire mux_tmp_268;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10408" *)
  wire mux_tmp_281;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10411" *)
  wire mux_tmp_296;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10441" *)
  wire mux_tmp_311;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10466" *)
  wire mux_tmp_323;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11127" *)
  wire mux_tmp_348;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11128" *)
  wire mux_tmp_349;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11129" *)
  wire mux_tmp_350;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10366" *)
  wire mux_tmp_53;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11078" *)
  wire nand_109_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11834" *)
  wire nand_17_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11219" *)
  wire nand_18_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11460" *)
  wire nand_29_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11605" *)
  wire nand_30_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11629" *)
  wire nand_35_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11632" *)
  wire nand_36_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11639" *)
  wire nand_37_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11642" *)
  wire nand_38_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11203" *)
  wire nand_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10381" *)
  wire nand_tmp_13;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10400" *)
  wire nand_tmp_20;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11888" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 24 25" *)
  wire [25:0] nl_FpAdd_8U_23U_is_a_greater_oif_aelse_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11890" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 24 25" *)
  wire [25:0] nl_FpAdd_8U_23U_is_a_greater_oif_aelse_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11892" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 24 25" *)
  wire [25:0] nl_FpAdd_8U_23U_is_a_greater_oif_aelse_acc_3_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11886" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 24 25" *)
  wire [25:0] nl_FpAdd_8U_23U_is_a_greater_oif_aelse_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11786" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 9 10" *)
  wire [10:0] nl_FpCmp_8U_23U_false_else_if_acc_10_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11765" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 9 10" *)
  wire [10:0] nl_FpCmp_8U_23U_false_else_if_acc_4_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11820" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 9 10" *)
  wire [10:0] nl_FpCmp_8U_23U_false_else_if_acc_6_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11778" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 9 10" *)
  wire [10:0] nl_FpCmp_8U_23U_false_else_if_acc_8_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11822" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 24 25" *)
  wire [25:0] nl_FpCmp_8U_23U_true_else_else_if_acc_4_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11784" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 24 25" *)
  wire [25:0] nl_FpCmp_8U_23U_true_else_else_if_acc_6_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11776" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 24 25" *)
  wire [25:0] nl_FpCmp_8U_23U_true_else_else_if_acc_7_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11767" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 24 25" *)
  wire [25:0] nl_FpCmp_8U_23U_true_else_else_if_acc_8_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11827" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 9 10" *)
  wire [10:0] nl_FpCmp_8U_23U_true_if_acc_10_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11816" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 9 10" *)
  wire [10:0] nl_FpCmp_8U_23U_true_if_acc_4_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11818" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 9 10" *)
  wire [10:0] nl_FpCmp_8U_23U_true_if_acc_6_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11825" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 9 10" *)
  wire [10:0] nl_FpCmp_8U_23U_true_if_acc_8_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12030" *)
  wire [127:0] nl_Y_alu_core_chn_alu_out_rsci_inst_chn_alu_out_rsci_d;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11729" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31 32 34" *)
  wire [34:0] nl_acc_10_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11733" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31 32 34" *)
  wire [34:0] nl_acc_11_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11910" *)
  (* unused_bits = "0 51" *)
  wire [51:0] nl_acc_12_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11914" *)
  (* unused_bits = "0 51" *)
  wire [51:0] nl_acc_13_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11918" *)
  (* unused_bits = "0 51" *)
  wire [51:0] nl_acc_14_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11922" *)
  (* unused_bits = "0 51" *)
  wire [51:0] nl_acc_15_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11674" *)
  (* unused_bits = "0 9" *)
  wire [9:0] nl_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11678" *)
  (* unused_bits = "0 9" *)
  wire [9:0] nl_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11682" *)
  (* unused_bits = "0 9" *)
  wire [9:0] nl_acc_3_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11894" *)
  (* unused_bits = "0 9" *)
  wire [9:0] nl_acc_4_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11898" *)
  (* unused_bits = "0 9" *)
  wire [9:0] nl_acc_5_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11902" *)
  (* unused_bits = "0 9" *)
  wire [9:0] nl_acc_6_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11906" *)
  (* unused_bits = "0 9" *)
  wire [9:0] nl_acc_7_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11725" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31 32 34" *)
  wire [34:0] nl_acc_8_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11737" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31 32 34" *)
  wire [34:0] nl_acc_9_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11670" *)
  (* unused_bits = "0 9" *)
  wire [9:0] nl_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12003" *)
  wire [23:0] nl_alu_loop_op_1_FpAdd_8U_23U_a_int_mant_p1_lshift_rg_a;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12008" *)
  wire [8:0] nl_alu_loop_op_1_FpAdd_8U_23U_a_int_mant_p1_lshift_rg_s;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12007" *)
  (* unused_bits = "8" *)
  wire [8:0] nl_alu_loop_op_1_FpAdd_8U_23U_a_left_shift_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11926" *)
  wire [23:0] nl_alu_loop_op_1_FpAdd_8U_23U_b_int_mant_p1_lshift_rg_a;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11931" *)
  wire [8:0] nl_alu_loop_op_1_FpAdd_8U_23U_b_int_mant_p1_lshift_rg_s;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11930" *)
  (* unused_bits = "8" *)
  wire [8:0] nl_alu_loop_op_1_FpAdd_8U_23U_b_left_shift_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11702" *)
  (* unused_bits = "0 1 2 3 4 5 6 8" *)
  wire [8:0] nl_alu_loop_op_1_FpAdd_8U_23U_if_3_if_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11741" *)
  (* unused_bits = "0 1 2 3 4 5 6 8" *)
  wire [8:0] nl_alu_loop_op_1_FpAdd_8U_23U_if_4_if_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11179" *)
  (* unused_bits = "8" *)
  wire [8:0] nl_alu_loop_op_1_FpAdd_8U_23U_if_4_if_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11362" *)
  (* unused_bits = "23" *)
  wire [23:0] nl_alu_loop_op_1_FpMantRNE_49U_24U_else_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11808" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 9 10" *)
  wire [10:0] nl_alu_loop_op_1_FpNormalize_8U_49U_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12028" *)
  wire [48:0] nl_alu_loop_op_1_FpNormalize_8U_49U_else_lshift_rg_a;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11757" *)
  (* unused_bits = "0 1 3" *)
  wire [3:0] nl_alu_loop_op_1_IntSaturation_33U_32U_else_if_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11700" *)
  (* unused_bits = "0 1 3" *)
  wire [3:0] nl_alu_loop_op_1_IntSaturation_33U_32U_if_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12014" *)
  wire [48:0] nl_alu_loop_op_1_leading_sign_49_0_rg_mantissa;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11992" *)
  wire [23:0] nl_alu_loop_op_2_FpAdd_8U_23U_a_int_mant_p1_lshift_2_rg_a;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11997" *)
  wire [8:0] nl_alu_loop_op_2_FpAdd_8U_23U_a_int_mant_p1_lshift_2_rg_s;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11996" *)
  (* unused_bits = "8" *)
  wire [8:0] nl_alu_loop_op_2_FpAdd_8U_23U_a_left_shift_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11937" *)
  wire [23:0] nl_alu_loop_op_2_FpAdd_8U_23U_b_int_mant_p1_lshift_2_rg_a;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11942" *)
  wire [8:0] nl_alu_loop_op_2_FpAdd_8U_23U_b_int_mant_p1_lshift_2_rg_s;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11941" *)
  (* unused_bits = "8" *)
  wire [8:0] nl_alu_loop_op_2_FpAdd_8U_23U_b_left_shift_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11704" *)
  (* unused_bits = "0 1 2 3 4 5 6 8" *)
  wire [8:0] nl_alu_loop_op_2_FpAdd_8U_23U_if_3_if_acc_4_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11743" *)
  (* unused_bits = "0 1 2 3 4 5 6 8" *)
  wire [8:0] nl_alu_loop_op_2_FpAdd_8U_23U_if_4_if_acc_4_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11194" *)
  (* unused_bits = "8" *)
  wire [8:0] nl_alu_loop_op_2_FpAdd_8U_23U_if_4_if_acc_5_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11353" *)
  (* unused_bits = "23" *)
  wire [23:0] nl_alu_loop_op_2_FpMantRNE_49U_24U_else_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11810" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 9 10" *)
  wire [10:0] nl_alu_loop_op_2_FpNormalize_8U_49U_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12026" *)
  wire [48:0] nl_alu_loop_op_2_FpNormalize_8U_49U_else_lshift_2_rg_a;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11759" *)
  (* unused_bits = "0 1 3" *)
  wire [3:0] nl_alu_loop_op_2_IntSaturation_33U_32U_else_if_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11690" *)
  (* unused_bits = "0 1 3" *)
  wire [3:0] nl_alu_loop_op_2_IntSaturation_33U_32U_if_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12016" *)
  wire [48:0] nl_alu_loop_op_2_leading_sign_49_0_2_rg_mantissa;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11981" *)
  wire [23:0] nl_alu_loop_op_3_FpAdd_8U_23U_a_int_mant_p1_lshift_1_rg_a;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11986" *)
  wire [8:0] nl_alu_loop_op_3_FpAdd_8U_23U_a_int_mant_p1_lshift_1_rg_s;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11985" *)
  (* unused_bits = "8" *)
  wire [8:0] nl_alu_loop_op_3_FpAdd_8U_23U_a_left_shift_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11948" *)
  wire [23:0] nl_alu_loop_op_3_FpAdd_8U_23U_b_int_mant_p1_lshift_1_rg_a;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11953" *)
  wire [8:0] nl_alu_loop_op_3_FpAdd_8U_23U_b_int_mant_p1_lshift_1_rg_s;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11952" *)
  (* unused_bits = "8" *)
  wire [8:0] nl_alu_loop_op_3_FpAdd_8U_23U_b_left_shift_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11706" *)
  (* unused_bits = "0 1 2 3 4 5 6 8" *)
  wire [8:0] nl_alu_loop_op_3_FpAdd_8U_23U_if_3_if_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11745" *)
  (* unused_bits = "0 1 2 3 4 5 6 8" *)
  wire [8:0] nl_alu_loop_op_3_FpAdd_8U_23U_if_4_if_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11657" *)
  (* unused_bits = "8" *)
  wire [8:0] nl_alu_loop_op_3_FpAdd_8U_23U_if_4_if_acc_3_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11344" *)
  (* unused_bits = "23" *)
  wire [23:0] nl_alu_loop_op_3_FpMantRNE_49U_24U_else_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11812" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 9 10" *)
  wire [10:0] nl_alu_loop_op_3_FpNormalize_8U_49U_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12024" *)
  wire [48:0] nl_alu_loop_op_3_FpNormalize_8U_49U_else_lshift_1_rg_a;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11761" *)
  (* unused_bits = "0 1 3" *)
  wire [3:0] nl_alu_loop_op_3_IntSaturation_33U_32U_else_if_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11698" *)
  (* unused_bits = "0 1 3" *)
  wire [3:0] nl_alu_loop_op_3_IntSaturation_33U_32U_if_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12018" *)
  wire [48:0] nl_alu_loop_op_3_leading_sign_49_0_1_rg_mantissa;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11970" *)
  wire [23:0] nl_alu_loop_op_4_FpAdd_8U_23U_a_int_mant_p1_lshift_3_rg_a;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11975" *)
  wire [8:0] nl_alu_loop_op_4_FpAdd_8U_23U_a_int_mant_p1_lshift_3_rg_s;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11974" *)
  (* unused_bits = "8" *)
  wire [8:0] nl_alu_loop_op_4_FpAdd_8U_23U_a_left_shift_acc_3_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11959" *)
  wire [23:0] nl_alu_loop_op_4_FpAdd_8U_23U_b_int_mant_p1_lshift_3_rg_a;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11964" *)
  wire [8:0] nl_alu_loop_op_4_FpAdd_8U_23U_b_int_mant_p1_lshift_3_rg_s;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11963" *)
  (* unused_bits = "8" *)
  wire [8:0] nl_alu_loop_op_4_FpAdd_8U_23U_b_left_shift_acc_3_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11708" *)
  (* unused_bits = "0 1 2 3 4 5 6 8" *)
  wire [8:0] nl_alu_loop_op_4_FpAdd_8U_23U_if_3_if_acc_6_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11747" *)
  (* unused_bits = "0 1 2 3 4 5 6 8" *)
  wire [8:0] nl_alu_loop_op_4_FpAdd_8U_23U_if_4_if_acc_6_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11717" *)
  (* unused_bits = "8" *)
  wire [8:0] nl_alu_loop_op_4_FpAdd_8U_23U_if_4_if_acc_7_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11323" *)
  (* unused_bits = "23" *)
  wire [23:0] nl_alu_loop_op_4_FpMantRNE_49U_24U_else_acc_3_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11814" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 9 10" *)
  wire [10:0] nl_alu_loop_op_4_FpNormalize_8U_49U_acc_3_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12022" *)
  wire [48:0] nl_alu_loop_op_4_FpNormalize_8U_49U_else_lshift_3_rg_a;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11763" *)
  (* unused_bits = "0 1 3" *)
  wire [3:0] nl_alu_loop_op_4_IntSaturation_33U_32U_else_if_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11696" *)
  (* unused_bits = "0 1 3" *)
  wire [3:0] nl_alu_loop_op_4_IntSaturation_33U_32U_if_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12020" *)
  wire [48:0] nl_alu_loop_op_4_leading_sign_49_0_3_rg_mantissa;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11028" *)
  (* unused_bits = "33" *)
  wire [33:0] nl_alu_loop_op_else_else_else_else_ac_int_cctor_1_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11031" *)
  (* unused_bits = "33" *)
  wire [33:0] nl_alu_loop_op_else_else_else_else_ac_int_cctor_2_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11034" *)
  (* unused_bits = "33" *)
  wire [33:0] nl_alu_loop_op_else_else_else_else_ac_int_cctor_3_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11037" *)
  (* unused_bits = "33" *)
  wire [33:0] nl_alu_loop_op_else_else_else_else_ac_int_cctor_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11802" *)
  wire nor_156_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11798" *)
  wire nor_159_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11794" *)
  wire nor_162_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11789" *)
  wire nor_163_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11781" *)
  wire nor_165_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11770" *)
  wire nor_168_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11641" *)
  wire nor_176_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10853" *)
  wire nor_177_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11631" *)
  wire nor_178_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11861" *)
  wire nor_187_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11569" *)
  wire nor_192_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11567" *)
  wire nor_195_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10839" *)
  wire nor_197_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11565" *)
  wire nor_200_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10856" *)
  wire nor_201_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10826" *)
  wire nor_202_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11563" *)
  wire nor_203_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11547" *)
  wire nor_204_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11549" *)
  wire nor_205_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11543" *)
  wire nor_206_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11541" *)
  wire nor_207_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11538" *)
  wire nor_208_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11539" *)
  wire nor_210_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11530" *)
  wire nor_213_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11531" *)
  wire nor_214_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11527" *)
  wire nor_215_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11528" *)
  wire nor_216_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11524" *)
  wire nor_217_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11525" *)
  wire nor_218_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11521" *)
  wire nor_219_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11522" *)
  wire nor_220_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11516" *)
  wire nor_222_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11517" *)
  wire nor_223_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11512" *)
  wire nor_227_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11513" *)
  wire nor_228_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11508" *)
  wire nor_232_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11509" *)
  wire nor_233_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10821" *)
  wire nor_236_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11501" *)
  wire nor_237_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11502" *)
  wire nor_238_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11466" *)
  wire nor_241_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11467" *)
  wire nor_243_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11847" *)
  wire nor_248_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11453" *)
  wire nor_249_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11450" *)
  wire nor_250_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11447" *)
  wire nor_251_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11444" *)
  wire nor_252_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11441" *)
  wire nor_254_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11442" *)
  wire nor_256_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11437" *)
  wire nor_257_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11438" *)
  wire nor_259_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11433" *)
  wire nor_260_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11434" *)
  wire nor_262_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11429" *)
  wire nor_263_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10816" *)
  wire nor_264_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11430" *)
  wire nor_265_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11401" *)
  wire nor_267_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11402" *)
  wire nor_268_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10820" *)
  wire nor_269_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11388" *)
  wire nor_270_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11389" *)
  wire nor_271_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11385" *)
  wire nor_272_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11386" *)
  wire nor_273_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11380" *)
  wire nor_274_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11381" *)
  wire nor_275_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11331" *)
  wire nor_290_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11332" *)
  wire nor_291_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11333" *)
  wire nor_292_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11335" *)
  wire nor_293_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11317" *)
  wire nor_298_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11318" *)
  wire nor_299_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11319" *)
  wire nor_300_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11312" *)
  wire nor_301_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11313" *)
  wire nor_302_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11314" *)
  wire nor_303_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11307" *)
  wire nor_304_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11308" *)
  wire nor_305_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11309" *)
  wire nor_306_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11302" *)
  wire nor_307_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11303" *)
  wire nor_308_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11304" *)
  wire nor_309_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11293" *)
  wire nor_310_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11294" *)
  wire nor_311_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11295" *)
  wire nor_312_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11296" *)
  wire nor_313_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11278" *)
  wire nor_314_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11282" *)
  wire nor_316_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11283" *)
  wire nor_317_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11284" *)
  wire nor_318_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11285" *)
  wire nor_319_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11287" *)
  wire nor_320_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11288" *)
  wire nor_322_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11266" *)
  wire nor_324_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11270" *)
  wire nor_326_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11271" *)
  wire nor_327_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11272" *)
  wire nor_328_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11273" *)
  wire nor_329_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11275" *)
  wire nor_330_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11276" *)
  wire nor_332_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11254" *)
  wire nor_334_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11258" *)
  wire nor_336_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11259" *)
  wire nor_337_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11260" *)
  wire nor_338_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11261" *)
  wire nor_339_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10832" *)
  wire nor_33_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11263" *)
  wire nor_340_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11264" *)
  wire nor_342_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11251" *)
  wire nor_344_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11247" *)
  wire nor_345_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11248" *)
  wire nor_346_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11249" *)
  wire nor_347_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11242" *)
  wire nor_348_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11243" *)
  wire nor_349_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11244" *)
  wire nor_350_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11237" *)
  wire nor_351_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11238" *)
  wire nor_352_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11239" *)
  wire nor_353_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11232" *)
  wire nor_354_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11233" *)
  wire nor_355_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11234" *)
  wire nor_356_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11837" *)
  wire nor_357_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11224" *)
  wire nor_367_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11225" *)
  wire nor_368_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11835" *)
  wire nor_371_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11836" *)
  wire nor_372_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11851" *)
  wire nor_379_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10833" *)
  wire nor_37_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10858" *)
  wire nor_397_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11185" *)
  wire nor_406_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11200" *)
  wire nor_407_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11663" *)
  wire nor_408_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10834" *)
  wire nor_41_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11079" *)
  wire nor_430_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11684" *)
  wire nor_433_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11680" *)
  wire nor_434_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11676" *)
  wire nor_435_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11672" *)
  wire nor_436_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11135" *)
  wire nor_437_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10835" *)
  wire nor_45_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10854" *)
  wire nor_71_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10409" *)
  wire nor_tmp_126;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10442" *)
  wire nor_tmp_144;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10385" *)
  wire nor_tmp_74;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10379" *)
  wire not_tmp_152;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10382" *)
  wire not_tmp_157;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10394" *)
  wire not_tmp_232;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10359" *)
  wire not_tmp_24;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10402" *)
  wire not_tmp_259;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10405" *)
  wire not_tmp_261;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10361" *)
  wire not_tmp_29;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10362" *)
  wire not_tmp_38;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10364" *)
  wire not_tmp_57;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10270" *)
  input nvdla_core_clk;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10271" *)
  input nvdla_core_rstn;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11411" *)
  wire or_1046_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11413" *)
  wire or_1048_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11104" *)
  wire or_1050_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11105" *)
  wire or_1055_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11573" *)
  wire or_1069_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11575" *)
  wire or_1076_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11137" *)
  wire or_1087_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11375" *)
  wire or_1100_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11376" *)
  wire or_1106_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10857" *)
  wire or_16_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11298" *)
  wire or_182_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11336" *)
  wire or_225_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11840" *)
  wire or_230_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11842" *)
  wire or_233_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11340" *)
  wire or_236_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11338" *)
  wire or_239_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11369" *)
  wire or_270_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11372" *)
  wire or_273_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11373" *)
  wire or_275_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11378" *)
  wire or_280_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11383" *)
  wire or_288_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10846" *)
  wire or_28_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11392" *)
  wire or_299_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11393" *)
  wire or_301_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11396" *)
  wire or_304_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11397" *)
  wire or_307_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11399" *)
  wire or_312_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11844" *)
  wire or_323_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11416" *)
  wire or_333_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11419" *)
  wire or_334_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11422" *)
  wire or_335_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11425" *)
  wire or_336_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10841" *)
  wire or_381_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11849" *)
  wire or_383_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11846" *)
  wire or_386_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10840" *)
  wire or_391_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11463" *)
  wire or_400_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11853" *)
  wire or_417_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11854" *)
  wire or_419_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11472" *)
  wire or_420_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11471" *)
  wire or_422_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11475" *)
  wire or_426_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11855" *)
  wire or_428_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11857" *)
  wire or_432_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11481" *)
  wire or_438_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11222" *)
  wire or_43_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11482" *)
  wire or_440_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11485" *)
  wire or_441_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11486" *)
  wire or_443_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11490" *)
  wire or_444_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11488" *)
  wire or_446_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11493" *)
  wire or_450_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11497" *)
  wire or_453_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11505" *)
  wire or_463_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11866" *)
  wire or_601_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11869" *)
  wire or_607_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11862" *)
  wire or_609_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11873" *)
  wire or_610_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11878" *)
  wire or_612_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11623" *)
  wire or_619_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11622" *)
  wire or_624_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11880" *)
  wire or_629_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10845" *)
  wire or_632_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11327" *)
  wire or_735_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11348" *)
  wire or_741_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11357" *)
  wire or_744_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11366" *)
  wire or_747_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10836" *)
  wire or_861_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11774" *)
  wire or_864_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10837" *)
  wire or_867_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10838" *)
  wire or_871_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11791" *)
  wire or_876_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11839" *)
  wire or_87_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11795" *)
  wire or_880_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11799" *)
  wire or_884_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10827" *)
  wire or_937_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11454" *)
  wire or_958_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11451" *)
  wire or_959_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11448" *)
  wire or_960_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11445" *)
  wire or_961_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11299" *)
  wire or_962_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10824" *)
  wire or_963_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11831" *)
  wire or_965_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11829" *)
  wire or_967_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10865" *)
  wire or_996_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10864" *)
  wire or_997_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10866" *)
  wire or_998_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11125" *)
  wire or_dcpl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10448" *)
  wire or_dcpl_100;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10449" *)
  wire or_dcpl_109;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10450" *)
  wire or_dcpl_117;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10451" *)
  wire or_dcpl_119;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10452" *)
  wire or_dcpl_121;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10453" *)
  wire or_dcpl_123;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10460" *)
  wire or_dcpl_125;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10461" *)
  wire or_dcpl_127;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10412" *)
  wire or_dcpl_14;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10472" *)
  wire or_dcpl_154;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10418" *)
  wire or_dcpl_20;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10422" *)
  wire or_dcpl_23;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11130" *)
  wire or_dcpl_272;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10429" *)
  wire or_dcpl_46;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10430" *)
  wire or_dcpl_49;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10444" *)
  wire or_dcpl_85;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10445" *)
  wire or_dcpl_86;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10446" *)
  wire or_dcpl_89;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10447" *)
  wire or_dcpl_91;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10365" *)
  wire or_tmp_103;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10356" *)
  wire or_tmp_15;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10358" *)
  wire or_tmp_20;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10367" *)
  wire or_tmp_218;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10368" *)
  wire or_tmp_224;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10360" *)
  wire or_tmp_23;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10369" *)
  wire or_tmp_251;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10370" *)
  wire or_tmp_261;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10371" *)
  wire or_tmp_269;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10372" *)
  wire or_tmp_280;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10373" *)
  wire or_tmp_293;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10374" *)
  wire or_tmp_305;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10375" *)
  wire or_tmp_309;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10376" *)
  wire or_tmp_312;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10377" *)
  wire or_tmp_315;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10378" *)
  wire or_tmp_347;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10383" *)
  wire or_tmp_382;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10384" *)
  wire or_tmp_386;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10386" *)
  wire or_tmp_395;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10389" *)
  wire or_tmp_402;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10391" *)
  wire or_tmp_409;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10393" *)
  wire or_tmp_416;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10395" *)
  wire or_tmp_577;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10397" *)
  wire or_tmp_583;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10398" *)
  wire or_tmp_585;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10403" *)
  wire or_tmp_596;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10404" *)
  wire or_tmp_597;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10440" *)
  wire or_tmp_657;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10480" *)
  wire or_tmp_668;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10481" *)
  wire or_tmp_674;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10482" *)
  wire or_tmp_678;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10483" *)
  wire or_tmp_695;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10363" *)
  wire or_tmp_75;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10354" *)
  wire or_tmp_9;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10886" *)
  reg [22:0] reg_AluIn_data_sva_4_126_96_1_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10885" *)
  reg [7:0] reg_AluIn_data_sva_4_126_96_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10895" *)
  reg [22:0] reg_AluIn_data_sva_4_30_0_1_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10894" *)
  reg [7:0] reg_AluIn_data_sva_4_30_0_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10892" *)
  reg [22:0] reg_AluIn_data_sva_4_62_32_1_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10891" *)
  reg [7:0] reg_AluIn_data_sva_4_62_32_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10889" *)
  reg [22:0] reg_AluIn_data_sva_4_94_64_1_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10888" *)
  reg [7:0] reg_AluIn_data_sva_4_94_64_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11124" *)
  reg reg_alu_loop_op_1_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_1_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11123" *)
  reg reg_alu_loop_op_2_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_2_svs_1_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11122" *)
  reg reg_alu_loop_op_3_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_1_svs_1_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11070" *)
  reg reg_alu_loop_op_4_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_3_svs_1_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10898" *)
  reg [30:0] reg_alu_loop_op_else_o_32_1_1_lpi_1_dfm_3_1_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10897" *)
  reg reg_alu_loop_op_else_o_32_1_1_lpi_1_dfm_3_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10901" *)
  reg [30:0] reg_alu_loop_op_else_o_32_1_2_lpi_1_dfm_4_1_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10900" *)
  reg reg_alu_loop_op_else_o_32_1_2_lpi_1_dfm_4_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10904" *)
  reg [30:0] reg_alu_loop_op_else_o_32_1_3_lpi_1_dfm_3_1_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10903" *)
  reg reg_alu_loop_op_else_o_32_1_3_lpi_1_dfm_3_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10907" *)
  reg [30:0] reg_alu_loop_op_else_o_32_1_lpi_1_dfm_4_1_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10906" *)
  reg reg_alu_loop_op_else_o_32_1_lpi_1_dfm_4_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11114" *)
  reg [1:0] reg_cfg_alu_algo_1_sva_st_13_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10812" *)
  reg reg_cfg_alu_algo_rsc_triosy_obj_ld_core_psct_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10814" *)
  reg reg_chn_alu_out_rsci_ld_core_psct_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10929" *)
  wire [49:0] z_out_12;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10931" *)
  wire [49:0] z_out_13;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10933" *)
  wire [49:0] z_out_14;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10935" *)
  wire [49:0] z_out_15;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10921" *)
  wire [7:0] z_out_4;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10923" *)
  wire [7:0] z_out_5;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10925" *)
  wire [7:0] z_out_6;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10927" *)
  wire [7:0] z_out_7;
  assign alu_loop_op_1_FpAdd_8U_23U_b_left_shift_acc_nl = { 1'b1, _1174_ } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11933" *) 4'b1101;
  assign alu_loop_op_2_FpAdd_8U_23U_b_left_shift_acc_2_nl = { 1'b1, _1175_ } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11944" *) 4'b1101;
  assign alu_loop_op_3_FpAdd_8U_23U_b_left_shift_acc_1_nl = { 1'b1, _1176_ } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11955" *) 4'b1101;
  assign alu_loop_op_4_FpAdd_8U_23U_b_left_shift_acc_3_nl = { 1'b1, _1177_ } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11966" *) 4'b1101;
  assign alu_loop_op_4_FpAdd_8U_23U_a_left_shift_acc_3_nl = { 1'b1, _1178_ } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11977" *) 4'b1101;
  assign alu_loop_op_3_FpAdd_8U_23U_a_left_shift_acc_1_nl = { 1'b1, _1179_ } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11988" *) 4'b1101;
  assign alu_loop_op_2_FpAdd_8U_23U_a_left_shift_acc_2_nl = { 1'b1, _1180_ } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11999" *) 4'b1101;
  assign alu_loop_op_1_FpAdd_8U_23U_a_left_shift_acc_nl = { 1'b1, _1181_ } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12010" *) 4'b1101;
  assign alu_loop_op_4_FpMantRNE_49U_24U_else_acc_3_nl = FpAdd_8U_23U_int_mant_1_lpi_1_dfm_2_mx0[47:25] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12318" *) FpMantRNE_49U_24U_else_carry_sva;
  assign alu_loop_op_3_FpMantRNE_49U_24U_else_acc_1_nl = FpAdd_8U_23U_int_mant_4_lpi_1_dfm_2_mx0[47:25] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12358" *) FpMantRNE_49U_24U_else_carry_3_sva;
  assign alu_loop_op_2_FpMantRNE_49U_24U_else_acc_2_nl = FpAdd_8U_23U_int_mant_3_lpi_1_dfm_2_mx0[47:25] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12374" *) FpMantRNE_49U_24U_else_carry_2_sva;
  assign alu_loop_op_1_FpMantRNE_49U_24U_else_acc_nl = FpAdd_8U_23U_int_mant_2_lpi_1_dfm_2_mx0[47:25] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12390" *) FpMantRNE_49U_24U_else_carry_1_sva;
  assign alu_loop_op_3_FpAdd_8U_23U_if_4_if_acc_3_nl = FpAdd_8U_23U_o_expo_3_lpi_1_dfm_13 + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12620" *) 1'b1;
  assign acc_nl = { FpAdd_8U_23U_qr_2_lpi_1_dfm_7, _0045_[8] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12709" *) { _0045_[8], _0045_[8], FpNormalize_8U_49U_else_mux_4_nl, 1'b1 };
  assign acc_1_nl = { FpAdd_8U_23U_qr_3_lpi_1_dfm_7, _0046_[8] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12721" *) { _0046_[8], _0046_[8], FpNormalize_8U_49U_else_mux_5_nl, 1'b1 };
  assign acc_2_nl = { FpAdd_8U_23U_qr_4_lpi_1_dfm_7, _0047_[8] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12733" *) { _0047_[8], _0047_[8], FpNormalize_8U_49U_else_mux_6_nl, 1'b1 };
  assign acc_3_nl = { FpAdd_8U_23U_qr_lpi_1_dfm_7, _0048_[8] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12745" *) { _0048_[8], _0048_[8], FpNormalize_8U_49U_else_mux_7_nl, 1'b1 };
  assign alu_loop_op_2_IntSaturation_33U_32U_if_acc_1_nl = { _0041_[2], _0041_[2], _0041_[0] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12780" *) 1'b1;
  assign alu_loop_op_4_IntSaturation_33U_32U_if_acc_1_nl = { _0042_[2], _0042_[2], _0042_[0] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12794" *) 1'b1;
  assign alu_loop_op_3_IntSaturation_33U_32U_if_acc_nl = { _0043_[2], _0043_[2], _0043_[0] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12798" *) 1'b1;
  assign alu_loop_op_1_IntSaturation_33U_32U_if_acc_nl = { _0044_[2], _0044_[2], _0044_[0] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12802" *) 1'b1;
  assign alu_loop_op_1_FpAdd_8U_23U_if_3_if_acc_1_nl = { 1'b1, FpAdd_8U_23U_qr_2_lpi_1_dfm_7[7:1] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12864" *) 1'b1;
  assign alu_loop_op_2_FpAdd_8U_23U_if_3_if_acc_4_nl = { 1'b1, FpAdd_8U_23U_qr_3_lpi_1_dfm_7[7:1] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12868" *) 1'b1;
  assign alu_loop_op_3_FpAdd_8U_23U_if_3_if_acc_2_nl = { 1'b1, FpAdd_8U_23U_qr_4_lpi_1_dfm_7[7:1] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12872" *) 1'b1;
  assign alu_loop_op_4_FpAdd_8U_23U_if_3_if_acc_6_nl = { 1'b1, FpAdd_8U_23U_qr_lpi_1_dfm_7[7:1] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12876" *) 1'b1;
  assign alu_loop_op_4_FpAdd_8U_23U_if_4_if_acc_7_nl = FpAdd_8U_23U_o_expo_lpi_1_dfm_13 + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12971" *) 1'b1;
  assign acc_8_nl = { alu_loop_op_else_if_mux_8_nl[31], alu_loop_op_else_if_mux_8_nl, 1'b1 } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13015" *) { alu_loop_op_else_if_mux_9_nl[31], alu_loop_op_else_if_mux_9_nl, 1'b1 };
  assign alu_loop_op_else_else_else_else_ac_int_cctor_1_sva = { AluIn_data_sva_127[31], AluIn_data_sva_127[31:0] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13020" *) { else_AluOp_data_0_lpi_1_dfm_mx0[31], else_AluOp_data_0_lpi_1_dfm_mx0 };
  assign acc_10_nl = { alu_loop_op_else_if_mux_12_nl[31], alu_loop_op_else_if_mux_12_nl, 1'b1 } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13027" *) { alu_loop_op_else_if_mux_13_nl[31], alu_loop_op_else_if_mux_13_nl, 1'b1 };
  assign alu_loop_op_else_else_else_else_ac_int_cctor_2_sva = { AluIn_data_sva_127[63], AluIn_data_sva_127[63:32] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13032" *) { else_AluOp_data_1_lpi_1_dfm_mx0[31], else_AluOp_data_1_lpi_1_dfm_mx0 };
  assign acc_11_nl = { alu_loop_op_else_if_mux_14_nl[31], alu_loop_op_else_if_mux_14_nl, 1'b1 } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13039" *) { alu_loop_op_else_if_mux_15_nl[31], alu_loop_op_else_if_mux_15_nl, 1'b1 };
  assign alu_loop_op_else_else_else_else_ac_int_cctor_3_sva = { AluIn_data_sva_127[95], AluIn_data_sva_127[95:64] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13044" *) { else_AluOp_data_2_lpi_1_dfm_mx0[31], else_AluOp_data_2_lpi_1_dfm_mx0 };
  assign acc_9_nl = { alu_loop_op_else_if_mux_10_nl[31], alu_loop_op_else_if_mux_10_nl, 1'b1 } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13051" *) { alu_loop_op_else_if_mux_11_nl[31], alu_loop_op_else_if_mux_11_nl, 1'b1 };
  assign alu_loop_op_else_else_else_else_ac_int_cctor_sva = { AluIn_data_sva_127[127], AluIn_data_sva_127[127:96] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13056" *) { else_AluOp_data_3_lpi_1_dfm_mx0[31], else_AluOp_data_3_lpi_1_dfm_mx0 };
  assign alu_loop_op_1_FpAdd_8U_23U_if_4_if_acc_1_nl = { 1'b1, FpAdd_8U_23U_o_expo_1_lpi_1_dfm_2_mx0w0[7:1] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13059" *) 1'b1;
  assign alu_loop_op_2_FpAdd_8U_23U_if_4_if_acc_4_nl = { 1'b1, FpAdd_8U_23U_o_expo_2_lpi_1_dfm_2_mx0w0[7:1] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13063" *) 1'b1;
  assign alu_loop_op_3_FpAdd_8U_23U_if_4_if_acc_2_nl = { 1'b1, FpAdd_8U_23U_o_expo_3_lpi_1_dfm_2_mx0w0[7:1] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13067" *) 1'b1;
  assign alu_loop_op_4_FpAdd_8U_23U_if_4_if_acc_6_nl = { 1'b1, FpAdd_8U_23U_o_expo_lpi_1_dfm_2_mx0w0[7:1] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13071" *) 1'b1;
  assign alu_loop_op_1_IntSaturation_33U_32U_else_if_acc_nl = { reg_alu_loop_op_else_o_32_1_1_lpi_1_dfm_3_itm, reg_alu_loop_op_else_o_32_1_1_lpi_1_dfm_3_itm, reg_alu_loop_op_else_o_32_1_1_lpi_1_dfm_3_1_itm[30] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13103" *) 1'b1;
  assign alu_loop_op_2_IntSaturation_33U_32U_else_if_acc_1_nl = { reg_alu_loop_op_else_o_32_1_2_lpi_1_dfm_4_itm, reg_alu_loop_op_else_o_32_1_2_lpi_1_dfm_4_itm, reg_alu_loop_op_else_o_32_1_2_lpi_1_dfm_4_1_itm[30] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13107" *) 1'b1;
  assign alu_loop_op_3_IntSaturation_33U_32U_else_if_acc_nl = { reg_alu_loop_op_else_o_32_1_3_lpi_1_dfm_3_itm, reg_alu_loop_op_else_o_32_1_3_lpi_1_dfm_3_itm, reg_alu_loop_op_else_o_32_1_3_lpi_1_dfm_3_1_itm[30] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13111" *) 1'b1;
  assign alu_loop_op_4_IntSaturation_33U_32U_else_if_acc_1_nl = { reg_alu_loop_op_else_o_32_1_lpi_1_dfm_4_itm, reg_alu_loop_op_else_o_32_1_lpi_1_dfm_4_itm, reg_alu_loop_op_else_o_32_1_lpi_1_dfm_4_1_itm[30] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13115" *) 1'b1;
  assign _0460_ = { 1'b1, AluIn_data_sva_127[30:23] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13119" *) _0039_;
  assign FpCmp_8U_23U_false_else_if_acc_4_nl = _0460_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13119" *) 1'b1;
  assign _0461_ = { 1'b1, else_AluOp_data_0_lpi_1_dfm_mx3_30_0[22:0] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13122" *) _0049_;
  assign FpCmp_8U_23U_true_else_else_if_acc_8_nl = _0461_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13122" *) 1'b1;
  assign _0462_ = { 1'b1, else_AluOp_data_2_lpi_1_dfm_mx3_30_0[22:0] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13141" *) _0050_;
  assign FpCmp_8U_23U_true_else_else_if_acc_7_nl = _0462_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13141" *) 1'b1;
  assign _0463_ = { 1'b1, AluIn_data_sva_127[94:87] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13144" *) _0035_;
  assign FpCmp_8U_23U_false_else_if_acc_8_nl = _0463_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13144" *) 1'b1;
  assign _0464_ = { 1'b1, else_AluOp_data_3_lpi_1_dfm_mx0[22:0] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13155" *) _0051_;
  assign FpCmp_8U_23U_true_else_else_if_acc_6_nl = _0464_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13155" *) 1'b1;
  assign _0465_ = { 1'b1, AluIn_data_sva_127[126:119] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13158" *) _0033_;
  assign FpCmp_8U_23U_false_else_if_acc_10_nl = _0465_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13158" *) 1'b1;
  assign _0466_ = { 1'b1, _1136_ } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13208" *) libraries_leading_sign_49_0_78e877fc94067377fcee479dbb0ed8e083a3_4;
  assign alu_loop_op_1_FpNormalize_8U_49U_acc_nl = _0466_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13208" *) 1'b1;
  assign _0467_ = { 1'b1, _1312_ } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13213" *) libraries_leading_sign_49_0_78e877fc94067377fcee479dbb0ed8e083a3_5;
  assign alu_loop_op_2_FpNormalize_8U_49U_acc_2_nl = _0467_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13213" *) 1'b1;
  assign _0468_ = { 1'b1, _1313_ } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13218" *) libraries_leading_sign_49_0_78e877fc94067377fcee479dbb0ed8e083a3_6;
  assign alu_loop_op_3_FpNormalize_8U_49U_acc_1_nl = _0468_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13218" *) 1'b1;
  assign _0469_ = { 1'b1, _1137_ } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13223" *) libraries_leading_sign_49_0_78e877fc94067377fcee479dbb0ed8e083a3_7;
  assign alu_loop_op_4_FpNormalize_8U_49U_acc_3_nl = _0469_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13223" *) 1'b1;
  assign _0470_ = { 1'b1, else_AluOp_data_0_lpi_1_dfm_mx1_tmp_30_23 } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13228" *) _0040_;
  assign FpCmp_8U_23U_true_if_acc_4_nl = _0470_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13228" *) 1'b1;
  assign _0471_ = { 1'b1, else_AluOp_data_1_lpi_1_dfm_mx1_tmp_30_23 } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13233" *) _0038_;
  assign FpCmp_8U_23U_true_if_acc_6_nl = _0471_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13233" *) 1'b1;
  assign _0472_ = { 1'b1, AluIn_data_sva_127[62:55] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13237" *) _0037_;
  assign FpCmp_8U_23U_false_else_if_acc_6_nl = _0472_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13237" *) 1'b1;
  assign _0473_ = { 1'b1, else_else_mux_13_nl } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13244" *) _0052_;
  assign FpCmp_8U_23U_true_else_else_if_acc_4_nl = _0473_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13244" *) 1'b1;
  assign _0474_ = { 1'b1, else_AluOp_data_2_lpi_1_dfm_mx1_tmp_30_23 } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13248" *) _0036_;
  assign FpCmp_8U_23U_true_if_acc_8_nl = _0474_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13248" *) 1'b1;
  assign _0475_ = { 1'b1, else_AluOp_data_3_lpi_1_dfm_mx1_tmp_30_23 } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13253" *) _0034_;
  assign FpCmp_8U_23U_true_if_acc_10_nl = _0475_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13253" *) 1'b1;
  assign _0476_ = { 1'b1, AluIn_data_sva_127[22:0] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13561" *) _0053_;
  assign FpAdd_8U_23U_is_a_greater_oif_aelse_acc_nl = _0476_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13561" *) 1'b1;
  assign _0477_ = { 1'b1, AluIn_data_sva_127[54:32] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13565" *) _0054_;
  assign FpAdd_8U_23U_is_a_greater_oif_aelse_acc_1_nl = _0477_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13565" *) 1'b1;
  assign _0478_ = { 1'b1, AluIn_data_sva_127[86:64] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13569" *) _0055_;
  assign FpAdd_8U_23U_is_a_greater_oif_aelse_acc_2_nl = _0478_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13569" *) 1'b1;
  assign _0479_ = { 1'b1, AluIn_data_sva_127[118:96] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13573" *) _0056_;
  assign FpAdd_8U_23U_is_a_greater_oif_aelse_acc_3_nl = _0479_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13573" *) 1'b1;
  assign alu_loop_op_1_FpAdd_8U_23U_if_4_if_acc_nl = FpAdd_8U_23U_o_expo_1_lpi_1_dfm_13 + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15564" *) 1'b1;
  assign alu_loop_op_2_FpAdd_8U_23U_if_4_if_acc_5_nl = FpAdd_8U_23U_o_expo_2_lpi_1_dfm_13 + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15584" *) 1'b1;
  assign acc_4_nl = { FpAdd_8U_23U_b_right_shift_qif_mux_15_nl, 1'b1 } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16185" *) { FpAdd_8U_23U_b_right_shift_qif_mux_16_nl, 1'b1 };
  assign acc_5_nl = { FpAdd_8U_23U_b_right_shift_qif_mux_17_nl, 1'b1 } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16193" *) { FpAdd_8U_23U_b_right_shift_qif_mux_18_nl, 1'b1 };
  assign acc_6_nl = { FpAdd_8U_23U_b_right_shift_qif_mux_19_nl, 1'b1 } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16201" *) { FpAdd_8U_23U_b_right_shift_qif_mux_20_nl, 1'b1 };
  assign acc_7_nl = { FpAdd_8U_23U_b_right_shift_qif_mux_21_nl, 1'b1 } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16209" *) { FpAdd_8U_23U_b_right_shift_qif_mux_22_nl, 1'b1 };
  assign acc_12_nl = { _1474_, FpAdd_8U_23U_else_2_mux_8_nl, _1474_ } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16218" *) { FpAdd_8U_23U_else_2_mux_9_nl, 1'b1 };
  assign acc_13_nl = { _1475_, FpAdd_8U_23U_else_2_mux_10_nl, _1475_ } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16227" *) { FpAdd_8U_23U_else_2_mux_11_nl, 1'b1 };
  assign acc_14_nl = { _1476_, FpAdd_8U_23U_else_2_mux_12_nl, _1476_ } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16236" *) { FpAdd_8U_23U_else_2_mux_13_nl, 1'b1 };
  assign acc_15_nl = { _1477_, FpAdd_8U_23U_else_2_mux_14_nl, _1477_ } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16245" *) { FpAdd_8U_23U_else_2_mux_15_nl, 1'b1 };
  assign _0480_ = and_dcpl_37 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12265" *) or_1087_cse;
  assign chn_alu_out_and_cse = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12266" *) chn_alu_out_or_cse;
  assign chn_alu_out_and_1_cse = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12267" *) _1182_;
  assign _0481_ = _1482_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12272" *) or_1087_cse;
  assign _0482_ = _0481_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12272" *) main_stage_v_4;
  assign and_734_cse = _0482_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12272" *) core_wen;
  assign chn_alu_out_and_8_cse = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12273" *) _1184_;
  assign chn_alu_out_and_18_cse = chn_alu_out_and_8_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12274" *) _1182_;
  assign _0483_ = or_16_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12275" *) _1186_;
  assign and_502_nl = or_1087_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12276" *) chn_alu_in_rsci_bawt;
  assign _0484_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12278" *) _1187_;
  assign AluIn_data_and_cse = _0484_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12278" *) mux_15_nl;
  assign _0485_ = or_dcpl_14 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12282" *) and_dcpl_78;
  assign _0486_ = or_963_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12287" *) cfg_alu_bypass_rsc_triosy_obj_bawt;
  assign _0487_ = _0486_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12288" *) cfg_alu_src_rsc_triosy_obj_bawt;
  assign _0488_ = _0487_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12288" *) cfg_alu_op_rsc_triosy_obj_bawt;
  assign and_501_cse = _0488_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12288" *) cfg_alu_algo_rsc_triosy_obj_bawt;
  assign _0489_ = or_tmp_386 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12289" *) _1190_;
  assign _0490_ = _0489_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12290" *) main_stage_v_1;
  assign and_167_rgt = _0490_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12290" *) alu_loop_op_2_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_1_svs_2;
  assign _0491_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12291" *) _1191_;
  assign IsNaN_8U_23U_aelse_and_cse = _0491_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12291" *) not_tmp_29;
  assign _0492_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12295" *) FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_or_7_cse;
  assign FpAdd_8U_23U_is_addition_and_8_cse = _0492_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12295" *) not_tmp_29;
  assign and_dcpl_3 = cfg_alu_bypass_rsc_triosy_obj_bawt & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12297" *) cfg_alu_src_rsc_triosy_obj_bawt;
  assign and_dcpl_28 = and_dcpl_3 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12298" *) cfg_alu_op_rsc_triosy_obj_bawt;
  assign and_486_cse = and_dcpl_28 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12298" *) cfg_alu_algo_rsc_triosy_obj_bawt;
  assign _0493_ = and_486_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12298" *) or_963_cse;
  assign else_AluOp_data_and_10_cse = _0491_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12301" *) mux_43_nl;
  assign AluIn_data_and_1_cse = _0491_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12305" *) mux_46_nl;
  assign FpAdd_8U_23U_and_39_cse = _0491_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12306" *) not_tmp_57;
  assign FpAdd_8U_23U_int_mant_p1_and_4_cse = _0492_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12309" *) not_tmp_57;
  assign and_550_cse = _0491_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12310" *) mux_tmp_53;
  assign _0494_ = or_1087_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12312" *) _1196_;
  assign and_192_nl = or_1087_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12324" *) _1200_;
  assign _0495_ = _1201_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12333" *) FpAlu_8U_23U_equal_tmp_22;
  assign IsNaN_8U_23U_aelse_and_8_cse = _0491_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12348" *) mux_107_nl;
  assign IsNaN_8U_23U_1_aelse_and_cse = _0491_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12349" *) _1207_;
  assign FpMantRNE_49U_24U_else_and_4_cse = _0492_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12356" *) _1208_;
  assign and_196_nl = or_1087_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12364" *) _1209_;
  assign and_200_nl = or_1087_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12380" *) _1210_;
  assign and_204_nl = or_1087_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12396" *) _1211_;
  assign FpAlu_8U_23U_and_82_cse = _0491_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12408" *) _1212_;
  assign FpCmp_8U_23U_true_o_and_cse = _0491_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12416" *) _1214_;
  assign and_211_rgt = or_1087_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12417" *) _1215_;
  assign FpCmp_8U_23U_false_o_and_1_cse = _0491_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12421" *) _1217_;
  assign and_213_rgt = or_1087_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12422" *) _1218_;
  assign and_215_rgt = or_1087_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12423" *) _1219_;
  assign _0496_ = _1480_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12427" *) or_1087_cse;
  assign _0497_ = _0496_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12427" *) nor_397_cse;
  assign _0498_ = _0497_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12427" *) main_stage_v_4;
  assign and_524_cse = _0498_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12428" *) core_wen;
  assign and_217_rgt = or_1087_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12429" *) _1220_;
  assign and_cse = _0491_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12431" *) mux_140_nl;
  assign AluOut_data_and_8_cse = _0491_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12432" *) _1221_;
  assign IntSaturation_33U_32U_and_cse = _0491_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12434" *) _1222_;
  assign FpMantRNE_49U_24U_else_and_cse = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12435" *) _1223_;
  assign FpAdd_8U_23U_int_mant_p1_and_cse = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12439" *) _1224_;
  assign FpAdd_8U_23U_int_mant_p1_and_12_cse = FpAdd_8U_23U_int_mant_p1_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12441" *) _1225_;
  assign FpAdd_8U_23U_if_3_and_cse = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12442" *) _1226_;
  assign _0499_ = main_stage_v_1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12447" *) _1227_;
  assign _0500_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12450" *) cfg_alu_algo_cfg_alu_algo_or_3_cse;
  assign IsZero_8U_23U_and_4_cse = _0500_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12450" *) _1228_;
  assign IsZero_8U_23U_1_and_cse = chn_alu_out_and_8_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12451" *) _1229_;
  assign FpAdd_8U_23U_is_addition_and_cse = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12452" *) _1229_;
  assign _0501_ = or_16_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12455" *) cfg_alu_bypass_rsc_triosy_obj_bawt;
  assign _0502_ = _0501_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12456" *) cfg_alu_src_rsc_triosy_obj_bawt;
  assign _0503_ = _0502_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12456" *) cfg_alu_op_rsc_triosy_obj_bawt;
  assign _0504_ = _0503_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12456" *) cfg_alu_algo_rsc_triosy_obj_bawt;
  assign and_489_cse = _1230_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12456" *) main_stage_v_1;
  assign and_231_rgt = and_dcpl_78 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12457" *) FpAdd_8U_23U_is_a_greater_lor_1_lpi_1_dfm_1_mx0w0;
  assign _0505_ = and_dcpl_78 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12458" *) or_dcpl_117;
  assign and_233_rgt = _0505_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12458" *) _1231_;
  assign and_235_rgt = and_dcpl_78 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12459" *) FpAdd_8U_23U_is_a_greater_lor_2_lpi_1_dfm_1_mx0w0;
  assign _0506_ = and_dcpl_78 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12460" *) or_dcpl_119;
  assign and_237_rgt = _0506_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12460" *) _1232_;
  assign and_239_rgt = and_dcpl_78 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12461" *) FpAdd_8U_23U_is_a_greater_lor_3_lpi_1_dfm_1_mx0w0;
  assign _0507_ = and_dcpl_78 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12462" *) or_dcpl_121;
  assign and_241_rgt = _0507_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12462" *) _1233_;
  assign and_243_rgt = and_dcpl_78 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12463" *) FpAdd_8U_23U_is_a_greater_lor_lpi_1_dfm_1_mx0w0;
  assign _0508_ = and_dcpl_78 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12464" *) or_dcpl_123;
  assign and_245_rgt = _0508_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12464" *) _1234_;
  assign _0509_ = cfg_alu_algo_1_sva_st_24[1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12471" *) FpAlu_8U_23U_nor_dfs_5;
  assign _0510_ = FpAlu_8U_23U_equal_tmp_22 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12471" *) _1533_;
  assign IsNaN_8U_23U_aelse_and_12_cse = _0491_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12473" *) mux_177_nl;
  assign _0511_ = or_1087_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12474" *) _1237_;
  assign _0512_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12481" *) FpAlu_8U_23U_o_FpAlu_8U_23U_o_or_cse;
  assign AluOut_data_and_12_cse = _0512_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12481" *) _1238_;
  assign FpAlu_8U_23U_and_88_cse = _0491_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12482" *) _1239_;
  assign FpCmp_8U_23U_true_o_and_5_cse = _0491_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12489" *) _1241_;
  assign FpCmp_8U_23U_false_o_and_6_cse = _0491_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12496" *) _1244_;
  assign IntSaturation_33U_32U_and_11_cse = _0491_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12504" *) _1245_;
  assign alu_loop_bypass_if_and_6_cse = _1237_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12505" *) and_dcpl_171;
  assign alu_loop_bypass_if_and_7_cse = alu_loop_op_unequal_tmp_6 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12506" *) and_dcpl_171;
  assign _0513_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12508" *) _1547_;
  assign AluOut_data_and_15_cse = _0513_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12508" *) mux_tmp_53;
  assign _0514_ = or_963_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12509" *) and_dcpl_77;
  assign _0515_ = _0514_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12509" *) main_stage_v_1;
  assign _0516_ = _0515_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12510" *) cfg_alu_bypass_rsc_triosy_obj_bawt;
  assign _0517_ = _0516_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12510" *) cfg_alu_src_rsc_triosy_obj_bawt;
  assign _0518_ = _0517_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12510" *) cfg_alu_op_rsc_triosy_obj_bawt;
  assign _0519_ = _0518_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12511" *) cfg_alu_algo_rsc_triosy_obj_bawt;
  assign and_485_nl = _0519_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12511" *) _0009_;
  assign FpAlu_8U_23U_and_94_cse = _0491_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12514" *) mux_214_nl;
  assign _0520_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12517" *) _1246_;
  assign IsZero_8U_23U_and_6_cse = _0520_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12517" *) _1247_;
  assign _0521_ = cfg_alu_algo_1_sva_st_23[1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12524" *) FpAlu_8U_23U_nor_dfs_4;
  assign _0522_ = FpAlu_8U_23U_equal_tmp_21 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12524" *) _1557_;
  assign IsNaN_8U_23U_aelse_and_16_cse = _0491_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12526" *) mux_217_nl;
  assign _0523_ = _0515_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12528" *) _1190_;
  assign _0524_ = _0523_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12528" *) cfg_alu_bypass_rsc_triosy_obj_bawt;
  assign _0525_ = _0524_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12529" *) cfg_alu_src_rsc_triosy_obj_bawt;
  assign _0526_ = _0525_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12529" *) cfg_alu_op_rsc_triosy_obj_bawt;
  assign _0527_ = _0526_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12530" *) cfg_alu_algo_rsc_triosy_obj_bawt;
  assign _0528_ = _0527_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12530" *) FpAlu_8U_23U_equal_tmp_1_mx0w0;
  assign and_481_cse = _0528_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12530" *) _0009_;
  assign AluOut_data_and_5_cse = alu_loop_op_else_nor_dfs & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12531" *) and_dcpl_208;
  assign _0529_ = main_stage_v_1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12536" *) cfg_alu_bypass_rsc_triosy_obj_bawt;
  assign _0530_ = _0529_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12537" *) cfg_alu_src_rsc_triosy_obj_bawt;
  assign _0531_ = _0530_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12537" *) cfg_alu_op_rsc_triosy_obj_bawt;
  assign _0532_ = _0531_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12537" *) cfg_alu_algo_rsc_triosy_obj_bawt;
  assign and_484_cse = _0532_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12538" *) _0009_;
  assign and_478_nl = and_484_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12538" *) mux_221_nl;
  assign AluOut_data_and_17_cse = _0491_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12541" *) mux_222_nl;
  assign FpCmp_8U_23U_true_o_and_9_cse = _0491_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12550" *) mux_224_nl;
  assign and_293_rgt = or_1087_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12559" *) io_read_cfg_alu_bypass_rsc_svs_st_1;
  assign IntSaturation_33U_32U_if_and_9_cse = _0491_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12564" *) not_tmp_232;
  assign FpAlu_8U_23U_and_102_cse = _0491_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12570" *) _1256_;
  assign _0533_ = alu_loop_op_else_nor_dfs & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12571" *) and_dcpl_214;
  assign _0534_ = FpAlu_8U_23U_equal_tmp_2_mx0w0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12572" *) and_dcpl_214;
  assign and_297_m1c = _1257_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12573" *) or_1087_cse;
  assign IsNaN_8U_23U_2_and_cse = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12588" *) IsNaN_8U_23U_2_IsNaN_8U_23U_2_or_5_cse;
  assign IsNaN_8U_23U_2_and_6_cse = IsNaN_8U_23U_2_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12588" *) _1258_;
  assign _0535_ = chn_alu_out_and_8_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12600" *) IsNaN_8U_23U_2_IsNaN_8U_23U_2_or_3_cse;
  assign IsNaN_8U_23U_2_and_9_cse = _0535_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12600" *) _1259_;
  assign _0536_ = or_dcpl_14 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12603" *) and_dcpl_234;
  assign _0537_ = _0536_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12603" *) or_1087_cse;
  assign and_328_rgt = _0537_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12603" *) _0004_;
  assign _0538_ = _1260_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12623" *) FpAdd_8U_23U_FpAdd_8U_23U_nor_9_m1c;
  assign FpAdd_8U_23U_and_31_nl = _0538_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12623" *) FpAlu_8U_23U_nor_dfs_6;
  assign _0539_ = FpAdd_8U_23U_and_2_tmp_3 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12625" *) _1261_;
  assign _0540_ = _0539_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12625" *) FpAdd_8U_23U_FpAdd_8U_23U_nor_9_m1c;
  assign FpAdd_8U_23U_and_19_nl = _0540_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12625" *) FpAlu_8U_23U_nor_dfs_6;
  assign _0541_ = FpAdd_8U_23U_is_inf_3_lpi_1_dfm_8 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12627" *) FpAdd_8U_23U_FpAdd_8U_23U_nor_9_m1c;
  assign FpAdd_8U_23U_and_32_nl = _0541_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12627" *) FpAlu_8U_23U_nor_dfs_6;
  assign _0542_ = IsNaN_8U_23U_1_land_3_lpi_1_dfm_9 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12629" *) _1262_;
  assign FpAdd_8U_23U_and_21_nl = _0542_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12629" *) FpAlu_8U_23U_nor_dfs_6;
  assign _0543_ = _1263_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12659" *) alu_loop_op_4_FpAdd_8U_23U_is_a_greater_oif_equal_3_tmp;
  assign _0544_ = _1264_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12669" *) alu_loop_op_3_FpAdd_8U_23U_is_a_greater_oif_equal_1_tmp;
  assign _0545_ = _1265_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12680" *) alu_loop_op_2_FpAdd_8U_23U_is_a_greater_oif_equal_2_tmp;
  assign _0546_ = _1266_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12691" *) alu_loop_op_1_FpAdd_8U_23U_is_a_greater_oif_equal_tmp;
  assign FpAdd_8U_23U_and_4_tmp = _1267_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12704" *) FpAdd_8U_23U_int_mant_p1_1_lpi_1_dfm_5[49];
  assign FpAdd_8U_23U_and_10_tmp = _1268_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12716" *) FpAdd_8U_23U_int_mant_p1_2_lpi_1_dfm_5[49];
  assign FpAdd_8U_23U_and_16_tmp = _1269_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12728" *) FpAdd_8U_23U_int_mant_p1_3_lpi_1_dfm_5[49];
  assign FpAdd_8U_23U_and_22_tmp = _1270_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12740" *) FpAdd_8U_23U_int_mant_p1_lpi_1_dfm_5[49];
  assign _0547_ = FpCmp_8U_23U_true_else_else_if_acc_4_nl[23] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12823" *) _1277_;
  assign alu_loop_op_4_FpMantRNE_49U_24U_else_and_3_tmp = FpMantRNE_49U_24U_else_carry_sva & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12880" *) _1140_;
  assign FpMantRNE_49U_24U_else_carry_sva = FpAdd_8U_23U_int_mant_1_lpi_1_dfm_2_mx0[24] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12894" *) _1618_;
  assign alu_loop_op_3_FpMantRNE_49U_24U_else_and_1_tmp = FpMantRNE_49U_24U_else_carry_3_sva & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12900" *) _1141_;
  assign FpMantRNE_49U_24U_else_carry_3_sva = FpAdd_8U_23U_int_mant_4_lpi_1_dfm_2_mx0[24] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12914" *) _1642_;
  assign alu_loop_op_2_FpMantRNE_49U_24U_else_and_2_tmp = FpMantRNE_49U_24U_else_carry_2_sva & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12920" *) _1142_;
  assign FpMantRNE_49U_24U_else_carry_2_sva = FpAdd_8U_23U_int_mant_3_lpi_1_dfm_2_mx0[24] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12934" *) _1666_;
  assign alu_loop_op_1_FpMantRNE_49U_24U_else_and_tmp = FpMantRNE_49U_24U_else_carry_1_sva & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12940" *) _1143_;
  assign FpMantRNE_49U_24U_else_carry_1_sva = FpAdd_8U_23U_int_mant_2_lpi_1_dfm_2_mx0[24] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12954" *) _1690_;
  assign _0548_ = _1278_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12974" *) FpAdd_8U_23U_FpAdd_8U_23U_nor_11_m1c;
  assign FpAdd_8U_23U_and_33_nl = _0548_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12974" *) FpAlu_8U_23U_nor_dfs_6;
  assign _0549_ = FpAdd_8U_23U_and_3_tmp_3 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12976" *) _1279_;
  assign _0550_ = _0549_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12976" *) FpAdd_8U_23U_FpAdd_8U_23U_nor_11_m1c;
  assign FpAdd_8U_23U_and_25_nl = _0550_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12976" *) FpAlu_8U_23U_nor_dfs_6;
  assign _0551_ = FpAdd_8U_23U_is_inf_lpi_1_dfm_8 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12978" *) FpAdd_8U_23U_FpAdd_8U_23U_nor_11_m1c;
  assign FpAdd_8U_23U_and_34_nl = _0551_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12978" *) FpAlu_8U_23U_nor_dfs_6;
  assign _0552_ = IsNaN_8U_23U_1_land_lpi_1_dfm_9 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12980" *) _1280_;
  assign FpAdd_8U_23U_and_27_nl = _0552_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12980" *) FpAlu_8U_23U_nor_dfs_6;
  assign FpAlu_8U_23U_and_62_nl = IsNaN_8U_23U_land_lpi_1_dfm_11 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12981" *) FpAlu_8U_23U_nor_dfs_6;
  assign FpAlu_8U_23U_and_30_cse = _1281_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13000" *) FpAlu_8U_23U_equal_tmp_29;
  assign FpAlu_8U_23U_and_31_m1c = FpAlu_8U_23U_equal_tmp_32 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13001" *) FpAlu_8U_23U_equal_tmp_29;
  assign FpAlu_8U_23U_and_44_cse = _1282_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13002" *) FpAlu_8U_23U_equal_tmp_29;
  assign FpAlu_8U_23U_and_45_cse = FpAlu_8U_23U_and_12_tmp & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13003" *) FpAlu_8U_23U_equal_tmp_29;
  assign FpAlu_8U_23U_and_12_tmp = FpAlu_8U_23U_equal_tmp_35 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13004" *) FpAlu_8U_23U_equal_tmp_32;
  assign _0553_ = cfg_alu_src_1_sva_st_1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13006" *) _1190_;
  assign _0554_ = _0553_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13006" *) main_stage_v_1;
  assign _0555_ = chn_alu_in_rsci_bawt & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13006" *) _1695_;
  assign _0556_ = _0555_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13007" *) _1696_;
  assign _0557_ = _0556_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13008" *) _1697_;
  assign _0558_ = _0557_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13008" *) _1698_;
  assign _0559_ = _0558_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13009" *) _1699_;
  assign main_stage_en_1 = _0559_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13009" *) or_1087_cse;
  assign IntSaturation_33U_32U_and_3_nl = alu_loop_op_2_IntSaturation_33U_32U_else_if_acc_1_nl[2] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13077" *) _1284_;
  assign IntSaturation_33U_32U_and_7_nl = alu_loop_op_4_IntSaturation_33U_32U_else_if_acc_1_nl[2] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13084" *) _1285_;
  assign IntSaturation_33U_32U_and_5_nl = alu_loop_op_3_IntSaturation_33U_32U_else_if_acc_nl[2] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13091" *) _1286_;
  assign IntSaturation_33U_32U_and_1_nl = alu_loop_op_1_IntSaturation_33U_32U_else_if_acc_nl[2] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13098" *) _1287_;
  assign and_446_nl = else_mux_tmp_31_23[8] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13127" *) or_tmp_668;
  assign _0560_ = _1152_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13137" *) _1144_;
  assign and_444_nl = else_mux_2_tmp_31_23[8] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13149" *) or_tmp_674;
  assign and_443_nl = else_mux_3_tmp_31_23[8] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13163" *) or_tmp_678;
  assign and_336_nl = AluIn_data_sva_127[31] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13168" *) or_tmp_668;
  assign and_338_nl = AluIn_data_sva_127[95] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13174" *) or_tmp_674;
  assign and_340_nl = AluIn_data_sva_127[127] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13181" *) or_tmp_678;
  assign FpCmp_8U_23U_false_else_1_FpCmp_8U_23U_false_else_1_and_1_nl = _1302_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13189" *) else_AluOp_data_1_lpi_1_dfm_mx0[31];
  assign _0561_ = _1721_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13195" *) _1303_;
  assign FpAlu_8U_23U_and_61_nl = _0561_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13195" *) FpAlu_8U_23U_equal_tmp_2_mx0w0;
  assign FpAlu_8U_23U_and_48_m1c = _1304_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13198" *) FpAlu_8U_23U_and_34_m1c;
  assign FpAlu_8U_23U_and_34_m1c = _1305_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13199" *) FpAlu_8U_23U_nor_dfs_mx0w0;
  assign FpAlu_8U_23U_and_52_m1c = _1306_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13200" *) FpAlu_8U_23U_and_36_m1c;
  assign FpAlu_8U_23U_and_36_m1c = _1307_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13201" *) FpAlu_8U_23U_nor_dfs_mx0w0;
  assign FpAlu_8U_23U_and_56_m1c = _1308_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13202" *) FpAlu_8U_23U_and_38_m1c;
  assign FpAlu_8U_23U_and_38_m1c = _1309_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13203" *) FpAlu_8U_23U_nor_dfs_mx0w0;
  assign FpAlu_8U_23U_and_40_m1c = _1310_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13204" *) FpAlu_8U_23U_and_24_m1c;
  assign FpAlu_8U_23U_and_24_m1c = _1311_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13205" *) FpAlu_8U_23U_nor_dfs_mx0w0;
  assign FpNormalize_8U_49U_oelse_not_9 = FpNormalize_8U_49U_if_or_itm_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13210" *) alu_loop_op_1_FpNormalize_8U_49U_acc_nl[8];
  assign FpNormalize_8U_49U_oelse_not_11 = FpNormalize_8U_49U_if_or_1_itm_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13215" *) alu_loop_op_2_FpNormalize_8U_49U_acc_2_nl[8];
  assign FpNormalize_8U_49U_oelse_not_13 = FpNormalize_8U_49U_if_or_2_itm_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13220" *) alu_loop_op_3_FpNormalize_8U_49U_acc_1_nl[8];
  assign FpNormalize_8U_49U_oelse_not_15 = FpNormalize_8U_49U_if_or_3_itm_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13225" *) alu_loop_op_4_FpNormalize_8U_49U_acc_3_nl[8];
  assign asn_267 = alu_loop_op_unequal_tmp_8 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13226" *) _1314_;
  assign and_dcpl_2 = cfg_alu_op_rsc_triosy_obj_bawt & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13265" *) cfg_alu_algo_rsc_triosy_obj_bawt;
  assign and_dcpl_4 = and_dcpl_3 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13267" *) and_dcpl_2;
  assign and_tmp = and_501_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13269" *) or_1087_cse;
  assign and_37_cse = and_486_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13273" *) or_1087_cse;
  assign _0562_ = io_read_cfg_alu_bypass_rsc_svs_st_1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13286" *) _1317_;
  assign _0563_ = cfg_alu_src_rsci_d & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13290" *) chn_alu_in_rsci_bawt;
  assign _0564_ = cfg_alu_algo_1_sva_st_22[1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13294" *) cfg_alu_bypass_rsc_triosy_obj_bawt;
  assign _0565_ = _0564_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13294" *) cfg_alu_src_rsc_triosy_obj_bawt;
  assign _0566_ = _0565_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13294" *) cfg_alu_op_rsc_triosy_obj_bawt;
  assign _0567_ = _0566_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13295" *) cfg_alu_algo_rsc_triosy_obj_bawt;
  assign _0568_ = _0567_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13295" *) or_963_cse;
  assign _0569_ = main_stage_v_1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13352" *) _1323_;
  assign not_tmp_157 = main_stage_v_1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13356" *) mux_163_nl;
  assign nor_tmp_74 = io_read_cfg_alu_bypass_rsc_svs_5 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13361" *) io_read_cfg_alu_bypass_rsc_svs_st_1;
  assign _0570_ = or_963_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13383" *) or_1050_cse;
  assign _0571_ = _0570_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13383" *) main_stage_v_1;
  assign _0572_ = _0571_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13384" *) cfg_alu_bypass_rsc_triosy_obj_bawt;
  assign _0573_ = _0572_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13384" *) cfg_alu_src_rsc_triosy_obj_bawt;
  assign _0574_ = _0573_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13384" *) cfg_alu_op_rsc_triosy_obj_bawt;
  assign _0575_ = _0574_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13385" *) cfg_alu_algo_rsc_triosy_obj_bawt;
  assign and_474_nl = _0575_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13385" *) _0009_;
  assign _0002_ = main_stage_v_1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13412" *) _1324_;
  assign _0576_ = cfg_alu_algo_1_sva_st[0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13424" *) _1147_;
  assign and_tmp_35 = cfg_alu_algo_1_sva_st[0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13442" *) or_28_cse;
  assign _0577_ = and_dcpl_4 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13447" *) or_16_cse;
  assign _0578_ = _1326_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13447" *) main_stage_v_1;
  assign _0579_ = and_dcpl_28 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13450" *) _1779_;
  assign _0580_ = _0579_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13450" *) cfg_alu_algo_rsc_triosy_obj_bawt;
  assign _0581_ = _1327_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13450" *) main_stage_v_1;
  assign and_dcpl_30 = _1328_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13450" *) or_1087_cse;
  assign and_dcpl_32 = _1329_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13451" *) reg_chn_alu_out_rsci_ld_core_psct_cse;
  assign and_dcpl_33 = _1330_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13452" *) cfg_alu_src_1_sva_st_1;
  assign and_dcpl_34 = and_dcpl_33 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13453" *) _1190_;
  assign and_dcpl_35 = _1780_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13456" *) main_stage_v_1;
  assign and_dcpl_37 = main_stage_v_4 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13457" *) io_read_cfg_alu_bypass_rsc_svs_8;
  assign _0582_ = main_stage_v_4 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13458" *) _1314_;
  assign and_dcpl_40 = _0582_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13458" *) or_1087_cse;
  assign and_dcpl_43 = or_1087_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13460" *) main_stage_v_4;
  assign _0583_ = _1206_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13461" *) chn_alu_out_rsci_bawt;
  assign and_dcpl_45 = _0583_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13461" *) reg_chn_alu_out_rsci_ld_core_psct_cse;
  assign and_dcpl_46 = chn_alu_in_rsci_bawt & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13462" *) _1331_;
  assign and_dcpl_349 = cfg_alu_src_rsc_triosy_obj_bawt & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13464" *) cfg_alu_op_rsc_triosy_obj_bawt;
  assign and_dcpl_53 = and_dcpl_349 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13464" *) cfg_alu_algo_rsc_triosy_obj_bawt;
  assign _0584_ = or_16_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13465" *) or_1087_cse;
  assign _0585_ = _0584_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13465" *) and_dcpl_28;
  assign _0586_ = _0585_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13466" *) cfg_alu_algo_rsc_triosy_obj_bawt;
  assign and_dcpl_64 = _0586_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13466" *) main_stage_v_1;
  assign and_dcpl_70 = and_dcpl_28 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13467" *) or_1087_cse;
  assign and_dcpl_78 = and_dcpl_77 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13471" *) or_1087_cse;
  assign and_dcpl_80 = or_dcpl_14 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13472" *) or_1050_cse;
  assign and_dcpl_81 = and_dcpl_80 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13473" *) or_1087_cse;
  assign _0587_ = or_dcpl_14 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13474" *) and_dcpl_46;
  assign and_dcpl_83 = _0587_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13474" *) or_1087_cse;
  assign and_dcpl_89 = chn_alu_in_rsci_bawt & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13475" *) cfg_alu_bypass_rsci_d;
  assign and_dcpl_96 = or_1087_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13476" *) main_stage_v_2;
  assign and_dcpl_99 = or_1050_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13477" *) or_1087_cse;
  assign and_dcpl_108 = or_1087_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13478" *) alu_loop_op_unequal_tmp_7;
  assign nor_tmp_144 = alu_loop_op_unequal_tmp_7 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13482" *) main_stage_v_3;
  assign and_dcpl_127 = nor_tmp_144 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13483" *) or_1087_cse;
  assign and_dcpl_165 = or_1087_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13503" *) alu_loop_op_unequal_tmp_6;
  assign and_dcpl_167 = or_1087_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13504" *) cfg_precision[1];
  assign _0588_ = and_dcpl_167 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13505" *) _1337_;
  assign and_dcpl_168 = _0588_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13505" *) _1237_;
  assign and_dcpl_169 = and_dcpl_99 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13506" *) _1237_;
  assign and_dcpl_170 = or_1087_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13507" *) io_read_cfg_alu_bypass_rsc_svs_6;
  assign and_dcpl_171 = or_1087_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13508" *) _1338_;
  assign _0589_ = and_dcpl_70 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13513" *) cfg_alu_algo_rsc_triosy_obj_bawt;
  assign _0590_ = _0589_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13514" *) cfg_precision[1];
  assign and_dcpl_179 = _0590_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13514" *) or_963_cse;
  assign and_dcpl_207 = _0588_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13515" *) _1190_;
  assign and_dcpl_208 = _1797_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13516" *) or_1087_cse;
  assign and_dcpl_214 = mux_tmp_323 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13519" *) or_1087_cse;
  assign and_dcpl_217 = and_dcpl_77 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13520" *) _0004_;
  assign _0591_ = or_dcpl_14 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13521" *) and_dcpl_217;
  assign and_dcpl_229 = _0591_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13521" *) or_1087_cse;
  assign and_dcpl_219 = and_dcpl_229 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13521" *) _1340_;
  assign _0592_ = or_dcpl_14 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13522" *) and_dcpl_77;
  assign _0593_ = _0592_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13522" *) cfg_alu_algo_rsci_d[0];
  assign and_dcpl_222 = _0593_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13522" *) or_1087_cse;
  assign and_dcpl_225 = and_dcpl_229 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13523" *) cfg_alu_algo_rsci_d[1];
  assign and_dcpl_227 = and_dcpl_81 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13525" *) _1341_;
  assign and_dcpl_231 = and_dcpl_81 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13527" *) cfg_alu_algo_1_sva_st[1];
  assign and_dcpl_234 = and_dcpl_46 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13528" *) and_dcpl_77;
  assign _0594_ = _0536_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13530" *) _1145_;
  assign and_dcpl_236 = _0594_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13530" *) or_1087_cse;
  assign and_dcpl_239 = _0537_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13531" *) cfg_alu_algo_rsci_d[0];
  assign _0595_ = _0536_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13533" *) _1146_;
  assign and_dcpl_243 = _0595_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13533" *) or_1087_cse;
  assign _0596_ = or_dcpl_14 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13537" *) or_1087_cse;
  assign _0597_ = _0596_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13537" *) chn_alu_in_rsci_bawt;
  assign or_tmp_695 = _0597_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13537" *) fsm_output[1];
  assign _0598_ = _0596_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13538" *) and_dcpl_46;
  assign _0599_ = _0598_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13539" *) cfg_alu_src_rsci_d;
  assign and_357_cse = _0599_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13539" *) fsm_output[1];
  assign _0600_ = or_1087_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13542" *) cfg_alu_bypass_rsc_triosy_obj_bawt;
  assign _0601_ = _0600_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13542" *) chn_alu_op_rsci_bawt;
  assign _0602_ = _0601_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13542" *) cfg_alu_src_1_sva_st_1;
  assign _0603_ = _0602_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13543" *) _1190_;
  assign _0604_ = _0603_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13543" *) main_stage_v_1;
  assign _0605_ = _0604_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13543" *) and_dcpl_53;
  assign chn_alu_op_rsci_ld_core_psct_mx0c1 = _0605_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13543" *) _1798_;
  assign _0606_ = _0600_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13545" *) or_16_cse;
  assign _0607_ = _0606_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13545" *) and_dcpl_53;
  assign _0608_ = _0607_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13545" *) _1188_;
  assign main_stage_v_1_mx0c1 = _0608_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13545" *) main_stage_v_1;
  assign _0609_ = or_dcpl_14 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13546" *) and_dcpl_89;
  assign _0610_ = _0609_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13546" *) or_1087_cse;
  assign _0611_ = _0610_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13547" *) fsm_output[1];
  assign _0612_ = and_dcpl_30 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13547" *) and_dcpl_89;
  assign _0613_ = _0612_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13547" *) cfg_alu_src_1_sva_st_1;
  assign main_stage_v_2_mx0c1 = _1799_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13549" *) and_dcpl_96;
  assign _0614_ = main_stage_v_3 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13550" *) _1194_;
  assign main_stage_v_3_mx0c1 = _0614_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13550" *) or_1087_cse;
  assign _0615_ = _1203_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13551" *) main_stage_v_4;
  assign main_stage_v_4_mx0c1 = _0615_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13551" *) or_1087_cse;
  assign _0616_ = and_dcpl_179 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13552" *) and_dcpl_175;
  assign _0617_ = _0616_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13553" *) main_stage_v_1;
  assign _0618_ = _0617_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13553" *) _1231_;
  assign FpAdd_8U_23U_qr_2_lpi_1_dfm_mx0c1 = _0618_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13553" *) or_dcpl_117;
  assign _0619_ = _0617_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13555" *) _1232_;
  assign FpAdd_8U_23U_qr_3_lpi_1_dfm_mx0c1 = _0619_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13555" *) or_dcpl_119;
  assign _0620_ = _0617_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13557" *) _1233_;
  assign FpAdd_8U_23U_qr_4_lpi_1_dfm_mx0c1 = _0620_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13557" *) or_dcpl_121;
  assign _0621_ = _0617_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13559" *) _1234_;
  assign FpAdd_8U_23U_qr_lpi_1_dfm_mx0c1 = _0621_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13559" *) or_dcpl_123;
  assign _0622_ = _0589_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13578" *) chn_alu_op_rsci_bawt;
  assign _0623_ = _0622_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13578" *) cfg_alu_src_1_sva_st_1;
  assign _0624_ = _0623_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13579" *) _1190_;
  assign chn_alu_op_rsci_oswt_unreg = _0624_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13579" *) main_stage_v_1;
  assign chn_alu_out_rsci_oswt_unreg = chn_alu_out_rsci_bawt & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13580" *) reg_chn_alu_out_rsci_ld_core_psct_cse;
  assign and_dcpl_269 = nor_397_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13582" *) _1204_;
  assign _0625_ = and_dcpl_269 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13583" *) FpAlu_8U_23U_nor_dfs_6;
  assign _0626_ = _0625_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13583" *) IsNaN_8U_23U_land_1_lpi_1_dfm_11;
  assign _0627_ = _0625_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13585" *) IsNaN_8U_23U_land_2_lpi_1_dfm_11;
  assign _0628_ = and_dcpl_269 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13587" *) IsNaN_8U_23U_land_3_lpi_1_dfm_11;
  assign _0629_ = _0628_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13587" *) FpAlu_8U_23U_nor_dfs_6;
  assign and_dcpl = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13589" *) main_stage_v_3;
  assign FpAdd_8U_23U_if_3_if_and_tmp = fsm_output[1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13591" *) FpAdd_8U_23U_int_mant_p1_1_lpi_1_dfm_5[49];
  assign FpAdd_8U_23U_if_3_if_and_tmp_1 = fsm_output[1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13592" *) FpAdd_8U_23U_int_mant_p1_2_lpi_1_dfm_5[49];
  assign FpAdd_8U_23U_if_3_if_and_tmp_2 = fsm_output[1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13593" *) FpAdd_8U_23U_int_mant_p1_3_lpi_1_dfm_5[49];
  assign FpAdd_8U_23U_if_3_if_and_tmp_3 = fsm_output[1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13594" *) FpAdd_8U_23U_int_mant_p1_lpi_1_dfm_5[49];
  assign FpAdd_8U_23U_a_right_shift_qelse_and_tmp = fsm_output[1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13596" *) _1344_;
  assign FpAdd_8U_23U_a_right_shift_qelse_and_tmp_1 = fsm_output[1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13598" *) _1346_;
  assign FpAdd_8U_23U_a_right_shift_qelse_and_tmp_2 = fsm_output[1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13600" *) _1348_;
  assign FpAdd_8U_23U_a_right_shift_qelse_and_tmp_3 = fsm_output[1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13602" *) _1350_;
  assign alu_loop_op_else_else_if_and_cse = fsm_output[1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13603" *) _1149_;
  assign alu_loop_op_else_else_if_and_1_cse = fsm_output[1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13604" *) cfg_alu_algo_1_sva_2[0];
  assign FpAdd_8U_23U_if_2_and_tmp = fsm_output[1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13605" *) reg_alu_loop_op_1_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_1_cse;
  assign FpAdd_8U_23U_if_2_and_tmp_1 = fsm_output[1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13606" *) reg_alu_loop_op_2_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_2_svs_1_cse;
  assign FpAdd_8U_23U_if_2_and_tmp_2 = fsm_output[1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13607" *) reg_alu_loop_op_3_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_1_svs_1_cse;
  assign FpAdd_8U_23U_if_2_and_tmp_3 = fsm_output[1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13608" *) reg_alu_loop_op_4_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_3_svs_1_cse;
  assign _0630_ = _1351_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13628" *) fsm_output[1];
  assign _0631_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13638" *) chn_alu_in_rsci_ld_core_psct_mx0c0;
  assign _0632_ = chn_alu_out_and_8_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13701" *) chn_alu_out_or_cse;
  assign _0633_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13720" *) _1804_;
  assign _0634_ = and_dcpl_30 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13728" *) and_dcpl_46;
  assign _0635_ = _0634_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13729" *) cfg_alu_src_1_sva_st_1;
  assign _0636_ = _0635_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13729" *) cfg_alu_src_rsci_d;
  assign _0637_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13729" *) _1806_;
  assign _0638_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13737" *) _1807_;
  assign _0639_ = _0500_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13763" *) _1356_;
  assign _0640_ = _0500_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13771" *) _1357_;
  assign _0641_ = _0500_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13779" *) _1358_;
  assign _0642_ = chn_alu_out_and_8_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13788" *) _1808_;
  assign _0643_ = _0642_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13788" *) mux_38_nl;
  assign _0644_ = and_dcpl_83 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13798" *) fsm_output[1];
  assign _0645_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13799" *) _1810_;
  assign _0646_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13809" *) _1359_;
  assign _0647_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13817" *) _1813_;
  assign _0648_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13960" *) _1814_;
  assign _0649_ = _0492_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14021" *) mux_59_nl;
  assign _0650_ = _0492_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14031" *) mux_61_nl;
  assign _0651_ = _0492_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14041" *) mux_63_nl;
  assign _0652_ = _0492_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14051" *) mux_65_nl;
  assign _0653_ = _0491_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14060" *) mux_67_nl;
  assign _0654_ = or_1087_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14088" *) main_stage_v_3;
  assign _0655_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14089" *) _1815_;
  assign _0656_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14097" *) FpAdd_8U_23U_o_expo_FpAdd_8U_23U_o_expo_or_2_cse;
  assign _0657_ = _0656_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14098" *) mux_74_nl;
  assign _0658_ = _0656_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14108" *) mux_80_nl;
  assign _0659_ = _0656_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14118" *) mux_86_nl;
  assign _0660_ = _0491_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14127" *) mux_92_nl;
  assign _0661_ = _0492_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14137" *) mux_94_nl;
  assign _0662_ = _0492_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14149" *) mux_96_nl;
  assign _0663_ = _0492_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14161" *) mux_98_nl;
  assign _0664_ = _0492_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14173" *) mux_100_nl;
  assign _0665_ = nand_109_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14183" *) FpAlu_8U_23U_nor_dfs_5;
  assign _0666_ = _0665_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14183" *) nor_430_cse;
  assign _0667_ = _0666_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14183" *) IsNaN_8U_23U_land_lpi_1_dfm_10;
  assign _0668_ = _1816_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14184" *) and_dcpl;
  assign _0669_ = _0668_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14184" *) or_1087_cse;
  assign _0670_ = _1364_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14192" *) IsNaN_8U_23U_land_lpi_1_dfm_10;
  assign _0671_ = _1817_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14193" *) FpAlu_8U_23U_nor_dfs_5;
  assign _0672_ = _0671_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14193" *) _1196_;
  assign _0673_ = _0672_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14193" *) _1365_;
  assign _0674_ = _1818_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14194" *) and_dcpl;
  assign _0675_ = _0674_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14194" *) or_1087_cse;
  assign _0676_ = alu_loop_op_3_FpAdd_8U_23U_if_4_if_acc_2_nl[7] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14229" *) alu_loop_op_3_FpMantRNE_49U_24U_else_and_1_tmp;
  assign _0677_ = alu_loop_op_2_FpAdd_8U_23U_if_4_if_acc_4_nl[7] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14231" *) alu_loop_op_2_FpMantRNE_49U_24U_else_and_2_tmp;
  assign _0678_ = alu_loop_op_1_FpAdd_8U_23U_if_4_if_acc_1_nl[7] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14233" *) alu_loop_op_1_FpMantRNE_49U_24U_else_and_tmp;
  assign _0679_ = alu_loop_op_4_FpAdd_8U_23U_if_4_if_acc_6_nl[7] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14235" *) alu_loop_op_4_FpMantRNE_49U_24U_else_and_3_tmp;
  assign _0680_ = _0666_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14260" *) IsNaN_8U_23U_land_3_lpi_1_dfm_10;
  assign _0681_ = _1819_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14261" *) and_dcpl;
  assign _0682_ = _0681_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14261" *) or_1087_cse;
  assign _0683_ = _1364_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14269" *) IsNaN_8U_23U_land_3_lpi_1_dfm_10;
  assign _0684_ = _1820_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14270" *) FpAlu_8U_23U_nor_dfs_5;
  assign _0685_ = _0684_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14270" *) _1196_;
  assign _0686_ = _0685_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14270" *) _1365_;
  assign _0687_ = _1821_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14271" *) and_dcpl;
  assign _0688_ = _0687_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14271" *) or_1087_cse;
  assign _0689_ = _0666_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14279" *) IsNaN_8U_23U_land_2_lpi_1_dfm_10;
  assign _0690_ = _1822_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14280" *) and_dcpl;
  assign _0691_ = _0690_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14280" *) or_1087_cse;
  assign _0692_ = _1364_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14288" *) IsNaN_8U_23U_land_2_lpi_1_dfm_10;
  assign _0693_ = _1823_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14289" *) FpAlu_8U_23U_nor_dfs_5;
  assign _0694_ = _0693_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14289" *) _1196_;
  assign _0695_ = _0694_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14289" *) _1365_;
  assign _0696_ = _1824_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14290" *) and_dcpl;
  assign _0697_ = _0696_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14290" *) or_1087_cse;
  assign _0698_ = _0666_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14298" *) IsNaN_8U_23U_land_1_lpi_1_dfm_10;
  assign _0699_ = _1825_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14299" *) and_dcpl;
  assign _0700_ = _0699_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14299" *) or_1087_cse;
  assign _0701_ = _1364_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14307" *) IsNaN_8U_23U_land_1_lpi_1_dfm_10;
  assign _0702_ = _1826_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14308" *) FpAlu_8U_23U_nor_dfs_5;
  assign _0703_ = _0702_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14308" *) _1196_;
  assign _0704_ = _0703_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14308" *) _1365_;
  assign _0705_ = _1827_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14309" *) and_dcpl;
  assign _0706_ = _0705_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14309" *) or_1087_cse;
  assign _0707_ = _1828_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14345" *) main_stage_v_4;
  assign _0708_ = _1829_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14346" *) or_1087_cse;
  assign _0709_ = _0708_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14346" *) core_wen;
  assign _0710_ = _0491_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14355" *) _1366_;
  assign _0711_ = or_1087_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14363" *) alu_loop_op_3_FpMantRNE_49U_24U_else_and_1_tmp;
  assign _0712_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14364" *) _1830_;
  assign _0713_ = _0712_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14364" *) _1207_;
  assign _0714_ = _0491_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14373" *) mux_128_nl;
  assign _0715_ = _1482_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14383" *) main_stage_v_4;
  assign _0716_ = _1831_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14383" *) or_1087_cse;
  assign _0717_ = _0716_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14383" *) core_wen;
  assign _0718_ = or_1087_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14402" *) alu_loop_op_2_FpMantRNE_49U_24U_else_and_2_tmp;
  assign _0719_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14403" *) _1832_;
  assign _0720_ = _0719_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14403" *) _1207_;
  assign _0721_ = _0491_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14412" *) mux_130_nl;
  assign _0722_ = or_1087_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14420" *) alu_loop_op_1_FpMantRNE_49U_24U_else_and_tmp;
  assign _0723_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14421" *) _1833_;
  assign _0724_ = _0723_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14421" *) _1207_;
  assign _0725_ = _0491_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14430" *) mux_131_nl;
  assign _0726_ = _0491_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14438" *) _1367_;
  assign _0727_ = _0491_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14446" *) _1368_;
  assign _0728_ = _1370_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14456" *) _1314_;
  assign _0729_ = _0728_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14456" *) main_stage_v_4;
  assign _0730_ = _0729_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14456" *) core_wen;
  assign _0731_ = _0730_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14456" *) or_1087_cse;
  assign _0732_ = _0491_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14464" *) _1371_;
  assign _0733_ = or_1087_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14482" *) alu_loop_op_4_FpMantRNE_49U_24U_else_and_3_tmp;
  assign _0734_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14483" *) _1838_;
  assign _0735_ = _0734_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14483" *) _1207_;
  assign _0736_ = _0491_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14492" *) mux_137_nl;
  assign _0737_ = _0491_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14500" *) _1372_;
  assign _0738_ = _0491_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14508" *) _1373_;
  assign _0739_ = mux_362_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14558" *) core_wen;
  assign _0740_ = _0656_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14569" *) _1221_;
  assign _0741_ = FpMantRNE_49U_24U_else_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14579" *) mux_145_nl;
  assign _0742_ = FpMantRNE_49U_24U_else_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14589" *) mux_146_nl;
  assign _0743_ = FpMantRNE_49U_24U_else_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14599" *) mux_147_nl;
  assign _0744_ = FpMantRNE_49U_24U_else_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14609" *) mux_148_nl;
  assign _0745_ = _0491_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14632" *) mux_150_nl;
  assign _0746_ = _0491_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14640" *) mux_152_nl;
  assign _0747_ = _0491_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14648" *) mux_154_nl;
  assign _0748_ = _0491_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14656" *) mux_156_nl;
  assign _0749_ = chn_alu_out_and_8_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14664" *) _1226_;
  assign _0750_ = _0749_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14664" *) mux_157_nl;
  assign _0751_ = _0749_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14686" *) mux_158_nl;
  assign _0752_ = _0749_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14694" *) mux_159_nl;
  assign _0753_ = _0749_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14702" *) mux_160_nl;
  assign _0754_ = _0520_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14788" *) _1374_;
  assign _0755_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14796" *) _1375_;
  assign _0756_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14805" *) _1376_;
  assign _0757_ = _0484_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14813" *) _1358_;
  assign _0758_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14821" *) _1843_;
  assign _0759_ = _0758_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14821" *) not_tmp_29;
  assign _0760_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14832" *) _1845_;
  assign _0761_ = _0760_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14832" *) not_tmp_29;
  assign _0762_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14843" *) _1847_;
  assign _0763_ = _0762_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14843" *) not_tmp_29;
  assign _0764_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14854" *) _1849_;
  assign _0765_ = _0764_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14854" *) not_tmp_29;
  assign _0766_ = _0512_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14880" *) _1377_;
  assign _0767_ = _0491_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14920" *) _1378_;
  assign _0768_ = _0491_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14940" *) _1379_;
  assign _0769_ = _0491_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14948" *) _1380_;
  assign _0770_ = _0491_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14966" *) _1381_;
  assign _0771_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14974" *) IntSaturation_33U_32U_IntSaturation_33U_32U_or_7_cse;
  assign _0772_ = _0771_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14975" *) mux_200_nl;
  assign _0773_ = _0771_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15000" *) mux_204_nl;
  assign _0774_ = _0771_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15011" *) mux_206_nl;
  assign _0775_ = _0771_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15022" *) mux_208_nl;
  assign _0776_ = _0492_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15055" *) mux_209_nl;
  assign _0777_ = _0492_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15065" *) mux_210_nl;
  assign _0778_ = _0492_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15075" *) mux_211_nl;
  assign _0779_ = _0492_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15085" *) mux_212_nl;
  assign _0780_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15095" *) _1382_;
  assign _0781_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15104" *) _1383_;
  assign _0782_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15113" *) _1384_;
  assign _0783_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15122" *) _1385_;
  assign _0784_ = FpAlu_8U_23U_mux1h_144_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15154" *) _1386_;
  assign _0785_ = FpAlu_8U_23U_mux1h_148_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15155" *) _1386_;
  assign _0786_ = _0616_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15163" *) FpAdd_8U_23U_is_a_greater_lor_1_lpi_1_dfm_1_mx0w0;
  assign _0787_ = _0786_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15163" *) main_stage_v_1;
  assign _0788_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15163" *) _1856_;
  assign _0789_ = _0616_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15173" *) FpAdd_8U_23U_is_a_greater_lor_2_lpi_1_dfm_1_mx0w0;
  assign _0790_ = _0789_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15173" *) main_stage_v_1;
  assign _0791_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15173" *) _1857_;
  assign _0792_ = _0616_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15183" *) FpAdd_8U_23U_is_a_greater_lor_3_lpi_1_dfm_1_mx0w0;
  assign _0793_ = _0792_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15183" *) main_stage_v_1;
  assign _0794_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15183" *) _1858_;
  assign _0795_ = _0616_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15193" *) FpAdd_8U_23U_is_a_greater_lor_lpi_1_dfm_1_mx0w0;
  assign _0796_ = _0795_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15193" *) main_stage_v_1;
  assign _0797_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15193" *) _1859_;
  assign _0798_ = _0491_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15228" *) mux_218_nl;
  assign _0799_ = _0491_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15236" *) mux_219_nl;
  assign _0800_ = _0491_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15258" *) mux_223_nl;
  assign _0801_ = _0491_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15278" *) mux_225_nl;
  assign _0802_ = _0491_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15286" *) mux_226_nl;
  assign _0803_ = or_963_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15294" *) core_wen;
  assign _0804_ = _0803_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15295" *) _1387_;
  assign _0805_ = _0804_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15295" *) _0009_;
  assign _0806_ = _0805_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15296" *) cfg_alu_algo_rsc_triosy_obj_bawt;
  assign _0807_ = _0806_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15296" *) or_1050_cse;
  assign _0808_ = _0807_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15296" *) and_dcpl_349;
  assign _0809_ = _0808_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15296" *) cfg_alu_bypass_rsc_triosy_obj_bawt;
  assign _0810_ = _0809_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15297" *) _1190_;
  assign _0811_ = _0810_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15297" *) or_1087_cse;
  assign _0812_ = _0811_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15297" *) main_stage_v_1;
  assign _0813_ = _1388_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15305" *) core_wen;
  assign _0814_ = _0813_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15306" *) _0009_;
  assign _0815_ = _0814_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15306" *) and_dcpl_2;
  assign _0816_ = _0815_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15306" *) and_dcpl_3;
  assign _0817_ = _0816_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15306" *) _1190_;
  assign _0818_ = _0817_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15307" *) main_stage_v_1;
  assign _0819_ = _0818_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15307" *) or_1087_cse;
  assign _0820_ = _0803_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15316" *) _1389_;
  assign _0821_ = _0820_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15316" *) _0009_;
  assign _0822_ = _0821_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15317" *) cfg_alu_algo_rsc_triosy_obj_bawt;
  assign _0823_ = _0822_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15317" *) or_1050_cse;
  assign _0824_ = _0823_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15317" *) and_dcpl_349;
  assign _0825_ = _0824_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15317" *) cfg_alu_bypass_rsc_triosy_obj_bawt;
  assign _0826_ = _0825_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15318" *) _1190_;
  assign _0827_ = _0826_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15318" *) or_1087_cse;
  assign _0828_ = _0827_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15318" *) main_stage_v_1;
  assign _0829_ = _1390_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15326" *) core_wen;
  assign _0830_ = _0829_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15327" *) _0009_;
  assign _0831_ = _0830_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15327" *) and_dcpl_2;
  assign _0832_ = _0831_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15327" *) and_dcpl_3;
  assign _0833_ = _0832_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15327" *) _1190_;
  assign _0834_ = _0833_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15328" *) main_stage_v_1;
  assign _0835_ = _0834_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15328" *) or_1087_cse;
  assign _0836_ = or_1087_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15337" *) _1190_;
  assign _0837_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15338" *) _1862_;
  assign _0838_ = _0837_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15338" *) not_tmp_232;
  assign _0839_ = _0803_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15349" *) _1391_;
  assign _0840_ = _0839_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15349" *) _0009_;
  assign _0841_ = _0840_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15350" *) cfg_alu_algo_rsc_triosy_obj_bawt;
  assign _0842_ = _0841_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15350" *) or_1050_cse;
  assign _0843_ = _0842_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15350" *) and_dcpl_349;
  assign _0844_ = _0843_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15350" *) cfg_alu_bypass_rsc_triosy_obj_bawt;
  assign _0845_ = _0844_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15351" *) _1190_;
  assign _0846_ = _0845_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15351" *) or_1087_cse;
  assign _0847_ = _0846_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15351" *) main_stage_v_1;
  assign _0848_ = _1392_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15359" *) or_963_cse;
  assign _0849_ = _0848_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15359" *) core_wen;
  assign _0850_ = _0849_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15360" *) _0009_;
  assign _0851_ = _0850_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15360" *) cfg_alu_algo_rsc_triosy_obj_bawt;
  assign _0852_ = _0851_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15360" *) cfg_alu_op_rsc_triosy_obj_bawt;
  assign _0853_ = _0852_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15361" *) and_dcpl_3;
  assign _0854_ = _0853_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15361" *) _1190_;
  assign _0855_ = _0854_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15361" *) main_stage_v_1;
  assign _0856_ = _0855_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15362" *) or_1087_cse;
  assign _0857_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15370" *) _0009_;
  assign _0858_ = _0857_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15370" *) or_963_cse;
  assign _0859_ = _0858_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15371" *) and_dcpl_2;
  assign _0860_ = _0859_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15371" *) or_1050_cse;
  assign _0861_ = _0860_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15371" *) and_dcpl_3;
  assign _0862_ = _0861_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15371" *) _1190_;
  assign _0863_ = _0862_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15372" *) main_stage_v_1;
  assign _0864_ = _0863_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15372" *) _1393_;
  assign _0865_ = _1394_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15381" *) core_wen;
  assign _0866_ = _0865_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15382" *) _0009_;
  assign _0867_ = _0866_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15382" *) cfg_alu_algo_rsc_triosy_obj_bawt;
  assign _0868_ = _0867_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15382" *) and_dcpl_349;
  assign _0869_ = _0868_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15383" *) cfg_alu_bypass_rsc_triosy_obj_bawt;
  assign _0870_ = _0869_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15383" *) _1190_;
  assign _0871_ = _0870_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15383" *) main_stage_v_1;
  assign _0872_ = _0871_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15384" *) or_1087_cse;
  assign _0873_ = _0484_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15432" *) _1395_;
  assign _0874_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15475" *) _1396_;
  assign _0875_ = _0874_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15475" *) _1397_;
  assign _0876_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15483" *) IsNaN_8U_23U_2_IsNaN_8U_23U_4_or_2_cse;
  assign _0877_ = _0876_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15484" *) _1398_;
  assign _0878_ = _0876_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15495" *) _1399_;
  assign _0879_ = _0535_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15506" *) _1400_;
  assign _0880_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15534" *) _1871_;
  assign _0881_ = _0880_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15534" *) _1401_;
  assign _0882_ = _1402_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15567" *) FpAdd_8U_23U_FpAdd_8U_23U_nor_5_m1c;
  assign FpAdd_8U_23U_and_nl = _0882_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15567" *) FpAlu_8U_23U_nor_dfs_6;
  assign _0883_ = FpAdd_8U_23U_and_tmp_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15569" *) _1403_;
  assign _0884_ = _0883_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15569" *) FpAdd_8U_23U_FpAdd_8U_23U_nor_5_m1c;
  assign FpAdd_8U_23U_and_6_nl = _0884_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15569" *) FpAlu_8U_23U_nor_dfs_6;
  assign _0885_ = FpAdd_8U_23U_is_inf_1_lpi_1_dfm_8 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15571" *) FpAdd_8U_23U_FpAdd_8U_23U_nor_5_m1c;
  assign FpAdd_8U_23U_and_28_nl = _0885_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15571" *) FpAlu_8U_23U_nor_dfs_6;
  assign _0886_ = IsNaN_8U_23U_1_land_1_lpi_1_dfm_9 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15573" *) _1404_;
  assign FpAdd_8U_23U_and_9_nl = _0886_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15573" *) FpAlu_8U_23U_nor_dfs_6;
  assign _0887_ = _1405_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15587" *) FpAdd_8U_23U_FpAdd_8U_23U_nor_7_m1c;
  assign FpAdd_8U_23U_and_29_nl = _0887_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15587" *) FpAlu_8U_23U_nor_dfs_6;
  assign _0888_ = FpAdd_8U_23U_and_1_tmp_3 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15589" *) _1406_;
  assign _0889_ = _0888_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15589" *) FpAdd_8U_23U_FpAdd_8U_23U_nor_7_m1c;
  assign FpAdd_8U_23U_and_13_nl = _0889_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15589" *) FpAlu_8U_23U_nor_dfs_6;
  assign _0890_ = FpAdd_8U_23U_is_inf_2_lpi_1_dfm_8 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15591" *) FpAdd_8U_23U_FpAdd_8U_23U_nor_7_m1c;
  assign FpAdd_8U_23U_and_30_nl = _0890_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15591" *) FpAlu_8U_23U_nor_dfs_6;
  assign _0891_ = IsNaN_8U_23U_1_land_2_lpi_1_dfm_9 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15593" *) _1407_;
  assign FpAdd_8U_23U_and_15_nl = _0891_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15593" *) FpAlu_8U_23U_nor_dfs_6;
  assign _0892_ = and_486_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15616" *) _1408_;
  assign and_500_nl = _1921_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15671" *) mux_69_nl;
  assign and_499_nl = _1957_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15698" *) mux_75_nl;
  assign and_498_nl = _1991_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15725" *) mux_81_nl;
  assign and_497_nl = _2031_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15754" *) mux_87_nl;
  assign _0893_ = cfg_alu_algo_1_sva_st_25[1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15775" *) alu_loop_op_1_FpMantRNE_49U_24U_else_and_svs_st_2;
  assign _0894_ = cfg_alu_algo_1_sva_st_25[1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15783" *) alu_loop_op_2_FpMantRNE_49U_24U_else_and_2_svs_st_2;
  assign _0895_ = cfg_alu_algo_1_sva_st_25[1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15791" *) alu_loop_op_3_FpMantRNE_49U_24U_else_and_1_svs_st_2;
  assign _0896_ = cfg_alu_algo_1_sva_st_25[1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15799" *) alu_loop_op_4_FpMantRNE_49U_24U_else_and_3_svs_st_2;
  assign and_218_nl = _1441_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15858" *) and_dcpl_37;
  assign _0897_ = _1441_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15859" *) main_stage_v_4;
  assign _0898_ = _0897_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15859" *) or_1087_cse;
  assign and_220_nl = _0898_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15859" *) _1314_;
  assign and_496_nl = alu_loop_op_1_FpMantRNE_49U_24U_else_and_tmp & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15868" *) _1442_;
  assign and_495_nl = alu_loop_op_2_FpMantRNE_49U_24U_else_and_2_tmp & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15871" *) _1442_;
  assign and_494_nl = alu_loop_op_3_FpMantRNE_49U_24U_else_and_1_tmp & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15874" *) _1442_;
  assign and_493_nl = alu_loop_op_4_FpMantRNE_49U_24U_else_and_3_tmp & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15877" *) _1442_;
  assign _0899_ = FpAlu_8U_23U_equal_tmp_22 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15887" *) _2130_;
  assign _0900_ = FpAlu_8U_23U_equal_tmp_22 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15897" *) _2141_;
  assign _0901_ = FpAlu_8U_23U_equal_tmp_22 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15907" *) _2152_;
  assign _0902_ = FpAlu_8U_23U_equal_tmp_22 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15917" *) _2163_;
  assign _0903_ = AluOut_data_0_0_sva_9 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15943" *) _1447_;
  assign _0904_ = FpAlu_8U_23U_mux1h_33_itm_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15950" *) _1449_;
  assign _0905_ = FpAlu_8U_23U_mux1h_152_itm_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15952" *) _1450_;
  assign _0906_ = AluOut_data_1_0_sva_10 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15954" *) _1451_;
  assign FpAlu_8U_23U_and_9_nl = FpAlu_8U_23U_mux1h_152_itm_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16008" *) _1448_;
  assign FpAlu_8U_23U_and_nl = FpAlu_8U_23U_mux1h_33_itm_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16009" *) _1448_;
  assign _0907_ = _1466_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16047" *) FpAlu_8U_23U_and_52_m1c;
  assign _0908_ = IsNaN_8U_23U_1_land_1_lpi_1_dfm_mx0w0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16047" *) FpAlu_8U_23U_and_36_m1c;
  assign _0909_ = FpAdd_8U_23U_is_a_greater_lor_1_lpi_1_dfm_1_mx0w0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16049" *) FpAlu_8U_23U_and_52_m1c;
  assign _0910_ = IsNaN_8U_23U_land_1_lpi_1_dfm_8 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16049" *) FpAlu_8U_23U_nor_dfs_mx0w0;
  assign _0911_ = _1467_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16055" *) FpAlu_8U_23U_and_56_m1c;
  assign _0912_ = IsNaN_8U_23U_1_land_2_lpi_1_dfm_mx0w0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16055" *) FpAlu_8U_23U_and_38_m1c;
  assign _0913_ = FpAdd_8U_23U_is_a_greater_lor_2_lpi_1_dfm_1_mx0w0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16057" *) FpAlu_8U_23U_and_56_m1c;
  assign _0914_ = IsNaN_8U_23U_land_2_lpi_1_dfm_8 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16057" *) FpAlu_8U_23U_nor_dfs_mx0w0;
  assign _0915_ = alu_loop_op_else_mux_1_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16070" *) and_dcpl_208;
  assign _0916_ = alu_loop_op_else_mux_2_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16074" *) and_dcpl_208;
  assign AluOut_data_and_7_nl = alu_loop_op_else_mux_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16077" *) and_dcpl_208;
  assign _0917_ = FpAlu_8U_23U_mux_21_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16080" *) and_dcpl_208;
  assign _0918_ = FpAlu_8U_23U_mux_20_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16084" *) and_dcpl_208;
  assign AluOut_data_and_3_nl = alu_loop_op_else_mux_3_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16087" *) and_dcpl_208;
  assign _0919_ = _1468_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16115" *) FpAlu_8U_23U_and_40_m1c;
  assign _0920_ = IsNaN_8U_23U_1_land_lpi_1_dfm_mx0w0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16115" *) FpAlu_8U_23U_and_24_m1c;
  assign FpAlu_8U_23U_and_74_nl = _2300_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16116" *) and_dcpl_207;
  assign _0921_ = FpAdd_8U_23U_is_a_greater_lor_lpi_1_dfm_1_mx0w0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16118" *) FpAlu_8U_23U_and_40_m1c;
  assign _0922_ = IsNaN_8U_23U_land_lpi_1_dfm_8 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16118" *) FpAlu_8U_23U_nor_dfs_mx0w0;
  assign FpAlu_8U_23U_and_75_nl = _2301_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16119" *) and_dcpl_207;
  assign FpAlu_8U_23U_and_76_nl = FpAlu_8U_23U_equal_tmp_mx0w0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16120" *) and_dcpl_207;
  assign FpAlu_8U_23U_and_77_nl = FpAlu_8U_23U_equal_tmp_2_mx0w0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16121" *) and_dcpl_207;
  assign FpAlu_8U_23U_and_80_nl = alu_loop_op_else_mux_5_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16124" *) and_dcpl_214;
  assign FpAlu_8U_23U_and_81_nl = alu_loop_op_else_mux_4_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16127" *) and_dcpl_214;
  assign _0923_ = _1469_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16129" *) FpAlu_8U_23U_and_48_m1c;
  assign _0924_ = IsNaN_8U_23U_1_land_3_lpi_1_dfm_mx0w0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16129" *) FpAlu_8U_23U_and_34_m1c;
  assign FpAlu_8U_23U_and_66_nl = _2302_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16130" *) and_297_m1c;
  assign _0925_ = FpAdd_8U_23U_is_a_greater_lor_3_lpi_1_dfm_1_mx0w0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16132" *) FpAlu_8U_23U_and_48_m1c;
  assign _0926_ = IsNaN_8U_23U_land_3_lpi_1_dfm_8 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16132" *) FpAlu_8U_23U_nor_dfs_mx0w0;
  assign FpAlu_8U_23U_and_67_nl = _2303_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16133" *) and_297_m1c;
  assign FpAlu_8U_23U_and_68_nl = FpAlu_8U_23U_equal_tmp_mx0w0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16134" *) and_297_m1c;
  assign FpAlu_8U_23U_and_69_nl = FpAlu_8U_23U_equal_tmp_2_mx0w0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16135" *) and_297_m1c;
  assign FpAlu_8U_23U_and_72_nl = FpAlu_8U_23U_equal_tmp_1_mx0w0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16136" *) and_dcpl_214;
  assign FpAlu_8U_23U_and_73_nl = alu_loop_op_else_equal_tmp_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16137" *) and_dcpl_214;
  assign and_74_nl = or_16_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16138" *) or_tmp_386;
  assign _0927_ = main_stage_v_1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16141" *) _1470_;
  assign _0928_ = main_stage_v_1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16159" *) mux_287_nl;
  assign _0929_ = main_stage_v_1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16163" *) _1472_;
  assign _0930_ = main_stage_v_1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16170" *) mux_300_nl;
  assign _0931_ = main_stage_v_1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16174" *) _1473_;
  assign _0932_ = AluOut_data_2_0_sva_10 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16264" *) and_dcpl_127;
  assign _0933_ = IntSaturation_33U_32U_o_31_1_3_lpi_1_dfm_1[30] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16264" *) alu_loop_bypass_if_and_7_cse;
  assign _0934_ = IntSaturation_33U_32U_o_31_1_lpi_1_dfm_1[30] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16264" *) alu_loop_bypass_if_and_7_cse;
  assign _0935_ = IntSaturation_33U_32U_o_31_1_2_lpi_1_dfm_1[30] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16264" *) alu_loop_bypass_if_and_7_cse;
  assign _0936_ = IntSaturation_33U_32U_o_31_1_1_lpi_1_dfm_1[30] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16264" *) alu_loop_bypass_if_and_7_cse;
  assign _0937_ = alu_loop_op_else_else_else_else_ac_int_cctor_2_sva[0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16264" *) AluOut_data_and_7_nl;
  assign _0938_ = alu_loop_op_else_else_else_else_ac_int_cctor_1_sva[0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16264" *) AluOut_data_and_3_nl;
  assign _0939_ = IsNaN_8U_23U_2_IsNaN_8U_23U_2_nor_2_itm_mx0w0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16264" *) and_dcpl_243;
  assign _0940_ = IsNaN_8U_23U_2_IsNaN_8U_23U_2_nor_1_itm_mx0w0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16264" *) and_dcpl_243;
  assign _0941_ = IsNaN_8U_23U_2_IsNaN_8U_23U_2_nor_itm_mx0w0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16264" *) and_dcpl_243;
  assign _0942_ = IsNaN_8U_23U_2_IsNaN_8U_23U_2_nor_3_itm_mx0w0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16264" *) and_dcpl_243;
  assign _0943_ = alu_loop_op_mux_204_mx1w1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16265" *) and_220_nl;
  assign _0944_ = FpAlu_8U_23U_and_9_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16265" *) alu_loop_bypass_if_and_6_cse;
  assign _0945_ = FpAlu_8U_23U_and_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16265" *) alu_loop_bypass_if_and_6_cse;
  assign _0946_ = FpAlu_8U_23U_and_6_itm_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16265" *) alu_loop_bypass_if_and_6_cse;
  assign _0947_ = FpAlu_8U_23U_and_3_itm_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16265" *) alu_loop_bypass_if_and_6_cse;
  assign _0948_ = alu_loop_op_else_if_qr_31_0_2_lpi_1_dfm_mx0[0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16265" *) AluOut_data_or_2_nl;
  assign _0949_ = alu_loop_op_else_if_qr_31_0_1_lpi_1_dfm_mx0[0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16265" *) AluOut_data_or_3_nl;
  assign _0950_ = IsNaN_8U_23U_2_IsNaN_8U_23U_2_nor_itm_mx0w0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16265" *) and_dcpl_239;
  assign _0951_ = IsNaN_8U_23U_4_IsNaN_8U_23U_4_nand_3_itm_mx0w2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16265" *) and_dcpl_239;
  assign _0952_ = IsNaN_8U_23U_4_IsNaN_8U_23U_4_nand_2_itm_mx0w2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16265" *) and_dcpl_239;
  assign _0953_ = IsNaN_8U_23U_2_nor_2_mx0w0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16265" *) and_dcpl_239;
  assign _0954_ = reg_AluIn_data_sva_4_94_64_1_itm[0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16266" *) and_218_nl;
  assign _0955_ = AluIn_data_sva_128[95] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16266" *) and_dcpl_170;
  assign _0956_ = AluIn_data_sva_128[127] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16266" *) and_dcpl_170;
  assign _0957_ = AluIn_data_sva_128[63] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16266" *) and_dcpl_170;
  assign _0958_ = AluIn_data_sva_128[31] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16266" *) and_dcpl_170;
  assign _0959_ = _1172_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16266" *) AluOut_data_or_1_nl;
  assign _0960_ = _1173_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16266" *) AluOut_data_or_nl;
  assign _0961_ = IsNaN_8U_23U_2_IsNaN_8U_23U_2_nor_3_itm_mx0w0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16266" *) and_dcpl_236;
  assign _0962_ = IsNaN_8U_23U_2_IsNaN_8U_23U_2_nor_2_itm_mx0w0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16266" *) and_dcpl_236;
  assign _0963_ = IsNaN_8U_23U_2_IsNaN_8U_23U_2_nor_1_itm_mx0w0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16266" *) and_dcpl_236;
  assign _0964_ = IsNaN_8U_23U_2_IsNaN_8U_23U_2_nor_itm_mx0w0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16266" *) and_dcpl_236;
  assign _0965_ = IsNaN_8U_23U_2_IsNaN_8U_23U_2_nor_2_itm_mx0w0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16278" *) and_dcpl_225;
  assign _0966_ = IsNaN_8U_23U_2_IsNaN_8U_23U_2_nor_3_itm_mx0w0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16278" *) and_dcpl_225;
  assign _0967_ = IsNaN_8U_23U_2_IsNaN_8U_23U_2_nor_1_itm_mx0w0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16278" *) and_dcpl_225;
  assign _0968_ = IsNaN_8U_23U_2_IsNaN_8U_23U_2_nor_itm_mx0w0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16278" *) and_dcpl_225;
  assign _0969_ = alu_loop_op_2_FpAdd_8U_23U_IsZero_8U_23U_or_itm_3 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16278" *) and_dcpl_231;
  assign _0970_ = IsNaN_8U_23U_4_nor_3_itm_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16278" *) and_dcpl_231;
  assign _0971_ = FpCmp_8U_23U_false_o_1_lpi_1_dfm_7_30_0_1[0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16278" *) FpAlu_8U_23U_equal_tmp_29;
  assign _0972_ = FpCmp_8U_23U_false_o_2_lpi_1_dfm_8_30_0_1[0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16278" *) FpAlu_8U_23U_equal_tmp_29;
  assign _0973_ = FpCmp_8U_23U_false_o_1_lpi_1_dfm_1_mx0[31] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16278" *) FpAlu_8U_23U_equal_tmp_2_mx0w0;
  assign _0974_ = FpCmp_8U_23U_false_o_2_lpi_1_dfm_2[31] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16278" *) FpAlu_8U_23U_equal_tmp_2_mx0w0;
  assign _0975_ = IsNaN_8U_23U_2_IsNaN_8U_23U_2_nor_itm_mx0w0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16279" *) and_dcpl_222;
  assign _0976_ = IsNaN_8U_23U_2_IsNaN_8U_23U_2_nor_1_itm_mx0w0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16279" *) and_dcpl_222;
  assign _0977_ = IsNaN_8U_23U_4_IsNaN_8U_23U_4_nand_3_itm_mx0w2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16279" *) and_dcpl_222;
  assign _0978_ = IsNaN_8U_23U_4_IsNaN_8U_23U_4_nand_2_itm_mx0w2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16279" *) and_dcpl_222;
  assign _0979_ = alu_loop_op_2_FpAdd_8U_23U_IsZero_8U_23U_or_itm_mx0w0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16279" *) and_dcpl_229;
  assign _0980_ = alu_loop_op_1_FpAdd_8U_23U_IsZero_8U_23U_or_itm_mx0w2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16279" *) and_dcpl_229;
  assign _0981_ = AluOut_data_0_0_sva_11 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16279" *) FpAlu_8U_23U_equal_tmp_23;
  assign _0982_ = AluOut_data_1_0_sva_12 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16279" *) FpAlu_8U_23U_equal_tmp_23;
  assign _0983_ = FpCmp_8U_23U_true_o_1_lpi_1_dfm_1_mx0[31] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16279" *) FpAlu_8U_23U_equal_tmp_mx0w0;
  assign _0984_ = FpCmp_8U_23U_true_o_2_lpi_1_dfm_1_mx0[31] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16279" *) FpAlu_8U_23U_equal_tmp_mx0w0;
  assign _0985_ = IsNaN_8U_23U_2_IsNaN_8U_23U_2_nor_3_itm & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16280" *) and_dcpl_81;
  assign _0986_ = IsNaN_8U_23U_2_IsNaN_8U_23U_2_nor_itm & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16280" *) and_dcpl_81;
  assign _0987_ = IsNaN_8U_23U_2_IsNaN_8U_23U_2_nor_2_itm & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16280" *) and_dcpl_81;
  assign _0988_ = IsNaN_8U_23U_2_IsNaN_8U_23U_2_nor_1_itm & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16280" *) and_dcpl_81;
  assign _0989_ = IsNaN_8U_23U_4_nor_3_itm_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16280" *) and_dcpl_227;
  assign _0990_ = IsNaN_8U_23U_2_IsNaN_8U_23U_2_nor_itm & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16280" *) and_dcpl_227;
  assign _0991_ = FpCmp_8U_23U_true_o_1_lpi_1_dfm_7_30_0_1[0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16280" *) FpAlu_8U_23U_equal_tmp_26;
  assign _0992_ = FpCmp_8U_23U_true_o_2_lpi_1_dfm_7_30_0_1[0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16280" *) FpAlu_8U_23U_equal_tmp_26;
  assign _0993_ = AluIn_data_sva_127[31] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16280" *) FpAlu_8U_23U_or_146_nl;
  assign _0994_ = AluIn_data_sva_127[63] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16280" *) FpAlu_8U_23U_or_148_nl;
  assign _0995_ = IsNaN_8U_23U_2_IsNaN_8U_23U_2_nor_3_itm_mx0w0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16281" *) and_dcpl_219;
  assign _0996_ = IsNaN_8U_23U_2_IsNaN_8U_23U_2_nor_itm_mx0w0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16281" *) and_dcpl_219;
  assign _0997_ = IsNaN_8U_23U_2_IsNaN_8U_23U_2_nor_2_itm_mx0w0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16281" *) and_dcpl_219;
  assign _0998_ = IsNaN_8U_23U_2_IsNaN_8U_23U_2_nor_1_itm_mx0w0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16281" *) and_dcpl_219;
  assign _0999_ = IsNaN_8U_23U_2_nor_3_mx0w0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16281" *) and_dcpl_222;
  assign _1000_ = IsNaN_8U_23U_2_nor_2_mx0w0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16281" *) and_dcpl_222;
  assign _1001_ = reg_AluIn_data_sva_4_30_0_1_itm[0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16281" *) FpAlu_8U_23U_nor_dfs_6;
  assign _1002_ = reg_AluIn_data_sva_4_62_32_1_itm[0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16281" *) FpAlu_8U_23U_nor_dfs_6;
  assign _1003_ = else_AluOp_data_0_lpi_1_dfm_mx0[31] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16281" *) FpAlu_8U_23U_or_145_nl;
  assign _1004_ = else_AluOp_data_1_lpi_1_dfm_mx0[31] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16281" *) FpAlu_8U_23U_or_147_nl;
  assign _1005_ = FpCmp_8U_23U_false_o_3_lpi_1_dfm_8_30_0_1[0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16294" *) FpAlu_8U_23U_and_31_m1c;
  assign _1006_ = FpCmp_8U_23U_false_o_lpi_1_dfm_9_30_0_1[0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16294" *) FpAlu_8U_23U_and_45_cse;
  assign _1007_ = AluOut_data_2_0_lpi_1_dfm_3 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16295" *) FpAlu_8U_23U_and_30_cse;
  assign _1008_ = FpAlu_8U_23U_o_0_lpi_1_dfm_4 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16295" *) FpAlu_8U_23U_and_44_cse;
  assign _1009_ = AluOut_data_2_0_sva_11 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16296" *) FpAlu_8U_23U_equal_tmp_23;
  assign _1010_ = FpAlu_8U_23U_o_0_sva_9 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16296" *) FpAlu_8U_23U_equal_tmp_23;
  assign _1011_ = FpCmp_8U_23U_true_o_3_lpi_1_dfm_7_30_0_1[0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16297" *) FpAlu_8U_23U_equal_tmp_26;
  assign _1012_ = FpCmp_8U_23U_true_o_lpi_1_dfm_7_30_0_1[0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16297" *) FpAlu_8U_23U_equal_tmp_26;
  assign _1013_ = reg_AluIn_data_sva_4_94_64_1_itm[0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16298" *) FpAlu_8U_23U_nor_dfs_6;
  assign _1014_ = reg_AluIn_data_sva_4_126_96_1_itm[0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16298" *) FpAlu_8U_23U_nor_dfs_6;
  assign _1015_ = alu_loop_op_else_else_else_else_ac_int_cctor_sva[0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16313" *) FpAlu_8U_23U_and_81_nl;
  assign _1016_ = alu_loop_op_else_else_else_else_ac_int_cctor_3_sva[0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16313" *) FpAlu_8U_23U_and_73_nl;
  assign _1017_ = FpAlu_8U_23U_o_0_sva_2_mx0w0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16314" *) FpAlu_8U_23U_and_80_nl;
  assign _1018_ = AluOut_data_2_0_sva_3_mx0w0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16314" *) FpAlu_8U_23U_and_72_nl;
  assign _1019_ = alu_loop_op_else_if_qr_31_0_lpi_1_dfm_mx0[0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16315" *) FpAlu_8U_23U_or_cse;
  assign _1020_ = alu_loop_op_else_if_qr_31_0_3_lpi_1_dfm_mx0[0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16315" *) FpAlu_8U_23U_or_cse;
  assign _1021_ = FpCmp_8U_23U_false_o_lpi_1_dfm_1_mx0[31] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16316" *) FpAlu_8U_23U_and_77_nl;
  assign _1022_ = FpCmp_8U_23U_false_o_3_lpi_1_dfm_1_mx0[31] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16316" *) FpAlu_8U_23U_and_69_nl;
  assign _1023_ = FpCmp_8U_23U_true_o_lpi_1_dfm_1_mx0[31] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16317" *) FpAlu_8U_23U_and_76_nl;
  assign _1024_ = FpCmp_8U_23U_true_o_3_lpi_1_dfm_1_mx0[31] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16317" *) FpAlu_8U_23U_and_68_nl;
  assign _1025_ = AluIn_data_sva_127[127] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16318" *) FpAlu_8U_23U_and_75_nl;
  assign _1026_ = AluIn_data_sva_127[95] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16318" *) FpAlu_8U_23U_and_67_nl;
  assign _1027_ = else_AluOp_data_3_lpi_1_dfm_mx0[31] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16319" *) FpAlu_8U_23U_and_74_nl;
  assign _1028_ = else_AluOp_data_2_lpi_1_dfm_mx0[31] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16319" *) FpAlu_8U_23U_and_66_nl;
  assign _1029_ = reg_AluIn_data_sva_4_30_0_1_itm[22:1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16330" *) { or_dcpl, or_dcpl, or_dcpl, or_dcpl, or_dcpl, or_dcpl, or_dcpl, or_dcpl, or_dcpl, or_dcpl, or_dcpl, or_dcpl, or_dcpl, or_dcpl, or_dcpl, or_dcpl, or_dcpl, or_dcpl, or_dcpl, or_dcpl, or_dcpl, or_dcpl };
  assign _1030_ = reg_AluIn_data_sva_4_62_32_1_itm[22:1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16330" *) { or_dcpl, or_dcpl, or_dcpl, or_dcpl, or_dcpl, or_dcpl, or_dcpl, or_dcpl, or_dcpl, or_dcpl, or_dcpl, or_dcpl, or_dcpl, or_dcpl, or_dcpl, or_dcpl, or_dcpl, or_dcpl, or_dcpl, or_dcpl, or_dcpl, or_dcpl };
  assign _1031_ = reg_AluIn_data_sva_4_126_96_1_itm[22:1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16330" *) { io_read_cfg_alu_bypass_rsc_svs_8, io_read_cfg_alu_bypass_rsc_svs_8, io_read_cfg_alu_bypass_rsc_svs_8, io_read_cfg_alu_bypass_rsc_svs_8, io_read_cfg_alu_bypass_rsc_svs_8, io_read_cfg_alu_bypass_rsc_svs_8, io_read_cfg_alu_bypass_rsc_svs_8, io_read_cfg_alu_bypass_rsc_svs_8, io_read_cfg_alu_bypass_rsc_svs_8, io_read_cfg_alu_bypass_rsc_svs_8, io_read_cfg_alu_bypass_rsc_svs_8, io_read_cfg_alu_bypass_rsc_svs_8, io_read_cfg_alu_bypass_rsc_svs_8, io_read_cfg_alu_bypass_rsc_svs_8, io_read_cfg_alu_bypass_rsc_svs_8, io_read_cfg_alu_bypass_rsc_svs_8, io_read_cfg_alu_bypass_rsc_svs_8, io_read_cfg_alu_bypass_rsc_svs_8, io_read_cfg_alu_bypass_rsc_svs_8, io_read_cfg_alu_bypass_rsc_svs_8, io_read_cfg_alu_bypass_rsc_svs_8, io_read_cfg_alu_bypass_rsc_svs_8 };
  assign _1032_ = FpCmp_8U_23U_false_o_3_lpi_1_dfm_8_30_0_1[22:1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16330" *) { FpAlu_8U_23U_and_31_m1c, FpAlu_8U_23U_and_31_m1c, FpAlu_8U_23U_and_31_m1c, FpAlu_8U_23U_and_31_m1c, FpAlu_8U_23U_and_31_m1c, FpAlu_8U_23U_and_31_m1c, FpAlu_8U_23U_and_31_m1c, FpAlu_8U_23U_and_31_m1c, FpAlu_8U_23U_and_31_m1c, FpAlu_8U_23U_and_31_m1c, FpAlu_8U_23U_and_31_m1c, FpAlu_8U_23U_and_31_m1c, FpAlu_8U_23U_and_31_m1c, FpAlu_8U_23U_and_31_m1c, FpAlu_8U_23U_and_31_m1c, FpAlu_8U_23U_and_31_m1c, FpAlu_8U_23U_and_31_m1c, FpAlu_8U_23U_and_31_m1c, FpAlu_8U_23U_and_31_m1c, FpAlu_8U_23U_and_31_m1c, FpAlu_8U_23U_and_31_m1c, FpAlu_8U_23U_and_31_m1c };
  assign _1033_ = reg_AluIn_data_sva_4_94_64_1_itm[22:1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16330" *) { or_dcpl, or_dcpl, or_dcpl, or_dcpl, or_dcpl, or_dcpl, or_dcpl, or_dcpl, or_dcpl, or_dcpl, or_dcpl, or_dcpl, or_dcpl, or_dcpl, or_dcpl, or_dcpl, or_dcpl, or_dcpl, or_dcpl, or_dcpl, or_dcpl, or_dcpl };
  assign _1034_ = AluOut_data_2_22_1_lpi_1_dfm_3 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16331" *) { asn_267, asn_267, asn_267, asn_267, asn_267, asn_267, asn_267, asn_267, asn_267, asn_267, asn_267, asn_267, asn_267, asn_267, asn_267, asn_267, asn_267, asn_267, asn_267, asn_267, asn_267, asn_267 };
  assign _1035_ = IntSaturation_33U_32U_slc_IntSaturation_33U_32U_o_31_1_2_21_0_itm_4 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16331" *) { asn_267, asn_267, asn_267, asn_267, asn_267, asn_267, asn_267, asn_267, asn_267, asn_267, asn_267, asn_267, asn_267, asn_267, asn_267, asn_267, asn_267, asn_267, asn_267, asn_267, asn_267, asn_267 };
  assign _1036_ = IntSaturation_33U_32U_slc_IntSaturation_33U_32U_o_31_1_21_0_itm_4 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16331" *) { asn_267, asn_267, asn_267, asn_267, asn_267, asn_267, asn_267, asn_267, asn_267, asn_267, asn_267, asn_267, asn_267, asn_267, asn_267, asn_267, asn_267, asn_267, asn_267, asn_267, asn_267, asn_267 };
  assign _1037_ = AluOut_data_2_22_1_lpi_1_dfm_3 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16331" *) { FpAlu_8U_23U_and_30_cse, FpAlu_8U_23U_and_30_cse, FpAlu_8U_23U_and_30_cse, FpAlu_8U_23U_and_30_cse, FpAlu_8U_23U_and_30_cse, FpAlu_8U_23U_and_30_cse, FpAlu_8U_23U_and_30_cse, FpAlu_8U_23U_and_30_cse, FpAlu_8U_23U_and_30_cse, FpAlu_8U_23U_and_30_cse, FpAlu_8U_23U_and_30_cse, FpAlu_8U_23U_and_30_cse, FpAlu_8U_23U_and_30_cse, FpAlu_8U_23U_and_30_cse, FpAlu_8U_23U_and_30_cse, FpAlu_8U_23U_and_30_cse, FpAlu_8U_23U_and_30_cse, FpAlu_8U_23U_and_30_cse, FpAlu_8U_23U_and_30_cse, FpAlu_8U_23U_and_30_cse, FpAlu_8U_23U_and_30_cse, FpAlu_8U_23U_and_30_cse };
  assign _1038_ = IntSaturation_33U_32U_slc_IntSaturation_33U_32U_o_31_1_3_21_0_itm_4 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16331" *) { asn_267, asn_267, asn_267, asn_267, asn_267, asn_267, asn_267, asn_267, asn_267, asn_267, asn_267, asn_267, asn_267, asn_267, asn_267, asn_267, asn_267, asn_267, asn_267, asn_267, asn_267, asn_267 };
  assign _1039_ = FpAlu_8U_23U_and_5_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16332" *) { nor_437_cse, nor_437_cse, nor_437_cse, nor_437_cse, nor_437_cse, nor_437_cse, nor_437_cse, nor_437_cse, nor_437_cse, nor_437_cse, nor_437_cse, nor_437_cse, nor_437_cse, nor_437_cse, nor_437_cse, nor_437_cse, nor_437_cse, nor_437_cse, nor_437_cse, nor_437_cse, nor_437_cse, nor_437_cse };
  assign _1040_ = FpAlu_8U_23U_and_8_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16332" *) { nor_437_cse, nor_437_cse, nor_437_cse, nor_437_cse, nor_437_cse, nor_437_cse, nor_437_cse, nor_437_cse, nor_437_cse, nor_437_cse, nor_437_cse, nor_437_cse, nor_437_cse, nor_437_cse, nor_437_cse, nor_437_cse, nor_437_cse, nor_437_cse, nor_437_cse, nor_437_cse, nor_437_cse, nor_437_cse };
  assign _1041_ = FpAlu_8U_23U_o_22_1_lpi_1_dfm_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16332" *) { nor_397_cse, nor_397_cse, nor_397_cse, nor_397_cse, nor_397_cse, nor_397_cse, nor_397_cse, nor_397_cse, nor_397_cse, nor_397_cse, nor_397_cse, nor_397_cse, nor_397_cse, nor_397_cse, nor_397_cse, nor_397_cse, nor_397_cse, nor_397_cse, nor_397_cse, nor_397_cse, nor_397_cse, nor_397_cse };
  assign _1042_ = FpCmp_8U_23U_true_o_3_lpi_1_dfm_7_30_0_1[22:1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16332" *) { FpAlu_8U_23U_equal_tmp_26, FpAlu_8U_23U_equal_tmp_26, FpAlu_8U_23U_equal_tmp_26, FpAlu_8U_23U_equal_tmp_26, FpAlu_8U_23U_equal_tmp_26, FpAlu_8U_23U_equal_tmp_26, FpAlu_8U_23U_equal_tmp_26, FpAlu_8U_23U_equal_tmp_26, FpAlu_8U_23U_equal_tmp_26, FpAlu_8U_23U_equal_tmp_26, FpAlu_8U_23U_equal_tmp_26, FpAlu_8U_23U_equal_tmp_26, FpAlu_8U_23U_equal_tmp_26, FpAlu_8U_23U_equal_tmp_26, FpAlu_8U_23U_equal_tmp_26, FpAlu_8U_23U_equal_tmp_26, FpAlu_8U_23U_equal_tmp_26, FpAlu_8U_23U_equal_tmp_26, FpAlu_8U_23U_equal_tmp_26, FpAlu_8U_23U_equal_tmp_26, FpAlu_8U_23U_equal_tmp_26, FpAlu_8U_23U_equal_tmp_26 };
  assign _1043_ = FpAlu_8U_23U_and_11_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16332" *) { nor_437_cse, nor_437_cse, nor_437_cse, nor_437_cse, nor_437_cse, nor_437_cse, nor_437_cse, nor_437_cse, nor_437_cse, nor_437_cse, nor_437_cse, nor_437_cse, nor_437_cse, nor_437_cse, nor_437_cse, nor_437_cse, nor_437_cse, nor_437_cse, nor_437_cse, nor_437_cse, nor_437_cse, nor_437_cse };
  assign _1044_ = FpCmp_8U_23U_false_o_lpi_1_dfm_9_30_0_1[22:1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16344" *) { FpAlu_8U_23U_and_45_cse, FpAlu_8U_23U_and_45_cse, FpAlu_8U_23U_and_45_cse, FpAlu_8U_23U_and_45_cse, FpAlu_8U_23U_and_45_cse, FpAlu_8U_23U_and_45_cse, FpAlu_8U_23U_and_45_cse, FpAlu_8U_23U_and_45_cse, FpAlu_8U_23U_and_45_cse, FpAlu_8U_23U_and_45_cse, FpAlu_8U_23U_and_45_cse, FpAlu_8U_23U_and_45_cse, FpAlu_8U_23U_and_45_cse, FpAlu_8U_23U_and_45_cse, FpAlu_8U_23U_and_45_cse, FpAlu_8U_23U_and_45_cse, FpAlu_8U_23U_and_45_cse, FpAlu_8U_23U_and_45_cse, FpAlu_8U_23U_and_45_cse, FpAlu_8U_23U_and_45_cse, FpAlu_8U_23U_and_45_cse, FpAlu_8U_23U_and_45_cse };
  assign _1045_ = FpAlu_8U_23U_o_22_1_lpi_1_dfm_4 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16345" *) { FpAlu_8U_23U_and_44_cse, FpAlu_8U_23U_and_44_cse, FpAlu_8U_23U_and_44_cse, FpAlu_8U_23U_and_44_cse, FpAlu_8U_23U_and_44_cse, FpAlu_8U_23U_and_44_cse, FpAlu_8U_23U_and_44_cse, FpAlu_8U_23U_and_44_cse, FpAlu_8U_23U_and_44_cse, FpAlu_8U_23U_and_44_cse, FpAlu_8U_23U_and_44_cse, FpAlu_8U_23U_and_44_cse, FpAlu_8U_23U_and_44_cse, FpAlu_8U_23U_and_44_cse, FpAlu_8U_23U_and_44_cse, FpAlu_8U_23U_and_44_cse, FpAlu_8U_23U_and_44_cse, FpAlu_8U_23U_and_44_cse, FpAlu_8U_23U_and_44_cse, FpAlu_8U_23U_and_44_cse, FpAlu_8U_23U_and_44_cse, FpAlu_8U_23U_and_44_cse };
  assign _1046_ = FpCmp_8U_23U_true_o_lpi_1_dfm_7_30_0_1[22:1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16346" *) { FpAlu_8U_23U_equal_tmp_26, FpAlu_8U_23U_equal_tmp_26, FpAlu_8U_23U_equal_tmp_26, FpAlu_8U_23U_equal_tmp_26, FpAlu_8U_23U_equal_tmp_26, FpAlu_8U_23U_equal_tmp_26, FpAlu_8U_23U_equal_tmp_26, FpAlu_8U_23U_equal_tmp_26, FpAlu_8U_23U_equal_tmp_26, FpAlu_8U_23U_equal_tmp_26, FpAlu_8U_23U_equal_tmp_26, FpAlu_8U_23U_equal_tmp_26, FpAlu_8U_23U_equal_tmp_26, FpAlu_8U_23U_equal_tmp_26, FpAlu_8U_23U_equal_tmp_26, FpAlu_8U_23U_equal_tmp_26, FpAlu_8U_23U_equal_tmp_26, FpAlu_8U_23U_equal_tmp_26, FpAlu_8U_23U_equal_tmp_26, FpAlu_8U_23U_equal_tmp_26, FpAlu_8U_23U_equal_tmp_26, FpAlu_8U_23U_equal_tmp_26 };
  assign _1047_ = reg_AluIn_data_sva_4_126_96_1_itm[22:1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16347" *) { FpAlu_8U_23U_nor_dfs_6, FpAlu_8U_23U_nor_dfs_6, FpAlu_8U_23U_nor_dfs_6, FpAlu_8U_23U_nor_dfs_6, FpAlu_8U_23U_nor_dfs_6, FpAlu_8U_23U_nor_dfs_6, FpAlu_8U_23U_nor_dfs_6, FpAlu_8U_23U_nor_dfs_6, FpAlu_8U_23U_nor_dfs_6, FpAlu_8U_23U_nor_dfs_6, FpAlu_8U_23U_nor_dfs_6, FpAlu_8U_23U_nor_dfs_6, FpAlu_8U_23U_nor_dfs_6, FpAlu_8U_23U_nor_dfs_6, FpAlu_8U_23U_nor_dfs_6, FpAlu_8U_23U_nor_dfs_6, FpAlu_8U_23U_nor_dfs_6, FpAlu_8U_23U_nor_dfs_6, FpAlu_8U_23U_nor_dfs_6, FpAlu_8U_23U_nor_dfs_6, FpAlu_8U_23U_nor_dfs_6, FpAlu_8U_23U_nor_dfs_6 };
  assign _1048_ = 30'b111111111111111111111111111111 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16358" *) { alu_loop_op_2_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_1_svs_3, alu_loop_op_2_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_1_svs_3, alu_loop_op_2_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_1_svs_3, alu_loop_op_2_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_1_svs_3, alu_loop_op_2_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_1_svs_3, alu_loop_op_2_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_1_svs_3, alu_loop_op_2_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_1_svs_3, alu_loop_op_2_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_1_svs_3, alu_loop_op_2_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_1_svs_3, alu_loop_op_2_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_1_svs_3, alu_loop_op_2_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_1_svs_3, alu_loop_op_2_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_1_svs_3, alu_loop_op_2_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_1_svs_3, alu_loop_op_2_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_1_svs_3, alu_loop_op_2_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_1_svs_3, alu_loop_op_2_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_1_svs_3, alu_loop_op_2_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_1_svs_3, alu_loop_op_2_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_1_svs_3, alu_loop_op_2_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_1_svs_3, alu_loop_op_2_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_1_svs_3, alu_loop_op_2_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_1_svs_3, alu_loop_op_2_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_1_svs_3, alu_loop_op_2_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_1_svs_3, alu_loop_op_2_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_1_svs_3, alu_loop_op_2_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_1_svs_3, alu_loop_op_2_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_1_svs_3, alu_loop_op_2_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_1_svs_3, alu_loop_op_2_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_1_svs_3, alu_loop_op_2_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_1_svs_3, alu_loop_op_2_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_1_svs_3, alu_loop_op_2_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_1_svs_3 };
  assign _1049_ = 30'b111111111111111111111111111111 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16358" *) { alu_loop_op_4_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_1_svs_2, alu_loop_op_4_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_1_svs_2, alu_loop_op_4_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_1_svs_2, alu_loop_op_4_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_1_svs_2, alu_loop_op_4_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_1_svs_2, alu_loop_op_4_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_1_svs_2, alu_loop_op_4_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_1_svs_2, alu_loop_op_4_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_1_svs_2, alu_loop_op_4_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_1_svs_2, alu_loop_op_4_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_1_svs_2, alu_loop_op_4_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_1_svs_2, alu_loop_op_4_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_1_svs_2, alu_loop_op_4_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_1_svs_2, alu_loop_op_4_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_1_svs_2, alu_loop_op_4_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_1_svs_2, alu_loop_op_4_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_1_svs_2, alu_loop_op_4_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_1_svs_2, alu_loop_op_4_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_1_svs_2, alu_loop_op_4_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_1_svs_2, alu_loop_op_4_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_1_svs_2, alu_loop_op_4_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_1_svs_2, alu_loop_op_4_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_1_svs_2, alu_loop_op_4_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_1_svs_2, alu_loop_op_4_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_1_svs_2, alu_loop_op_4_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_1_svs_2, alu_loop_op_4_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_1_svs_2, alu_loop_op_4_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_1_svs_2, alu_loop_op_4_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_1_svs_2, alu_loop_op_4_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_1_svs_2, alu_loop_op_4_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_1_svs_2, alu_loop_op_4_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_1_svs_2 };
  assign _1050_ = 30'b111111111111111111111111111111 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16358" *) { alu_loop_op_3_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_svs_2, alu_loop_op_3_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_svs_2, alu_loop_op_3_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_svs_2, alu_loop_op_3_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_svs_2, alu_loop_op_3_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_svs_2, alu_loop_op_3_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_svs_2, alu_loop_op_3_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_svs_2, alu_loop_op_3_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_svs_2, alu_loop_op_3_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_svs_2, alu_loop_op_3_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_svs_2, alu_loop_op_3_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_svs_2, alu_loop_op_3_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_svs_2, alu_loop_op_3_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_svs_2, alu_loop_op_3_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_svs_2, alu_loop_op_3_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_svs_2, alu_loop_op_3_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_svs_2, alu_loop_op_3_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_svs_2, alu_loop_op_3_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_svs_2, alu_loop_op_3_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_svs_2, alu_loop_op_3_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_svs_2, alu_loop_op_3_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_svs_2, alu_loop_op_3_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_svs_2, alu_loop_op_3_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_svs_2, alu_loop_op_3_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_svs_2, alu_loop_op_3_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_svs_2, alu_loop_op_3_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_svs_2, alu_loop_op_3_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_svs_2, alu_loop_op_3_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_svs_2, alu_loop_op_3_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_svs_2, alu_loop_op_3_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_svs_2, alu_loop_op_3_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_svs_2 };
  assign _1051_ = 30'b111111111111111111111111111111 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16358" *) { alu_loop_op_1_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_svs_2, alu_loop_op_1_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_svs_2, alu_loop_op_1_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_svs_2, alu_loop_op_1_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_svs_2, alu_loop_op_1_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_svs_2, alu_loop_op_1_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_svs_2, alu_loop_op_1_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_svs_2, alu_loop_op_1_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_svs_2, alu_loop_op_1_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_svs_2, alu_loop_op_1_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_svs_2, alu_loop_op_1_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_svs_2, alu_loop_op_1_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_svs_2, alu_loop_op_1_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_svs_2, alu_loop_op_1_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_svs_2, alu_loop_op_1_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_svs_2, alu_loop_op_1_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_svs_2, alu_loop_op_1_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_svs_2, alu_loop_op_1_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_svs_2, alu_loop_op_1_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_svs_2, alu_loop_op_1_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_svs_2, alu_loop_op_1_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_svs_2, alu_loop_op_1_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_svs_2, alu_loop_op_1_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_svs_2, alu_loop_op_1_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_svs_2, alu_loop_op_1_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_svs_2, alu_loop_op_1_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_svs_2, alu_loop_op_1_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_svs_2, alu_loop_op_1_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_svs_2, alu_loop_op_1_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_svs_2, alu_loop_op_1_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_svs_2, alu_loop_op_1_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_svs_2 };
  assign _1052_ = 31'b1000000000000000000000000000000 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16359" *) { IntSaturation_33U_32U_and_3_nl, IntSaturation_33U_32U_and_3_nl, IntSaturation_33U_32U_and_3_nl, IntSaturation_33U_32U_and_3_nl, IntSaturation_33U_32U_and_3_nl, IntSaturation_33U_32U_and_3_nl, IntSaturation_33U_32U_and_3_nl, IntSaturation_33U_32U_and_3_nl, IntSaturation_33U_32U_and_3_nl, IntSaturation_33U_32U_and_3_nl, IntSaturation_33U_32U_and_3_nl, IntSaturation_33U_32U_and_3_nl, IntSaturation_33U_32U_and_3_nl, IntSaturation_33U_32U_and_3_nl, IntSaturation_33U_32U_and_3_nl, IntSaturation_33U_32U_and_3_nl, IntSaturation_33U_32U_and_3_nl, IntSaturation_33U_32U_and_3_nl, IntSaturation_33U_32U_and_3_nl, IntSaturation_33U_32U_and_3_nl, IntSaturation_33U_32U_and_3_nl, IntSaturation_33U_32U_and_3_nl, IntSaturation_33U_32U_and_3_nl, IntSaturation_33U_32U_and_3_nl, IntSaturation_33U_32U_and_3_nl, IntSaturation_33U_32U_and_3_nl, IntSaturation_33U_32U_and_3_nl, IntSaturation_33U_32U_and_3_nl, IntSaturation_33U_32U_and_3_nl, IntSaturation_33U_32U_and_3_nl, IntSaturation_33U_32U_and_3_nl };
  assign _1053_ = 31'b1000000000000000000000000000000 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16359" *) { IntSaturation_33U_32U_and_7_nl, IntSaturation_33U_32U_and_7_nl, IntSaturation_33U_32U_and_7_nl, IntSaturation_33U_32U_and_7_nl, IntSaturation_33U_32U_and_7_nl, IntSaturation_33U_32U_and_7_nl, IntSaturation_33U_32U_and_7_nl, IntSaturation_33U_32U_and_7_nl, IntSaturation_33U_32U_and_7_nl, IntSaturation_33U_32U_and_7_nl, IntSaturation_33U_32U_and_7_nl, IntSaturation_33U_32U_and_7_nl, IntSaturation_33U_32U_and_7_nl, IntSaturation_33U_32U_and_7_nl, IntSaturation_33U_32U_and_7_nl, IntSaturation_33U_32U_and_7_nl, IntSaturation_33U_32U_and_7_nl, IntSaturation_33U_32U_and_7_nl, IntSaturation_33U_32U_and_7_nl, IntSaturation_33U_32U_and_7_nl, IntSaturation_33U_32U_and_7_nl, IntSaturation_33U_32U_and_7_nl, IntSaturation_33U_32U_and_7_nl, IntSaturation_33U_32U_and_7_nl, IntSaturation_33U_32U_and_7_nl, IntSaturation_33U_32U_and_7_nl, IntSaturation_33U_32U_and_7_nl, IntSaturation_33U_32U_and_7_nl, IntSaturation_33U_32U_and_7_nl, IntSaturation_33U_32U_and_7_nl, IntSaturation_33U_32U_and_7_nl };
  assign _1054_ = 31'b1000000000000000000000000000000 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16359" *) { IntSaturation_33U_32U_and_5_nl, IntSaturation_33U_32U_and_5_nl, IntSaturation_33U_32U_and_5_nl, IntSaturation_33U_32U_and_5_nl, IntSaturation_33U_32U_and_5_nl, IntSaturation_33U_32U_and_5_nl, IntSaturation_33U_32U_and_5_nl, IntSaturation_33U_32U_and_5_nl, IntSaturation_33U_32U_and_5_nl, IntSaturation_33U_32U_and_5_nl, IntSaturation_33U_32U_and_5_nl, IntSaturation_33U_32U_and_5_nl, IntSaturation_33U_32U_and_5_nl, IntSaturation_33U_32U_and_5_nl, IntSaturation_33U_32U_and_5_nl, IntSaturation_33U_32U_and_5_nl, IntSaturation_33U_32U_and_5_nl, IntSaturation_33U_32U_and_5_nl, IntSaturation_33U_32U_and_5_nl, IntSaturation_33U_32U_and_5_nl, IntSaturation_33U_32U_and_5_nl, IntSaturation_33U_32U_and_5_nl, IntSaturation_33U_32U_and_5_nl, IntSaturation_33U_32U_and_5_nl, IntSaturation_33U_32U_and_5_nl, IntSaturation_33U_32U_and_5_nl, IntSaturation_33U_32U_and_5_nl, IntSaturation_33U_32U_and_5_nl, IntSaturation_33U_32U_and_5_nl, IntSaturation_33U_32U_and_5_nl, IntSaturation_33U_32U_and_5_nl };
  assign _1055_ = 31'b1000000000000000000000000000000 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16359" *) { IntSaturation_33U_32U_and_1_nl, IntSaturation_33U_32U_and_1_nl, IntSaturation_33U_32U_and_1_nl, IntSaturation_33U_32U_and_1_nl, IntSaturation_33U_32U_and_1_nl, IntSaturation_33U_32U_and_1_nl, IntSaturation_33U_32U_and_1_nl, IntSaturation_33U_32U_and_1_nl, IntSaturation_33U_32U_and_1_nl, IntSaturation_33U_32U_and_1_nl, IntSaturation_33U_32U_and_1_nl, IntSaturation_33U_32U_and_1_nl, IntSaturation_33U_32U_and_1_nl, IntSaturation_33U_32U_and_1_nl, IntSaturation_33U_32U_and_1_nl, IntSaturation_33U_32U_and_1_nl, IntSaturation_33U_32U_and_1_nl, IntSaturation_33U_32U_and_1_nl, IntSaturation_33U_32U_and_1_nl, IntSaturation_33U_32U_and_1_nl, IntSaturation_33U_32U_and_1_nl, IntSaturation_33U_32U_and_1_nl, IntSaturation_33U_32U_and_1_nl, IntSaturation_33U_32U_and_1_nl, IntSaturation_33U_32U_and_1_nl, IntSaturation_33U_32U_and_1_nl, IntSaturation_33U_32U_and_1_nl, IntSaturation_33U_32U_and_1_nl, IntSaturation_33U_32U_and_1_nl, IntSaturation_33U_32U_and_1_nl, IntSaturation_33U_32U_and_1_nl };
  assign _1056_ = reg_alu_loop_op_else_o_32_1_2_lpi_1_dfm_4_1_itm & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16360" *) { IntSaturation_33U_32U_IntSaturation_33U_32U_nor_1_nl, IntSaturation_33U_32U_IntSaturation_33U_32U_nor_1_nl, IntSaturation_33U_32U_IntSaturation_33U_32U_nor_1_nl, IntSaturation_33U_32U_IntSaturation_33U_32U_nor_1_nl, IntSaturation_33U_32U_IntSaturation_33U_32U_nor_1_nl, IntSaturation_33U_32U_IntSaturation_33U_32U_nor_1_nl, IntSaturation_33U_32U_IntSaturation_33U_32U_nor_1_nl, IntSaturation_33U_32U_IntSaturation_33U_32U_nor_1_nl, IntSaturation_33U_32U_IntSaturation_33U_32U_nor_1_nl, IntSaturation_33U_32U_IntSaturation_33U_32U_nor_1_nl, IntSaturation_33U_32U_IntSaturation_33U_32U_nor_1_nl, IntSaturation_33U_32U_IntSaturation_33U_32U_nor_1_nl, IntSaturation_33U_32U_IntSaturation_33U_32U_nor_1_nl, IntSaturation_33U_32U_IntSaturation_33U_32U_nor_1_nl, IntSaturation_33U_32U_IntSaturation_33U_32U_nor_1_nl, IntSaturation_33U_32U_IntSaturation_33U_32U_nor_1_nl, IntSaturation_33U_32U_IntSaturation_33U_32U_nor_1_nl, IntSaturation_33U_32U_IntSaturation_33U_32U_nor_1_nl, IntSaturation_33U_32U_IntSaturation_33U_32U_nor_1_nl, IntSaturation_33U_32U_IntSaturation_33U_32U_nor_1_nl, IntSaturation_33U_32U_IntSaturation_33U_32U_nor_1_nl, IntSaturation_33U_32U_IntSaturation_33U_32U_nor_1_nl, IntSaturation_33U_32U_IntSaturation_33U_32U_nor_1_nl, IntSaturation_33U_32U_IntSaturation_33U_32U_nor_1_nl, IntSaturation_33U_32U_IntSaturation_33U_32U_nor_1_nl, IntSaturation_33U_32U_IntSaturation_33U_32U_nor_1_nl, IntSaturation_33U_32U_IntSaturation_33U_32U_nor_1_nl, IntSaturation_33U_32U_IntSaturation_33U_32U_nor_1_nl, IntSaturation_33U_32U_IntSaturation_33U_32U_nor_1_nl, IntSaturation_33U_32U_IntSaturation_33U_32U_nor_1_nl, IntSaturation_33U_32U_IntSaturation_33U_32U_nor_1_nl };
  assign _1057_ = reg_alu_loop_op_else_o_32_1_lpi_1_dfm_4_1_itm & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16360" *) { IntSaturation_33U_32U_IntSaturation_33U_32U_nor_3_nl, IntSaturation_33U_32U_IntSaturation_33U_32U_nor_3_nl, IntSaturation_33U_32U_IntSaturation_33U_32U_nor_3_nl, IntSaturation_33U_32U_IntSaturation_33U_32U_nor_3_nl, IntSaturation_33U_32U_IntSaturation_33U_32U_nor_3_nl, IntSaturation_33U_32U_IntSaturation_33U_32U_nor_3_nl, IntSaturation_33U_32U_IntSaturation_33U_32U_nor_3_nl, IntSaturation_33U_32U_IntSaturation_33U_32U_nor_3_nl, IntSaturation_33U_32U_IntSaturation_33U_32U_nor_3_nl, IntSaturation_33U_32U_IntSaturation_33U_32U_nor_3_nl, IntSaturation_33U_32U_IntSaturation_33U_32U_nor_3_nl, IntSaturation_33U_32U_IntSaturation_33U_32U_nor_3_nl, IntSaturation_33U_32U_IntSaturation_33U_32U_nor_3_nl, IntSaturation_33U_32U_IntSaturation_33U_32U_nor_3_nl, IntSaturation_33U_32U_IntSaturation_33U_32U_nor_3_nl, IntSaturation_33U_32U_IntSaturation_33U_32U_nor_3_nl, IntSaturation_33U_32U_IntSaturation_33U_32U_nor_3_nl, IntSaturation_33U_32U_IntSaturation_33U_32U_nor_3_nl, IntSaturation_33U_32U_IntSaturation_33U_32U_nor_3_nl, IntSaturation_33U_32U_IntSaturation_33U_32U_nor_3_nl, IntSaturation_33U_32U_IntSaturation_33U_32U_nor_3_nl, IntSaturation_33U_32U_IntSaturation_33U_32U_nor_3_nl, IntSaturation_33U_32U_IntSaturation_33U_32U_nor_3_nl, IntSaturation_33U_32U_IntSaturation_33U_32U_nor_3_nl, IntSaturation_33U_32U_IntSaturation_33U_32U_nor_3_nl, IntSaturation_33U_32U_IntSaturation_33U_32U_nor_3_nl, IntSaturation_33U_32U_IntSaturation_33U_32U_nor_3_nl, IntSaturation_33U_32U_IntSaturation_33U_32U_nor_3_nl, IntSaturation_33U_32U_IntSaturation_33U_32U_nor_3_nl, IntSaturation_33U_32U_IntSaturation_33U_32U_nor_3_nl, IntSaturation_33U_32U_IntSaturation_33U_32U_nor_3_nl };
  assign _1058_ = reg_alu_loop_op_else_o_32_1_3_lpi_1_dfm_3_1_itm & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16360" *) { IntSaturation_33U_32U_IntSaturation_33U_32U_nor_2_nl, IntSaturation_33U_32U_IntSaturation_33U_32U_nor_2_nl, IntSaturation_33U_32U_IntSaturation_33U_32U_nor_2_nl, IntSaturation_33U_32U_IntSaturation_33U_32U_nor_2_nl, IntSaturation_33U_32U_IntSaturation_33U_32U_nor_2_nl, IntSaturation_33U_32U_IntSaturation_33U_32U_nor_2_nl, IntSaturation_33U_32U_IntSaturation_33U_32U_nor_2_nl, IntSaturation_33U_32U_IntSaturation_33U_32U_nor_2_nl, IntSaturation_33U_32U_IntSaturation_33U_32U_nor_2_nl, IntSaturation_33U_32U_IntSaturation_33U_32U_nor_2_nl, IntSaturation_33U_32U_IntSaturation_33U_32U_nor_2_nl, IntSaturation_33U_32U_IntSaturation_33U_32U_nor_2_nl, IntSaturation_33U_32U_IntSaturation_33U_32U_nor_2_nl, IntSaturation_33U_32U_IntSaturation_33U_32U_nor_2_nl, IntSaturation_33U_32U_IntSaturation_33U_32U_nor_2_nl, IntSaturation_33U_32U_IntSaturation_33U_32U_nor_2_nl, IntSaturation_33U_32U_IntSaturation_33U_32U_nor_2_nl, IntSaturation_33U_32U_IntSaturation_33U_32U_nor_2_nl, IntSaturation_33U_32U_IntSaturation_33U_32U_nor_2_nl, IntSaturation_33U_32U_IntSaturation_33U_32U_nor_2_nl, IntSaturation_33U_32U_IntSaturation_33U_32U_nor_2_nl, IntSaturation_33U_32U_IntSaturation_33U_32U_nor_2_nl, IntSaturation_33U_32U_IntSaturation_33U_32U_nor_2_nl, IntSaturation_33U_32U_IntSaturation_33U_32U_nor_2_nl, IntSaturation_33U_32U_IntSaturation_33U_32U_nor_2_nl, IntSaturation_33U_32U_IntSaturation_33U_32U_nor_2_nl, IntSaturation_33U_32U_IntSaturation_33U_32U_nor_2_nl, IntSaturation_33U_32U_IntSaturation_33U_32U_nor_2_nl, IntSaturation_33U_32U_IntSaturation_33U_32U_nor_2_nl, IntSaturation_33U_32U_IntSaturation_33U_32U_nor_2_nl, IntSaturation_33U_32U_IntSaturation_33U_32U_nor_2_nl };
  assign { _1135_[30:7], _1059_ } = reg_alu_loop_op_else_o_32_1_1_lpi_1_dfm_3_1_itm & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16360" *) { IntSaturation_33U_32U_IntSaturation_33U_32U_nor_nl, IntSaturation_33U_32U_IntSaturation_33U_32U_nor_nl, IntSaturation_33U_32U_IntSaturation_33U_32U_nor_nl, IntSaturation_33U_32U_IntSaturation_33U_32U_nor_nl, IntSaturation_33U_32U_IntSaturation_33U_32U_nor_nl, IntSaturation_33U_32U_IntSaturation_33U_32U_nor_nl, IntSaturation_33U_32U_IntSaturation_33U_32U_nor_nl, IntSaturation_33U_32U_IntSaturation_33U_32U_nor_nl, IntSaturation_33U_32U_IntSaturation_33U_32U_nor_nl, IntSaturation_33U_32U_IntSaturation_33U_32U_nor_nl, IntSaturation_33U_32U_IntSaturation_33U_32U_nor_nl, IntSaturation_33U_32U_IntSaturation_33U_32U_nor_nl, IntSaturation_33U_32U_IntSaturation_33U_32U_nor_nl, IntSaturation_33U_32U_IntSaturation_33U_32U_nor_nl, IntSaturation_33U_32U_IntSaturation_33U_32U_nor_nl, IntSaturation_33U_32U_IntSaturation_33U_32U_nor_nl, IntSaturation_33U_32U_IntSaturation_33U_32U_nor_nl, IntSaturation_33U_32U_IntSaturation_33U_32U_nor_nl, IntSaturation_33U_32U_IntSaturation_33U_32U_nor_nl, IntSaturation_33U_32U_IntSaturation_33U_32U_nor_nl, IntSaturation_33U_32U_IntSaturation_33U_32U_nor_nl, IntSaturation_33U_32U_IntSaturation_33U_32U_nor_nl, IntSaturation_33U_32U_IntSaturation_33U_32U_nor_nl, IntSaturation_33U_32U_IntSaturation_33U_32U_nor_nl, IntSaturation_33U_32U_IntSaturation_33U_32U_nor_nl, IntSaturation_33U_32U_IntSaturation_33U_32U_nor_nl, IntSaturation_33U_32U_IntSaturation_33U_32U_nor_nl, IntSaturation_33U_32U_IntSaturation_33U_32U_nor_nl, IntSaturation_33U_32U_IntSaturation_33U_32U_nor_nl, IntSaturation_33U_32U_IntSaturation_33U_32U_nor_nl, IntSaturation_33U_32U_IntSaturation_33U_32U_nor_nl };
  assign _1060_ = reg_AluIn_data_sva_4_30_0_itm & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16371" *) { or_996_tmp, or_996_tmp, or_996_tmp, or_996_tmp, or_996_tmp, or_996_tmp, or_996_tmp, or_996_tmp };
  assign _1061_ = reg_AluIn_data_sva_4_62_32_itm & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16371" *) { or_997_tmp, or_997_tmp, or_997_tmp, or_997_tmp, or_997_tmp, or_997_tmp, or_997_tmp, or_997_tmp };
  assign _1062_ = reg_AluIn_data_sva_4_126_96_itm & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16371" *) { io_read_cfg_alu_bypass_rsc_svs_8, io_read_cfg_alu_bypass_rsc_svs_8, io_read_cfg_alu_bypass_rsc_svs_8, io_read_cfg_alu_bypass_rsc_svs_8, io_read_cfg_alu_bypass_rsc_svs_8, io_read_cfg_alu_bypass_rsc_svs_8, io_read_cfg_alu_bypass_rsc_svs_8, io_read_cfg_alu_bypass_rsc_svs_8 };
  assign _1063_ = FpAdd_8U_23U_qr_2_lpi_1_dfm & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16371" *) { and_dcpl_99, and_dcpl_99, and_dcpl_99, and_dcpl_99, and_dcpl_99, and_dcpl_99, and_dcpl_99, and_dcpl_99 };
  assign _1064_ = FpAdd_8U_23U_qr_3_lpi_1_dfm & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16371" *) { and_dcpl_99, and_dcpl_99, and_dcpl_99, and_dcpl_99, and_dcpl_99, and_dcpl_99, and_dcpl_99, and_dcpl_99 };
  assign _1065_ = FpAdd_8U_23U_qr_4_lpi_1_dfm & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16371" *) { and_dcpl_99, and_dcpl_99, and_dcpl_99, and_dcpl_99, and_dcpl_99, and_dcpl_99, and_dcpl_99, and_dcpl_99 };
  assign _1066_ = FpAdd_8U_23U_qr_lpi_1_dfm & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16371" *) { and_dcpl_99, and_dcpl_99, and_dcpl_99, and_dcpl_99, and_dcpl_99, and_dcpl_99, and_dcpl_99, and_dcpl_99 };
  assign _1067_ = else_AluOp_data_slc_else_AluOp_data_2_30_23_21_itm & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16371" *) { and_dcpl_169, and_dcpl_169, and_dcpl_169, and_dcpl_169, and_dcpl_169, and_dcpl_169, and_dcpl_169, and_dcpl_169 };
  assign _1068_ = else_AluOp_data_slc_else_AluOp_data_3_30_23_35_itm & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16371" *) { and_dcpl_169, and_dcpl_169, and_dcpl_169, and_dcpl_169, and_dcpl_169, and_dcpl_169, and_dcpl_169, and_dcpl_169 };
  assign _1069_ = else_AluOp_data_slc_else_AluOp_data_1_30_23_21_itm & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16371" *) { and_dcpl_169, and_dcpl_169, and_dcpl_169, and_dcpl_169, and_dcpl_169, and_dcpl_169, and_dcpl_169, and_dcpl_169 };
  assign _1070_ = else_AluOp_data_slc_else_AluOp_data_0_30_23_7_itm & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16371" *) { and_dcpl_169, and_dcpl_169, and_dcpl_169, and_dcpl_169, and_dcpl_169, and_dcpl_169, and_dcpl_169, and_dcpl_169 };
  assign _1071_ = reg_AluIn_data_sva_4_94_64_itm & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16371" *) { or_998_tmp, or_998_tmp, or_998_tmp, or_998_tmp, or_998_tmp, or_998_tmp, or_998_tmp, or_998_tmp };
  assign _1072_ = acc_nl[8:1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16371" *) { mux_tmp, mux_tmp, mux_tmp, mux_tmp, mux_tmp, mux_tmp, mux_tmp, mux_tmp };
  assign _1073_ = acc_1_nl[8:1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16371" *) { mux_tmp_348, mux_tmp_348, mux_tmp_348, mux_tmp_348, mux_tmp_348, mux_tmp_348, mux_tmp_348, mux_tmp_348 };
  assign _1074_ = acc_2_nl[8:1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16371" *) { mux_tmp_349, mux_tmp_349, mux_tmp_349, mux_tmp_349, mux_tmp_349, mux_tmp_349, mux_tmp_349, mux_tmp_349 };
  assign _1075_ = acc_3_nl[8:1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16371" *) { mux_tmp_350, mux_tmp_350, mux_tmp_350, mux_tmp_350, mux_tmp_350, mux_tmp_350, mux_tmp_350, mux_tmp_350 };
  assign _1076_ = AluOut_data_2_30_23_lpi_1_dfm_3 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16372" *) { asn_267, asn_267, asn_267, asn_267, asn_267, asn_267, asn_267, asn_267 };
  assign _1077_ = FpAdd_8U_23U_o_expo_1_lpi_1_dfm_13 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16372" *) { asn_267, asn_267, asn_267, asn_267, asn_267, asn_267, asn_267, asn_267 };
  assign _1078_ = FpAdd_8U_23U_o_expo_3_lpi_1_dfm_13 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16372" *) { asn_267, asn_267, asn_267, asn_267, asn_267, asn_267, asn_267, asn_267 };
  assign _1079_ = else_AluOp_data_0_lpi_1_dfm_mx1_tmp_30_23 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16372" *) { and_233_rgt, and_233_rgt, and_233_rgt, and_233_rgt, and_233_rgt, and_233_rgt, and_233_rgt, and_233_rgt };
  assign _1080_ = else_AluOp_data_1_lpi_1_dfm_mx1_tmp_30_23 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16372" *) { and_237_rgt, and_237_rgt, and_237_rgt, and_237_rgt, and_237_rgt, and_237_rgt, and_237_rgt, and_237_rgt };
  assign _1081_ = else_AluOp_data_2_lpi_1_dfm_mx1_tmp_30_23 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16372" *) { and_241_rgt, and_241_rgt, and_241_rgt, and_241_rgt, and_241_rgt, and_241_rgt, and_241_rgt, and_241_rgt };
  assign _1082_ = else_AluOp_data_3_lpi_1_dfm_mx1_tmp_30_23 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16372" *) { and_245_rgt, and_245_rgt, and_245_rgt, and_245_rgt, and_245_rgt, and_245_rgt, and_245_rgt, and_245_rgt };
  assign _1083_ = else_AluOp_data_2_lpi_1_dfm_2_30_0_1[30:23] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16372" *) { and_dcpl_168, and_dcpl_168, and_dcpl_168, and_dcpl_168, and_dcpl_168, and_dcpl_168, and_dcpl_168, and_dcpl_168 };
  assign _1084_ = else_AluOp_data_3_lpi_1_dfm_2_30_0_1[30:23] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16372" *) { and_dcpl_168, and_dcpl_168, and_dcpl_168, and_dcpl_168, and_dcpl_168, and_dcpl_168, and_dcpl_168, and_dcpl_168 };
  assign _1085_ = else_AluOp_data_1_lpi_1_dfm_2_30_0_1[30:23] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16372" *) { and_dcpl_168, and_dcpl_168, and_dcpl_168, and_dcpl_168, and_dcpl_168, and_dcpl_168, and_dcpl_168, and_dcpl_168 };
  assign _1086_ = else_AluOp_data_0_lpi_1_dfm_2_30_0_1[30:23] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16372" *) { and_dcpl_168, and_dcpl_168, and_dcpl_168, and_dcpl_168, and_dcpl_168, and_dcpl_168, and_dcpl_168, and_dcpl_168 };
  assign _1087_ = FpAdd_8U_23U_o_expo_2_lpi_1_dfm_13 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16372" *) { asn_267, asn_267, asn_267, asn_267, asn_267, asn_267, asn_267, asn_267 };
  assign _1088_ = FpAdd_8U_23U_qr_2_lpi_1_dfm_7 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16372" *) { FpAdd_8U_23U_and_4_tmp, FpAdd_8U_23U_and_4_tmp, FpAdd_8U_23U_and_4_tmp, FpAdd_8U_23U_and_4_tmp, FpAdd_8U_23U_and_4_tmp, FpAdd_8U_23U_and_4_tmp, FpAdd_8U_23U_and_4_tmp, FpAdd_8U_23U_and_4_tmp };
  assign _1089_ = FpAdd_8U_23U_qr_3_lpi_1_dfm_7 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16372" *) { FpAdd_8U_23U_and_10_tmp, FpAdd_8U_23U_and_10_tmp, FpAdd_8U_23U_and_10_tmp, FpAdd_8U_23U_and_10_tmp, FpAdd_8U_23U_and_10_tmp, FpAdd_8U_23U_and_10_tmp, FpAdd_8U_23U_and_10_tmp, FpAdd_8U_23U_and_10_tmp };
  assign _1090_ = FpAdd_8U_23U_qr_4_lpi_1_dfm_7 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16372" *) { FpAdd_8U_23U_and_16_tmp, FpAdd_8U_23U_and_16_tmp, FpAdd_8U_23U_and_16_tmp, FpAdd_8U_23U_and_16_tmp, FpAdd_8U_23U_and_16_tmp, FpAdd_8U_23U_and_16_tmp, FpAdd_8U_23U_and_16_tmp, FpAdd_8U_23U_and_16_tmp };
  assign _1091_ = FpAdd_8U_23U_qr_lpi_1_dfm_7 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16372" *) { FpAdd_8U_23U_and_22_tmp, FpAdd_8U_23U_and_22_tmp, FpAdd_8U_23U_and_22_tmp, FpAdd_8U_23U_and_22_tmp, FpAdd_8U_23U_and_22_tmp, FpAdd_8U_23U_and_22_tmp, FpAdd_8U_23U_and_22_tmp, FpAdd_8U_23U_and_22_tmp };
  assign _1092_ = FpAlu_8U_23U_and_4_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16373" *) { nor_406_nl, nor_406_nl, nor_406_nl, nor_406_nl, nor_406_nl, nor_406_nl, nor_406_nl, nor_406_nl };
  assign _1093_ = FpAlu_8U_23U_and_7_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16373" *) { nor_407_nl, nor_407_nl, nor_407_nl, nor_407_nl, nor_407_nl, nor_407_nl, nor_407_nl, nor_407_nl };
  assign _1094_ = FpAlu_8U_23U_o_30_23_lpi_1_dfm_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16373" *) { nor_397_cse, nor_397_cse, nor_397_cse, nor_397_cse, nor_397_cse, nor_397_cse, nor_397_cse, nor_397_cse };
  assign _1095_ = AluIn_data_sva_127[30:23] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16373" *) { and_231_rgt, and_231_rgt, and_231_rgt, and_231_rgt, and_231_rgt, and_231_rgt, and_231_rgt, and_231_rgt };
  assign _1096_ = AluIn_data_sva_127[62:55] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16373" *) { and_235_rgt, and_235_rgt, and_235_rgt, and_235_rgt, and_235_rgt, and_235_rgt, and_235_rgt, and_235_rgt };
  assign _1097_ = AluIn_data_sva_127[94:87] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16373" *) { and_239_rgt, and_239_rgt, and_239_rgt, and_239_rgt, and_239_rgt, and_239_rgt, and_239_rgt, and_239_rgt };
  assign _1098_ = AluIn_data_sva_127[126:119] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16373" *) { and_243_rgt, and_243_rgt, and_243_rgt, and_243_rgt, and_243_rgt, and_243_rgt, and_243_rgt, and_243_rgt };
  assign _1099_ = IntSaturation_33U_32U_o_31_1_3_lpi_1_dfm_1[29:22] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16373" *) { and_dcpl_165, and_dcpl_165, and_dcpl_165, and_dcpl_165, and_dcpl_165, and_dcpl_165, and_dcpl_165, and_dcpl_165 };
  assign _1100_ = IntSaturation_33U_32U_o_31_1_lpi_1_dfm_1[29:22] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16373" *) { and_dcpl_165, and_dcpl_165, and_dcpl_165, and_dcpl_165, and_dcpl_165, and_dcpl_165, and_dcpl_165, and_dcpl_165 };
  assign _1101_ = IntSaturation_33U_32U_o_31_1_2_lpi_1_dfm_1[29:22] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16373" *) { and_dcpl_165, and_dcpl_165, and_dcpl_165, and_dcpl_165, and_dcpl_165, and_dcpl_165, and_dcpl_165, and_dcpl_165 };
  assign _1102_ = IntSaturation_33U_32U_o_31_1_1_lpi_1_dfm_1[29:22] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16373" *) { and_dcpl_165, and_dcpl_165, and_dcpl_165, and_dcpl_165, and_dcpl_165, and_dcpl_165, and_dcpl_165, and_dcpl_165 };
  assign _1103_ = FpAlu_8U_23U_and_10_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16373" *) { nor_408_nl, nor_408_nl, nor_408_nl, nor_408_nl, nor_408_nl, nor_408_nl, nor_408_nl, nor_408_nl };
  assign _1104_ = { FpNormalize_8U_49U_oelse_not_9, FpNormalize_8U_49U_oelse_not_9, FpNormalize_8U_49U_oelse_not_9, FpNormalize_8U_49U_oelse_not_9, FpNormalize_8U_49U_oelse_not_9, FpNormalize_8U_49U_oelse_not_9, FpNormalize_8U_49U_oelse_not_9, FpNormalize_8U_49U_oelse_not_9 } & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16373" *) { nor_436_nl, nor_436_nl, nor_436_nl, nor_436_nl, nor_436_nl, nor_436_nl, nor_436_nl, nor_436_nl };
  assign _1105_ = { FpNormalize_8U_49U_oelse_not_11, FpNormalize_8U_49U_oelse_not_11, FpNormalize_8U_49U_oelse_not_11, FpNormalize_8U_49U_oelse_not_11, FpNormalize_8U_49U_oelse_not_11, FpNormalize_8U_49U_oelse_not_11, FpNormalize_8U_49U_oelse_not_11, FpNormalize_8U_49U_oelse_not_11 } & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16373" *) { nor_435_nl, nor_435_nl, nor_435_nl, nor_435_nl, nor_435_nl, nor_435_nl, nor_435_nl, nor_435_nl };
  assign _1106_ = { FpNormalize_8U_49U_oelse_not_13, FpNormalize_8U_49U_oelse_not_13, FpNormalize_8U_49U_oelse_not_13, FpNormalize_8U_49U_oelse_not_13, FpNormalize_8U_49U_oelse_not_13, FpNormalize_8U_49U_oelse_not_13, FpNormalize_8U_49U_oelse_not_13, FpNormalize_8U_49U_oelse_not_13 } & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16373" *) { nor_434_nl, nor_434_nl, nor_434_nl, nor_434_nl, nor_434_nl, nor_434_nl, nor_434_nl, nor_434_nl };
  assign _1107_ = { FpNormalize_8U_49U_oelse_not_15, FpNormalize_8U_49U_oelse_not_15, FpNormalize_8U_49U_oelse_not_15, FpNormalize_8U_49U_oelse_not_15, FpNormalize_8U_49U_oelse_not_15, FpNormalize_8U_49U_oelse_not_15, FpNormalize_8U_49U_oelse_not_15, FpNormalize_8U_49U_oelse_not_15 } & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16373" *) { nor_433_nl, nor_433_nl, nor_433_nl, nor_433_nl, nor_433_nl, nor_433_nl, nor_433_nl, nor_433_nl };
  assign _1108_ = FpCmp_8U_23U_false_o_1_lpi_1_dfm_7_30_0_1[30:23] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16387" *) { FpAlu_8U_23U_equal_tmp_29, FpAlu_8U_23U_equal_tmp_29, FpAlu_8U_23U_equal_tmp_29, FpAlu_8U_23U_equal_tmp_29, FpAlu_8U_23U_equal_tmp_29, FpAlu_8U_23U_equal_tmp_29, FpAlu_8U_23U_equal_tmp_29, FpAlu_8U_23U_equal_tmp_29 };
  assign _1109_ = FpCmp_8U_23U_false_o_2_lpi_1_dfm_8_30_0_1[30:23] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16387" *) { FpAlu_8U_23U_equal_tmp_29, FpAlu_8U_23U_equal_tmp_29, FpAlu_8U_23U_equal_tmp_29, FpAlu_8U_23U_equal_tmp_29, FpAlu_8U_23U_equal_tmp_29, FpAlu_8U_23U_equal_tmp_29, FpAlu_8U_23U_equal_tmp_29, FpAlu_8U_23U_equal_tmp_29 };
  assign _1110_ = FpCmp_8U_23U_true_o_1_lpi_1_dfm_7_30_0_1[30:23] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16388" *) { FpAlu_8U_23U_equal_tmp_26, FpAlu_8U_23U_equal_tmp_26, FpAlu_8U_23U_equal_tmp_26, FpAlu_8U_23U_equal_tmp_26, FpAlu_8U_23U_equal_tmp_26, FpAlu_8U_23U_equal_tmp_26, FpAlu_8U_23U_equal_tmp_26, FpAlu_8U_23U_equal_tmp_26 };
  assign _1111_ = FpCmp_8U_23U_true_o_2_lpi_1_dfm_7_30_0_1[30:23] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16388" *) { FpAlu_8U_23U_equal_tmp_26, FpAlu_8U_23U_equal_tmp_26, FpAlu_8U_23U_equal_tmp_26, FpAlu_8U_23U_equal_tmp_26, FpAlu_8U_23U_equal_tmp_26, FpAlu_8U_23U_equal_tmp_26, FpAlu_8U_23U_equal_tmp_26, FpAlu_8U_23U_equal_tmp_26 };
  assign _1112_ = else_AluOp_data_slc_else_AluOp_data_0_30_23_7_itm_3 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16389" *) { FpAdd_8U_23U_and_9_nl, FpAdd_8U_23U_and_9_nl, FpAdd_8U_23U_and_9_nl, FpAdd_8U_23U_and_9_nl, FpAdd_8U_23U_and_9_nl, FpAdd_8U_23U_and_9_nl, FpAdd_8U_23U_and_9_nl, FpAdd_8U_23U_and_9_nl };
  assign _1113_ = else_AluOp_data_slc_else_AluOp_data_1_30_23_21_itm_3 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16389" *) { FpAdd_8U_23U_and_15_nl, FpAdd_8U_23U_and_15_nl, FpAdd_8U_23U_and_15_nl, FpAdd_8U_23U_and_15_nl, FpAdd_8U_23U_and_15_nl, FpAdd_8U_23U_and_15_nl, FpAdd_8U_23U_and_15_nl, FpAdd_8U_23U_and_15_nl };
  assign _1114_ = 8'b11111110 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16390" *) { FpAdd_8U_23U_and_28_nl, FpAdd_8U_23U_and_28_nl, FpAdd_8U_23U_and_28_nl, FpAdd_8U_23U_and_28_nl, FpAdd_8U_23U_and_28_nl, FpAdd_8U_23U_and_28_nl, FpAdd_8U_23U_and_28_nl, FpAdd_8U_23U_and_28_nl };
  assign _1115_ = 8'b11111110 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16390" *) { FpAdd_8U_23U_and_30_nl, FpAdd_8U_23U_and_30_nl, FpAdd_8U_23U_and_30_nl, FpAdd_8U_23U_and_30_nl, FpAdd_8U_23U_and_30_nl, FpAdd_8U_23U_and_30_nl, FpAdd_8U_23U_and_30_nl, FpAdd_8U_23U_and_30_nl };
  assign _1116_ = alu_loop_op_1_FpAdd_8U_23U_if_4_if_acc_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16391" *) { FpAdd_8U_23U_and_6_nl, FpAdd_8U_23U_and_6_nl, FpAdd_8U_23U_and_6_nl, FpAdd_8U_23U_and_6_nl, FpAdd_8U_23U_and_6_nl, FpAdd_8U_23U_and_6_nl, FpAdd_8U_23U_and_6_nl, FpAdd_8U_23U_and_6_nl };
  assign _1117_ = alu_loop_op_2_FpAdd_8U_23U_if_4_if_acc_5_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16391" *) { FpAdd_8U_23U_and_13_nl, FpAdd_8U_23U_and_13_nl, FpAdd_8U_23U_and_13_nl, FpAdd_8U_23U_and_13_nl, FpAdd_8U_23U_and_13_nl, FpAdd_8U_23U_and_13_nl, FpAdd_8U_23U_and_13_nl, FpAdd_8U_23U_and_13_nl };
  assign _1118_ = FpAdd_8U_23U_o_expo_1_lpi_1_dfm_13 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16392" *) { FpAdd_8U_23U_and_nl, FpAdd_8U_23U_and_nl, FpAdd_8U_23U_and_nl, FpAdd_8U_23U_and_nl, FpAdd_8U_23U_and_nl, FpAdd_8U_23U_and_nl, FpAdd_8U_23U_and_nl, FpAdd_8U_23U_and_nl };
  assign _1119_ = FpAdd_8U_23U_o_expo_2_lpi_1_dfm_13 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16392" *) { FpAdd_8U_23U_and_29_nl, FpAdd_8U_23U_and_29_nl, FpAdd_8U_23U_and_29_nl, FpAdd_8U_23U_and_29_nl, FpAdd_8U_23U_and_29_nl, FpAdd_8U_23U_and_29_nl, FpAdd_8U_23U_and_29_nl, FpAdd_8U_23U_and_29_nl };
  assign _1120_ = FpCmp_8U_23U_false_o_3_lpi_1_dfm_8_30_0_1[30:23] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16407" *) { FpAlu_8U_23U_and_31_m1c, FpAlu_8U_23U_and_31_m1c, FpAlu_8U_23U_and_31_m1c, FpAlu_8U_23U_and_31_m1c, FpAlu_8U_23U_and_31_m1c, FpAlu_8U_23U_and_31_m1c, FpAlu_8U_23U_and_31_m1c, FpAlu_8U_23U_and_31_m1c };
  assign _1121_ = AluOut_data_2_30_23_lpi_1_dfm_3 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16408" *) { FpAlu_8U_23U_and_30_cse, FpAlu_8U_23U_and_30_cse, FpAlu_8U_23U_and_30_cse, FpAlu_8U_23U_and_30_cse, FpAlu_8U_23U_and_30_cse, FpAlu_8U_23U_and_30_cse, FpAlu_8U_23U_and_30_cse, FpAlu_8U_23U_and_30_cse };
  assign _1122_ = FpCmp_8U_23U_true_o_3_lpi_1_dfm_7_30_0_1[30:23] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16409" *) { FpAlu_8U_23U_equal_tmp_26, FpAlu_8U_23U_equal_tmp_26, FpAlu_8U_23U_equal_tmp_26, FpAlu_8U_23U_equal_tmp_26, FpAlu_8U_23U_equal_tmp_26, FpAlu_8U_23U_equal_tmp_26, FpAlu_8U_23U_equal_tmp_26, FpAlu_8U_23U_equal_tmp_26 };
  assign _1123_ = else_AluOp_data_slc_else_AluOp_data_2_30_23_21_itm_3 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16410" *) { FpAdd_8U_23U_and_21_nl, FpAdd_8U_23U_and_21_nl, FpAdd_8U_23U_and_21_nl, FpAdd_8U_23U_and_21_nl, FpAdd_8U_23U_and_21_nl, FpAdd_8U_23U_and_21_nl, FpAdd_8U_23U_and_21_nl, FpAdd_8U_23U_and_21_nl };
  assign _1124_ = 8'b11111110 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16411" *) { FpAdd_8U_23U_and_32_nl, FpAdd_8U_23U_and_32_nl, FpAdd_8U_23U_and_32_nl, FpAdd_8U_23U_and_32_nl, FpAdd_8U_23U_and_32_nl, FpAdd_8U_23U_and_32_nl, FpAdd_8U_23U_and_32_nl, FpAdd_8U_23U_and_32_nl };
  assign _1125_ = alu_loop_op_3_FpAdd_8U_23U_if_4_if_acc_3_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16412" *) { FpAdd_8U_23U_and_19_nl, FpAdd_8U_23U_and_19_nl, FpAdd_8U_23U_and_19_nl, FpAdd_8U_23U_and_19_nl, FpAdd_8U_23U_and_19_nl, FpAdd_8U_23U_and_19_nl, FpAdd_8U_23U_and_19_nl, FpAdd_8U_23U_and_19_nl };
  assign _1126_ = FpAdd_8U_23U_o_expo_3_lpi_1_dfm_13 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16413" *) { FpAdd_8U_23U_and_31_nl, FpAdd_8U_23U_and_31_nl, FpAdd_8U_23U_and_31_nl, FpAdd_8U_23U_and_31_nl, FpAdd_8U_23U_and_31_nl, FpAdd_8U_23U_and_31_nl, FpAdd_8U_23U_and_31_nl, FpAdd_8U_23U_and_31_nl };
  assign _1127_ = FpCmp_8U_23U_false_o_lpi_1_dfm_9_30_0_1[30:23] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16429" *) { FpAlu_8U_23U_and_45_cse, FpAlu_8U_23U_and_45_cse, FpAlu_8U_23U_and_45_cse, FpAlu_8U_23U_and_45_cse, FpAlu_8U_23U_and_45_cse, FpAlu_8U_23U_and_45_cse, FpAlu_8U_23U_and_45_cse, FpAlu_8U_23U_and_45_cse };
  assign _1128_ = FpAlu_8U_23U_o_30_23_lpi_1_dfm_4 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16430" *) { FpAlu_8U_23U_and_44_cse, FpAlu_8U_23U_and_44_cse, FpAlu_8U_23U_and_44_cse, FpAlu_8U_23U_and_44_cse, FpAlu_8U_23U_and_44_cse, FpAlu_8U_23U_and_44_cse, FpAlu_8U_23U_and_44_cse, FpAlu_8U_23U_and_44_cse };
  assign _1129_ = FpCmp_8U_23U_true_o_lpi_1_dfm_7_30_0_1[30:23] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16431" *) { FpAlu_8U_23U_equal_tmp_26, FpAlu_8U_23U_equal_tmp_26, FpAlu_8U_23U_equal_tmp_26, FpAlu_8U_23U_equal_tmp_26, FpAlu_8U_23U_equal_tmp_26, FpAlu_8U_23U_equal_tmp_26, FpAlu_8U_23U_equal_tmp_26, FpAlu_8U_23U_equal_tmp_26 };
  assign _1130_ = reg_AluIn_data_sva_4_126_96_itm & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16432" *) { FpAlu_8U_23U_and_62_nl, FpAlu_8U_23U_and_62_nl, FpAlu_8U_23U_and_62_nl, FpAlu_8U_23U_and_62_nl, FpAlu_8U_23U_and_62_nl, FpAlu_8U_23U_and_62_nl, FpAlu_8U_23U_and_62_nl, FpAlu_8U_23U_and_62_nl };
  assign _1131_ = else_AluOp_data_slc_else_AluOp_data_3_30_23_35_itm_3 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16433" *) { FpAdd_8U_23U_and_27_nl, FpAdd_8U_23U_and_27_nl, FpAdd_8U_23U_and_27_nl, FpAdd_8U_23U_and_27_nl, FpAdd_8U_23U_and_27_nl, FpAdd_8U_23U_and_27_nl, FpAdd_8U_23U_and_27_nl, FpAdd_8U_23U_and_27_nl };
  assign _1132_ = 8'b11111110 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16434" *) { FpAdd_8U_23U_and_34_nl, FpAdd_8U_23U_and_34_nl, FpAdd_8U_23U_and_34_nl, FpAdd_8U_23U_and_34_nl, FpAdd_8U_23U_and_34_nl, FpAdd_8U_23U_and_34_nl, FpAdd_8U_23U_and_34_nl, FpAdd_8U_23U_and_34_nl };
  assign _1133_ = alu_loop_op_4_FpAdd_8U_23U_if_4_if_acc_7_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16435" *) { FpAdd_8U_23U_and_25_nl, FpAdd_8U_23U_and_25_nl, FpAdd_8U_23U_and_25_nl, FpAdd_8U_23U_and_25_nl, FpAdd_8U_23U_and_25_nl, FpAdd_8U_23U_and_25_nl, FpAdd_8U_23U_and_25_nl, FpAdd_8U_23U_and_25_nl };
  assign _1134_ = FpAdd_8U_23U_o_expo_lpi_1_dfm_13 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16436" *) { FpAdd_8U_23U_and_33_nl, FpAdd_8U_23U_and_33_nl, FpAdd_8U_23U_and_33_nl, FpAdd_8U_23U_and_33_nl, FpAdd_8U_23U_and_33_nl, FpAdd_8U_23U_and_33_nl, FpAdd_8U_23U_and_33_nl, FpAdd_8U_23U_and_33_nl };
  assign and_564_cse = cfg_alu_algo_1_sva_st_24 == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12333" *) 2'b10;
  assign and_dcpl_77 = cfg_precision == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12509" *) 2'b10;
  assign FpAlu_8U_23U_equal_tmp_1_mx0w0 = cfg_alu_algo_1_sva_2 == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12530" *) 2'b11;
  assign and_451_cse = cfg_alu_algo_rsci_d == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12595" *) 2'b11;
  assign alu_loop_op_1_FpAdd_8U_23U_is_a_greater_oif_equal_tmp = AluIn_data_sva_127[30:23] == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12649" *) else_AluOp_data_0_lpi_1_dfm_mx1_tmp_30_23;
  assign alu_loop_op_2_FpAdd_8U_23U_is_a_greater_oif_equal_2_tmp = AluIn_data_sva_127[62:55] == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12651" *) else_AluOp_data_1_lpi_1_dfm_mx1_tmp_30_23;
  assign alu_loop_op_3_FpAdd_8U_23U_is_a_greater_oif_equal_1_tmp = AluIn_data_sva_127[94:87] == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12653" *) else_AluOp_data_2_lpi_1_dfm_mx1_tmp_30_23;
  assign alu_loop_op_4_FpAdd_8U_23U_is_a_greater_oif_equal_3_tmp = AluIn_data_sva_127[126:119] == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12655" *) else_AluOp_data_3_lpi_1_dfm_mx1_tmp_30_23;
  assign FpAlu_8U_23U_equal_tmp_2_mx0w0 = cfg_alu_algo_1_sva_2 == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12768" *) 1'b1;
  assign alu_loop_op_else_equal_tmp_2 = cfg_alu_algo_1_sva_2 == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12819" *) 2'b10;
  assign _1138_ = chn_alu_in_rsci_d_mxwt[126:119] == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12820" *) 8'b11111111;
  assign _1139_ = chn_alu_in_rsci_d_mxwt[94:87] == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12821" *) 8'b11111111;
  assign _1140_ = FpAdd_8U_23U_int_mant_1_lpi_1_dfm_2_mx0[48:25] == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12880" *) 24'b111111111111111111111111;
  assign _1141_ = FpAdd_8U_23U_int_mant_4_lpi_1_dfm_2_mx0[48:25] == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12900" *) 24'b111111111111111111111111;
  assign _1142_ = FpAdd_8U_23U_int_mant_3_lpi_1_dfm_2_mx0[48:25] == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12920" *) 24'b111111111111111111111111;
  assign _1143_ = FpAdd_8U_23U_int_mant_2_lpi_1_dfm_2_mx0[48:25] == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12940" *) 24'b111111111111111111111111;
  assign _1144_ = else_mux_1_tmp_31_23[7:0] == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13137" *) 8'b11111111;
  assign nor_tmp_126 = cfg_alu_algo_1_sva_st == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13441" *) 2'b11;
  assign _1145_ = ! (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13529" *) cfg_alu_algo_rsci_d;
  assign _1146_ = cfg_alu_algo_rsci_d == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13532" *) 2'b10;
  assign or_1050_cse = cfg_precision != (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12279" *) 2'b10;
  assign _1147_ = cfg_alu_algo_1_sva_st_20 != (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12281" *) 1'b1;
  assign _1148_ = cfg_alu_algo_1_sva_st_24 != (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12336" *) 2'b10;
  assign or_236_nl = cfg_alu_algo_1_sva_st_25 != (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12353" *) 2'b10;
  assign or_dcpl_86 = cfg_alu_algo_1_sva_st_23 != (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12465" *) 2'b10;
  assign _1149_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12546" *) cfg_alu_algo_1_sva_2;
  assign or_1055_cse = cfg_alu_algo_1_sva_2 != (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12556" *) 1'b1;
  assign alu_loop_op_4_FpAdd_8U_23U_IsZero_8U_23U_1_or_itm_mx0w0 = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12660" *) else_AluOp_data_3_lpi_1_dfm_mx0[30:0];
  assign _1150_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12670" *) else_AluOp_data_2_lpi_1_dfm_mx0[22:0];
  assign _1151_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12671" *) else_AluOp_data_2_lpi_1_dfm_mx3_30_0[30:23];
  assign _1152_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12681" *) else_AluOp_data_1_lpi_1_dfm_mx2_30_0[22:0];
  assign _1153_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12682" *) else_AluOp_data_1_lpi_1_dfm_mx0[30:23];
  assign _1154_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12692" *) else_AluOp_data_0_lpi_1_dfm_mx0[22:0];
  assign _1155_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12693" *) else_AluOp_data_0_lpi_1_dfm_mx3_30_0[30:23];
  assign FpNormalize_8U_49U_if_or_itm_mx0w0 = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12699" *) acc_12_nl[49:1];
  assign FpNormalize_8U_49U_if_or_1_itm_mx0w0 = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12700" *) acc_13_nl[49:1];
  assign FpNormalize_8U_49U_if_or_2_itm_mx0w0 = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12701" *) acc_14_nl[49:1];
  assign FpNormalize_8U_49U_if_or_3_itm_mx0w0 = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12702" *) acc_15_nl[49:1];
  assign alu_loop_op_4_FpAdd_8U_23U_IsZero_8U_23U_or_itm_mx0w0 = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12755" *) chn_alu_in_rsci_d_mxwt[126:96];
  assign alu_loop_op_3_FpAdd_8U_23U_IsZero_8U_23U_or_itm_mx0w0 = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12756" *) chn_alu_in_rsci_d_mxwt[94:64];
  assign alu_loop_op_2_FpAdd_8U_23U_IsZero_8U_23U_or_itm_mx0w0 = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12758" *) chn_alu_in_rsci_d_mxwt[62:32];
  assign _1156_ = else_AluOp_data_3_lpi_1_dfm_mx0[30:23] != (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12759" *) 8'b11111111;
  assign _1157_ = else_AluOp_data_2_lpi_1_dfm_mx3_30_0[30:23] != (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12760" *) 8'b11111111;
  assign _1158_ = else_AluOp_data_1_lpi_1_dfm_mx0[30:23] != (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12761" *) 8'b11111111;
  assign _1159_ = else_AluOp_data_0_lpi_1_dfm_mx3_30_0[30:23] != (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12762" *) 8'b11111111;
  assign FpAlu_8U_23U_o_0_sva_2_mx0w0 = AluIn_data_sva_127[127:96] != (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12763" *) else_AluOp_data_3_lpi_1_dfm_mx0;
  assign AluOut_data_2_0_sva_3_mx0w0 = AluIn_data_sva_127[95:64] != (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12764" *) else_AluOp_data_2_lpi_1_dfm_mx0;
  assign _1160_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12811" *) chn_alu_in_rsci_d_mxwt[22:0];
  assign _1161_ = chn_alu_in_rsci_d_mxwt[30:23] != (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12812" *) 8'b11111111;
  assign _1162_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12813" *) chn_alu_in_rsci_d_mxwt[54:32];
  assign _1163_ = chn_alu_in_rsci_d_mxwt[62:55] != (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12814" *) 8'b11111111;
  assign _1164_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12826" *) chn_alu_in_rsci_d_mxwt[118:96];
  assign _1165_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12827" *) chn_alu_in_rsci_d_mxwt[86:64];
  assign alu_loop_op_1_FpAdd_8U_23U_IsZero_8U_23U_or_itm_mx0w2 = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12828" *) chn_alu_in_rsci_d_mxwt[30:0];
  assign _1166_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13256" *) else_AluOp_data_3_lpi_1_dfm_mx0[22:0];
  assign _1167_ = cfg_alu_algo_1_sva_st_22 != (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13270" *) 1'b1;
  assign or_dcpl_154 = reg_cfg_alu_algo_1_sva_st_13_cse != (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13271" *) 1'b1;
  assign or_632_cse = cfg_alu_algo_1_sva_st_22 != (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13345" *) 2'b10;
  assign or_391_cse = cfg_alu_algo_1_sva_st != (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13357" *) 2'b10;
  assign or_381_cse = cfg_alu_algo_rsci_d != (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13358" *) 2'b10;
  assign or_tmp_382 = cfg_alu_algo_1_sva_st != (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13359" *) 1'b1;
  assign or_400_nl = cfg_alu_algo_rsci_d != (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13429" *) 1'b1;
  assign _1168_ = cfg_alu_algo_1_sva_st_28 != (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13436" *) 1'b1;
  assign _1169_ = else_mux_tmp_31_23[7:0] != (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13534" *) 8'b11111111;
  assign _1170_ = else_mux_2_tmp_31_23[7:0] != (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13535" *) 8'b11111111;
  assign _1171_ = else_mux_3_tmp_31_23[7:0] != (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13536" *) 8'b11111111;
  assign _1172_ = AluIn_data_sva_127[63:32] != (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15246" *) else_AluOp_data_1_lpi_1_dfm_mx0;
  assign _1173_ = AluIn_data_sva_127[31:0] != (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15249" *) else_AluOp_data_0_lpi_1_dfm_mx0;
  assign _1174_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11932" *) FpAdd_8U_23U_b_right_shift_qr_1_lpi_1_dfm_5[7:1];
  assign nl_alu_loop_op_1_FpAdd_8U_23U_b_int_mant_p1_lshift_rg_s[0] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11936" *) FpAdd_8U_23U_b_right_shift_qr_1_lpi_1_dfm_5[0];
  assign _1175_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11943" *) FpAdd_8U_23U_b_right_shift_qr_2_lpi_1_dfm_5[7:1];
  assign nl_alu_loop_op_2_FpAdd_8U_23U_b_int_mant_p1_lshift_2_rg_s[0] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11947" *) FpAdd_8U_23U_b_right_shift_qr_2_lpi_1_dfm_5[0];
  assign _1176_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11954" *) FpAdd_8U_23U_b_right_shift_qr_3_lpi_1_dfm_5[7:1];
  assign nl_alu_loop_op_3_FpAdd_8U_23U_b_int_mant_p1_lshift_1_rg_s[0] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11958" *) FpAdd_8U_23U_b_right_shift_qr_3_lpi_1_dfm_5[0];
  assign _1177_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11965" *) FpAdd_8U_23U_b_right_shift_qr_lpi_1_dfm_5[7:1];
  assign nl_alu_loop_op_4_FpAdd_8U_23U_b_int_mant_p1_lshift_3_rg_s[0] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11969" *) FpAdd_8U_23U_b_right_shift_qr_lpi_1_dfm_5[0];
  assign _1178_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11976" *) FpAdd_8U_23U_a_right_shift_qr_lpi_1_dfm_5[7:1];
  assign nl_alu_loop_op_4_FpAdd_8U_23U_a_int_mant_p1_lshift_3_rg_s[0] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11980" *) FpAdd_8U_23U_a_right_shift_qr_lpi_1_dfm_5[0];
  assign _1179_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11987" *) FpAdd_8U_23U_a_right_shift_qr_3_lpi_1_dfm_5[7:1];
  assign nl_alu_loop_op_3_FpAdd_8U_23U_a_int_mant_p1_lshift_1_rg_s[0] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11991" *) FpAdd_8U_23U_a_right_shift_qr_3_lpi_1_dfm_5[0];
  assign _1180_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:11998" *) FpAdd_8U_23U_a_right_shift_qr_2_lpi_1_dfm_5[7:1];
  assign nl_alu_loop_op_2_FpAdd_8U_23U_a_int_mant_p1_lshift_2_rg_s[0] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12002" *) FpAdd_8U_23U_a_right_shift_qr_2_lpi_1_dfm_5[0];
  assign _1181_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12009" *) FpAdd_8U_23U_a_right_shift_qr_1_lpi_1_dfm_5[7:1];
  assign nl_alu_loop_op_1_FpAdd_8U_23U_a_int_mant_p1_lshift_rg_s[0] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12013" *) FpAdd_8U_23U_a_right_shift_qr_1_lpi_1_dfm_5[0];
  assign _1182_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12267" *) or_dcpl_23;
  assign nor_437_cse = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12268" *) _1478_;
  assign _1183_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12269" *) reg_chn_alu_out_rsci_ld_core_psct_cse;
  assign _1184_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12273" *) fsm_output[0];
  assign _1185_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12275" *) and_dcpl_4;
  assign _1186_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12275" *) _1484_;
  assign nand_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12275" *) _0483_;
  assign _1187_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12278" *) or_dcpl_49;
  assign _1188_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12280" *) chn_alu_in_rsci_bawt;
  assign _1189_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12285" *) cfg_alu_src_1_sva_st_1;
  assign _1190_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12289" *) io_read_cfg_alu_bypass_rsc_svs_st_1;
  assign _1191_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12291" *) and_dcpl_32;
  assign _1192_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12296" *) main_stage_v_1;
  assign _1193_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12298" *) _0493_;
  assign nor_367_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12298" *) _1486_;
  assign _1194_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12299" *) main_stage_v_2;
  assign nor_368_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12299" *) _1487_;
  assign _1195_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12311" *) FpAdd_8U_23U_int_mant_p1_1_lpi_1_dfm_5[49];
  assign nor_33_cse = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12311" *) _1488_;
  assign _1196_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12312" *) alu_loop_op_unequal_tmp_7;
  assign _1197_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12314" *) FpAdd_8U_23U_int_mant_p1_2_lpi_1_dfm_5[49];
  assign nor_37_cse = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12314" *) _1489_;
  assign _1198_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12315" *) FpAdd_8U_23U_int_mant_p1_3_lpi_1_dfm_5[49];
  assign nor_41_cse = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12315" *) _1490_;
  assign _1199_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12316" *) FpAdd_8U_23U_int_mant_p1_lpi_1_dfm_5[49];
  assign nor_45_cse = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12316" *) _1491_;
  assign _1200_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12324" *) IsNaN_8U_23U_1_land_lpi_1_dfm_8;
  assign _1201_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12333" *) and_564_cse;
  assign nand_109_cse = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12333" *) _0495_;
  assign nor_430_cse = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12334" *) _1494_;
  assign _1202_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12336" *) FpAlu_8U_23U_nor_dfs_5;
  assign _1203_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12337" *) main_stage_v_3;
  assign nor_290_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12338" *) _1499_;
  assign nor_291_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12340" *) _1501_;
  assign _1204_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12342" *) FpAlu_8U_23U_equal_tmp_23;
  assign nor_293_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12342" *) _1502_;
  assign _1205_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12343" *) FpAlu_8U_23U_nor_dfs_6;
  assign _1206_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12345" *) main_stage_v_4;
  assign nor_292_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12346" *) _1505_;
  assign _1207_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12349" *) mux_109_itm;
  assign _1208_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12356" *) mux_111_nl;
  assign _1209_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12364" *) IsNaN_8U_23U_1_land_3_lpi_1_dfm_8;
  assign _1210_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12380" *) IsNaN_8U_23U_1_land_2_lpi_1_dfm_8;
  assign _1211_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12396" *) IsNaN_8U_23U_1_land_1_lpi_1_dfm_8;
  assign _1212_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12408" *) mux_124_nl;
  assign _1213_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12409" *) FpAlu_8U_23U_equal_tmp_26;
  assign _1214_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12416" *) mux_126_nl;
  assign _1215_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12417" *) alu_loop_op_3_FpMantRNE_49U_24U_else_and_1_tmp;
  assign _1216_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12418" *) FpAlu_8U_23U_equal_tmp_29;
  assign _1217_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12421" *) mux_129_nl;
  assign _1218_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12422" *) alu_loop_op_2_FpMantRNE_49U_24U_else_and_2_tmp;
  assign _1219_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12423" *) alu_loop_op_1_FpMantRNE_49U_24U_else_and_tmp;
  assign nor_269_cse = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12424" *) or_1087_cse;
  assign nor_397_cse = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12425" *) _1514_;
  assign _1220_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12429" *) alu_loop_op_4_FpMantRNE_49U_24U_else_and_3_tmp;
  assign _1221_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12432" *) mux_143_itm;
  assign _1222_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12434" *) mux_144_nl;
  assign _1223_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12435" *) or_dcpl_85;
  assign nor_264_cse = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12437" *) _1523_;
  assign _1224_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12439" *) _1524_;
  assign _1225_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12441" *) or_dcpl_86;
  assign _1226_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12442" *) or_dcpl_89;
  assign _1227_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12447" *) mux_tmp_146;
  assign nand_29_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12447" *) _0499_;
  assign _1228_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12450" *) mux_168_nl;
  assign _1229_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12451" *) or_dcpl_100;
  assign nor_71_cse = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12454" *) _1527_;
  assign _1230_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12456" *) _0504_;
  assign _1231_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12458" *) FpCmp_8U_23U_true_if_acc_4_nl[8];
  assign _1232_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12460" *) FpCmp_8U_23U_true_if_acc_6_nl[8];
  assign _1233_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12462" *) FpCmp_8U_23U_true_if_acc_8_nl[8];
  assign _1234_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12464" *) FpCmp_8U_23U_true_if_acc_10_nl[8];
  assign _1235_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12465" *) FpAlu_8U_23U_nor_dfs_4;
  assign nor_241_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12467" *) _1532_;
  assign _1236_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12471" *) _0509_;
  assign nor_243_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12471" *) _1534_;
  assign _1237_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12474" *) alu_loop_op_unequal_tmp_6;
  assign _1238_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12481" *) mux_184_nl;
  assign _1239_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12482" *) mux_tmp_171;
  assign _1240_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12485" *) FpAlu_8U_23U_equal_tmp_25;
  assign _1241_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12489" *) mux_192_nl;
  assign _1242_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12492" *) FpAlu_8U_23U_equal_tmp_28;
  assign _1243_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12494" *) FpAlu_8U_23U_equal_tmp_27;
  assign _1244_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12496" *) mux_198_nl;
  assign nor_236_cse = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12497" *) or_tmp_395;
  assign _1245_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12504" *) mux_202_nl;
  assign _0009_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12511" *) io_read_cfg_alu_bypass_rsc_svs_5;
  assign _1246_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12517" *) or_dcpl_109;
  assign _1247_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12517" *) mux_216_nl;
  assign _1248_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12519" *) cfg_alu_bypass_rsc_triosy_obj_bawt;
  assign _1249_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12519" *) cfg_alu_src_rsc_triosy_obj_bawt;
  assign _1250_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12520" *) cfg_alu_op_rsc_triosy_obj_bawt;
  assign _1251_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12520" *) cfg_alu_algo_rsc_triosy_obj_bawt;
  assign nor_208_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12521" *) _1556_;
  assign _1252_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12524" *) _0521_;
  assign nor_210_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12524" *) _1558_;
  assign nor_202_cse = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12532" *) or_963_cse;
  assign nor_204_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12532" *) _1559_;
  assign _1253_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12533" *) _1560_;
  assign _1254_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12539" *) or_tmp_402;
  assign nor_205_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12539" *) _1563_;
  assign nor_201_cse = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12546" *) _1572_;
  assign _1255_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12548" *) FpAlu_8U_23U_equal_tmp_24;
  assign nor_200_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12548" *) _1574_;
  assign nor_197_cse = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12552" *) _1573_;
  assign _0000_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12565" *) mux_tmp_227;
  assign _1256_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12570" *) mux_247_nl;
  assign _0001_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12578" *) mux_tmp_246;
  assign _0003_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12583" *) mux_266_nl;
  assign _1258_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12588" *) mux_270_nl;
  assign nor_177_cse = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12590" *) _1577_;
  assign _1259_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12600" *) mux_307_nl;
  assign _0004_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12601" *) cfg_alu_algo_rsci_d[0];
  assign _1260_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12622" *) _1581_;
  assign _1261_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12624" *) FpAdd_8U_23U_is_inf_3_lpi_1_dfm_8;
  assign _1262_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12628" *) IsNaN_8U_23U_land_3_lpi_1_dfm_11;
  assign nor_408_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12639" *) _1582_;
  assign alu_loop_op_4_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_3_svs_mx0w0 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12657" *) _2435_;
  assign _1263_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12658" *) FpAdd_8U_23U_is_a_greater_oif_aelse_acc_3_nl[23];
  assign alu_loop_op_3_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_1_svs_mx0w0 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12667" *) _2436_;
  assign _1264_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12668" *) FpAdd_8U_23U_is_a_greater_oif_aelse_acc_2_nl[23];
  assign alu_loop_op_2_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_2_svs_mx0w0 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12678" *) _2437_;
  assign _1265_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12679" *) FpAdd_8U_23U_is_a_greater_oif_aelse_acc_1_nl[23];
  assign alu_loop_op_1_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_mx0w0 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12689" *) _2438_;
  assign _1266_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12690" *) FpAdd_8U_23U_is_a_greater_oif_aelse_acc_nl[23];
  assign _1267_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12703" *) alu_loop_op_1_FpAdd_8U_23U_if_3_if_acc_1_nl[7];
  assign _0029_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12705" *) libraries_leading_sign_49_0_78e877fc94067377fcee479dbb0ed8e083a3_4;
  assign _0045_[8] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12707" *) FpAdd_8U_23U_if_3_if_and_tmp;
  assign nor_436_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12711" *) _1583_;
  assign _1268_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12715" *) alu_loop_op_2_FpAdd_8U_23U_if_3_if_acc_4_nl[7];
  assign _0030_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12717" *) libraries_leading_sign_49_0_78e877fc94067377fcee479dbb0ed8e083a3_5;
  assign _0046_[8] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12719" *) FpAdd_8U_23U_if_3_if_and_tmp_1;
  assign nor_435_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12723" *) _1584_;
  assign _1269_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12727" *) alu_loop_op_3_FpAdd_8U_23U_if_3_if_acc_2_nl[7];
  assign _0031_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12729" *) libraries_leading_sign_49_0_78e877fc94067377fcee479dbb0ed8e083a3_6;
  assign _0047_[8] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12731" *) FpAdd_8U_23U_if_3_if_and_tmp_2;
  assign nor_434_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12735" *) _1585_;
  assign _1270_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12739" *) alu_loop_op_4_FpAdd_8U_23U_if_3_if_acc_6_nl[7];
  assign _0032_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12741" *) libraries_leading_sign_49_0_78e877fc94067377fcee479dbb0ed8e083a3_7;
  assign _0048_[8] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12743" *) FpAdd_8U_23U_if_3_if_and_tmp_3;
  assign nor_433_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12747" *) _1586_;
  assign _1271_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12751" *) alu_loop_op_3_FpAdd_8U_23U_if_4_if_acc_2_nl[7];
  assign _1272_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12752" *) alu_loop_op_2_FpAdd_8U_23U_if_4_if_acc_4_nl[7];
  assign _1273_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12753" *) alu_loop_op_1_FpAdd_8U_23U_if_4_if_acc_1_nl[7];
  assign _1274_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12754" *) alu_loop_op_4_FpAdd_8U_23U_if_4_if_acc_6_nl[7];
  assign IsNaN_8U_23U_1_land_lpi_1_dfm_mx0w0 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12759" *) _1310_;
  assign IsNaN_8U_23U_1_land_3_lpi_1_dfm_mx0w0 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12760" *) _1304_;
  assign IsNaN_8U_23U_1_land_2_lpi_1_dfm_mx0w0 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12761" *) _1308_;
  assign IsNaN_8U_23U_1_land_1_lpi_1_dfm_mx0w0 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12762" *) _1306_;
  assign FpAlu_8U_23U_equal_tmp_mx0w0 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12765" *) _1149_;
  assign FpAlu_8U_23U_nor_dfs_mx0w0 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12767" *) _1588_;
  assign { _0041_[2], _0041_[0] } = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12779" *) alu_loop_op_else_o_32_1_2_lpi_1_dfm_mx0w0[31:30];
  assign { _0042_[2], _0042_[0] } = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12793" *) alu_loop_op_else_o_32_1_lpi_1_dfm_mx0w0[31:30];
  assign { _0043_[2], _0043_[0] } = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12797" *) alu_loop_op_else_o_32_1_3_lpi_1_dfm_mx0w0[31:30];
  assign { _0044_[2], _0044_[0] } = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12801" *) alu_loop_op_else_o_32_1_1_lpi_1_dfm_mx0w0[31:30];
  assign IsNaN_8U_23U_2_IsNaN_8U_23U_2_nor_2_itm_mx0w0 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12810" *) _1589_;
  assign _1275_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12811" *) _1160_;
  assign IsNaN_8U_23U_2_IsNaN_8U_23U_2_nor_itm_mx0w0 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12812" *) _1590_;
  assign _1276_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12813" *) _1162_;
  assign IsNaN_8U_23U_2_IsNaN_8U_23U_2_nor_1_itm_mx0w0 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12814" *) _1591_;
  assign IsNaN_8U_23U_2_IsNaN_8U_23U_2_nor_3_itm_mx0w0 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12816" *) _1592_;
  assign alu_loop_op_else_nor_dfs = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12818" *) _1594_;
  assign IsNaN_8U_23U_4_IsNaN_8U_23U_4_nand_3_itm_mx0w2 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12820" *) _1138_;
  assign IsNaN_8U_23U_4_IsNaN_8U_23U_4_nand_2_itm_mx0w2 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12821" *) _1139_;
  assign _1277_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12823" *) FpCmp_8U_23U_false_else_if_acc_6_nl[8];
  assign IsNaN_8U_23U_2_nor_3_mx0w0 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12826" *) _1164_;
  assign IsNaN_8U_23U_2_nor_2_mx0w0 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12827" *) _1165_;
  assign _1278_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12973" *) _1691_;
  assign _1279_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12975" *) FpAdd_8U_23U_is_inf_lpi_1_dfm_8;
  assign _1280_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12979" *) IsNaN_8U_23U_land_lpi_1_dfm_11;
  assign FpAdd_8U_23U_FpAdd_8U_23U_nor_11_m1c = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12993" *) or_962_nl;
  assign FpAdd_8U_23U_FpAdd_8U_23U_nor_9_m1c = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12995" *) _1692_;
  assign FpAdd_8U_23U_FpAdd_8U_23U_nor_7_m1c = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12997" *) _1693_;
  assign FpAdd_8U_23U_FpAdd_8U_23U_nor_5_m1c = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12999" *) _1694_;
  assign _1281_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13000" *) FpAlu_8U_23U_equal_tmp_32;
  assign _1282_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13002" *) FpAlu_8U_23U_and_12_tmp;
  assign _1283_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13006" *) _0554_;
  assign _0017_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13012" *) AluIn_data_sva_127[31:0];
  assign _0018_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13013" *) else_AluOp_data_0_lpi_1_dfm_mx0;
  assign _0019_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13024" *) AluIn_data_sva_127[63:32];
  assign _0020_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13025" *) else_AluOp_data_1_lpi_1_dfm_mx0;
  assign _0021_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13036" *) AluIn_data_sva_127[95:64];
  assign _0022_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13037" *) else_AluOp_data_2_lpi_1_dfm_mx0;
  assign _0023_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13048" *) AluIn_data_sva_127[127:96];
  assign _0024_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13049" *) else_AluOp_data_3_lpi_1_dfm_mx0;
  assign IntSaturation_33U_32U_IntSaturation_33U_32U_nor_1_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13075" *) _1700_;
  assign _1284_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13077" *) alu_loop_op_2_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_1_svs_3;
  assign IntSaturation_33U_32U_IntSaturation_33U_32U_nor_3_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13082" *) _1701_;
  assign _1285_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13084" *) alu_loop_op_4_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_1_svs_2;
  assign IntSaturation_33U_32U_IntSaturation_33U_32U_nor_2_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13089" *) _1702_;
  assign _1286_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13091" *) alu_loop_op_3_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_svs_2;
  assign IntSaturation_33U_32U_IntSaturation_33U_32U_nor_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13096" *) _1703_;
  assign _1287_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13098" *) alu_loop_op_1_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_svs_2;
  assign _0039_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13119" *) else_AluOp_data_0_lpi_1_dfm_mx0[30:23];
  assign _0049_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13122" *) AluIn_data_sva_127[22:0];
  assign _1288_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13125" *) FpCmp_8U_23U_true_else_else_if_acc_8_nl[23];
  assign _1289_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13125" *) _1704_;
  assign _1290_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13126" *) or_tmp_668;
  assign nor_168_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13126" *) _1705_;
  assign _1291_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13132" *) FpCmp_8U_23U_true_else_else_if_acc_4_nl[23];
  assign _1292_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13132" *) _1707_;
  assign _0005_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13134" *) else_mux_1_tmp_31_23[8];
  assign _1293_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13137" *) _1708_;
  assign _0050_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13141" *) AluIn_data_sva_127[86:64];
  assign _0035_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13144" *) else_AluOp_data_2_lpi_1_dfm_mx0[30:23];
  assign _1294_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13146" *) FpCmp_8U_23U_true_else_else_if_acc_7_nl[23];
  assign _1295_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13147" *) _1710_;
  assign _1296_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13148" *) or_tmp_674;
  assign nor_165_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13148" *) _1711_;
  assign _0051_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13155" *) AluIn_data_sva_127[118:96];
  assign _0033_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13158" *) else_AluOp_data_3_lpi_1_dfm_mx0[30:23];
  assign _1297_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13160" *) FpCmp_8U_23U_true_else_else_if_acc_6_nl[23];
  assign _1298_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13161" *) _1713_;
  assign _1299_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13162" *) or_tmp_678;
  assign nor_163_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13162" *) _1714_;
  assign nor_162_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13169" *) _1716_;
  assign nor_159_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13175" *) _1717_;
  assign _1300_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13178" *) _1718_;
  assign nor_156_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13182" *) _1719_;
  assign _1301_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13185" *) _1720_;
  assign _1302_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13188" *) FpCmp_8U_23U_false_is_abs_a_greater_2_lpi_1_dfm_1_mx0;
  assign _1303_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13195" *) IsNaN_8U_23U_2_IsNaN_8U_23U_2_nor_itm_2;
  assign _1305_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13199" *) IsNaN_8U_23U_land_3_lpi_1_dfm_8;
  assign _1307_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13201" *) IsNaN_8U_23U_land_1_lpi_1_dfm_8;
  assign _1309_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13203" *) IsNaN_8U_23U_land_2_lpi_1_dfm_8;
  assign _1311_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13205" *) IsNaN_8U_23U_land_lpi_1_dfm_8;
  assign _1136_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13206" *) FpAdd_8U_23U_qr_2_lpi_1_dfm_7;
  assign _1312_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13211" *) FpAdd_8U_23U_qr_3_lpi_1_dfm_7;
  assign _1313_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13216" *) FpAdd_8U_23U_qr_4_lpi_1_dfm_7;
  assign _1137_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13221" *) FpAdd_8U_23U_qr_lpi_1_dfm_7;
  assign _1314_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13226" *) io_read_cfg_alu_bypass_rsc_svs_8;
  assign _0040_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13228" *) AluIn_data_sva_127[30:23];
  assign IsNaN_8U_23U_3_nor_4_tmp = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13231" *) _1154_;
  assign _0038_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13233" *) AluIn_data_sva_127[62:55];
  assign _0037_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13237" *) else_AluOp_data_1_lpi_1_dfm_mx2_30_0[30:23];
  assign IsNaN_8U_23U_3_nor_6_tmp = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13240" *) _1152_;
  assign _0052_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13244" *) AluIn_data_sva_127[54:32];
  assign _0036_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13248" *) AluIn_data_sva_127[94:87];
  assign IsNaN_8U_23U_3_nor_8_tmp = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13251" *) _1150_;
  assign _0034_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13253" *) AluIn_data_sva_127[126:119];
  assign IsNaN_8U_23U_3_nor_10_tmp = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13256" *) _1166_;
  assign _1315_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13274" *) _1724_;
  assign _1316_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13280" *) _1167_;
  assign _1317_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13286" *) and_37_cse;
  assign nand_17_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13286" *) _0562_;
  assign _0006_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13288" *) mux_32_nl;
  assign not_tmp_24 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13290" *) _0563_;
  assign _1318_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13295" *) _0568_;
  assign nor_371_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13295" *) _1727_;
  assign nor_372_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13297" *) _1728_;
  assign not_tmp_38 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13300" *) _1729_;
  assign nor_357_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13305" *) _1733_;
  assign _0007_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13306" *) or_tmp_75;
  assign _1319_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13323" *) FpAlu_8U_23U_equal_tmp_31;
  assign _1320_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13329" *) FpAlu_8U_23U_equal_tmp_34;
  assign _1321_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13332" *) _1740_;
  assign _1322_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13334" *) alu_loop_op_unequal_tmp_8;
  assign not_tmp_152 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13345" *) or_632_cse;
  assign nor_248_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13347" *) _1759_;
  assign _1323_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13352" *) mux_162_nl;
  assign nand_tmp_13 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13352" *) _0569_;
  assign nor_379_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13354" *) _1760_;
  assign nor_187_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13388" *) _1766_;
  assign _0008_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13395" *) cfg_alu_algo_1_sva_st_22[0];
  assign _1324_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13412" *) mux_254_nl;
  assign nand_tmp_20 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13412" *) _0002_;
  assign _0010_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13421" *) mux_tmp_237;
  assign not_tmp_259 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13424" *) _0576_;
  assign _1325_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13427" *) or_tmp_597;
  assign not_tmp_261 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13427" *) _1773_;
  assign _0012_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13428" *) cfg_alu_algo_1_sva_st[0];
  assign _0011_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13432" *) cfg_alu_algo_1_sva_st_22[1];
  assign _1326_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13447" *) _0577_;
  assign or_dcpl_14 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13447" *) _0578_;
  assign _1327_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13450" *) _0580_;
  assign _1328_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13450" *) _0581_;
  assign _1329_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13451" *) chn_alu_out_rsci_bawt;
  assign _1330_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13452" *) chn_alu_op_rsci_bawt;
  assign or_dcpl_20 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13455" *) and_486_cse;
  assign _1331_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13462" *) cfg_alu_bypass_rsci_d;
  assign _1332_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13493" *) cfg_precision[1];
  assign _1333_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13495" *) alu_loop_op_1_FpAdd_8U_23U_is_a_greater_oif_equal_tmp;
  assign _1334_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13497" *) alu_loop_op_2_FpAdd_8U_23U_is_a_greater_oif_equal_2_tmp;
  assign _1335_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13499" *) alu_loop_op_3_FpAdd_8U_23U_is_a_greater_oif_equal_1_tmp;
  assign _1336_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13501" *) alu_loop_op_4_FpAdd_8U_23U_is_a_greater_oif_equal_3_tmp;
  assign _1337_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13505" *) cfg_precision[0];
  assign _1338_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13508" *) io_read_cfg_alu_bypass_rsc_svs_6;
  assign _1339_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13509" *) cfg_alu_algo_1_sva_st_23[1];
  assign and_dcpl_175 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13512" *) _1796_;
  assign mux_tmp_323 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13518" *) _1257_;
  assign _1340_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13521" *) cfg_alu_algo_rsci_d[1];
  assign _1341_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13525" *) cfg_alu_algo_1_sva_st[1];
  assign _1342_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13543" *) cfg_alu_src_rsci_d;
  assign _0053_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13561" *) else_AluOp_data_0_lpi_1_dfm_mx0[22:0];
  assign _0054_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13565" *) else_AluOp_data_1_lpi_1_dfm_mx0[22:0];
  assign _0055_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13569" *) else_AluOp_data_2_lpi_1_dfm_mx0[22:0];
  assign _0056_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13573" *) else_AluOp_data_3_lpi_1_dfm_mx0[22:0];
  assign _1343_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13596" *) or_dcpl_123;
  assign _1344_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13596" *) _1800_;
  assign _1345_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13598" *) or_dcpl_121;
  assign _1346_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13598" *) _1801_;
  assign _1347_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13600" *) or_dcpl_119;
  assign _1348_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13600" *) _1802_;
  assign _1349_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13602" *) or_dcpl_117;
  assign _1350_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13602" *) _1803_;
  assign _1351_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13628" *) main_stage_en_1;
  assign _1352_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13628" *) _0630_;
  assign _1353_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13721" *) and_dcpl_45;
  assign _1354_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13730" *) chn_alu_op_rsci_ld_core_psct_mx0c1;
  assign _1355_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13738" *) main_stage_v_1_mx0c1;
  assign _1356_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13763" *) mux_23_nl;
  assign _1357_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13771" *) mux_31_nl;
  assign _1358_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13779" *) mux_34_itm;
  assign _1359_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13809" *) _1812_;
  assign _1360_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13818" *) main_stage_v_2_mx0c1;
  assign _1361_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13948" *) and_dcpl_77;
  assign _1362_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13961" *) main_stage_v_3_mx0c1;
  assign _1363_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14090" *) main_stage_v_4_mx0c1;
  assign _1364_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14192" *) FpAlu_8U_23U_equal_tmp_22;
  assign _1365_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14193" *) io_read_cfg_alu_bypass_rsc_svs_st_6;
  assign _1366_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14355" *) mux_127_nl;
  assign _1367_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14438" *) mux_133_nl;
  assign _1368_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14446" *) mux_135_nl;
  assign _1369_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14455" *) _1836_;
  assign _1370_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14455" *) _1837_;
  assign _1371_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14464" *) mux_136_nl;
  assign _1372_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14500" *) mux_138_nl;
  assign _1373_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14508" *) mux_139_nl;
  assign _1374_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14788" *) mux_172_nl;
  assign _1375_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14796" *) _1839_;
  assign _1376_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14804" *) _1841_;
  assign _1377_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14879" *) mux_182_nl;
  assign _1378_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14920" *) mux_190_nl;
  assign _1379_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14940" *) mux_194_nl;
  assign _1380_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14948" *) mux_196_nl;
  assign _1381_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14966" *) mux_tmp_173;
  assign _1382_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15095" *) _1852_;
  assign _1383_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15104" *) _1853_;
  assign _1384_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15113" *) _1854_;
  assign _1385_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15122" *) _1855_;
  assign _1386_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15154" *) FpAlu_8U_23U_equal_tmp_1_mx0w0;
  assign _1387_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15294" *) alu_loop_op_1_IntSaturation_33U_32U_if_acc_nl[2];
  assign _1388_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15305" *) _1860_;
  assign _1389_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15315" *) alu_loop_op_2_IntSaturation_33U_32U_if_acc_1_nl[2];
  assign _1390_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15326" *) _1861_;
  assign _1391_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15348" *) alu_loop_op_3_IntSaturation_33U_32U_if_acc_nl[2];
  assign _1392_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15359" *) mux_365_nl;
  assign _1393_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15372" *) _1863_;
  assign _1394_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15381" *) _1864_;
  assign _1395_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15432" *) mux_175_nl;
  assign _1396_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15475" *) _1870_;
  assign _1397_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15475" *) mux_277_nl;
  assign _1398_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15483" *) mux_290_nl;
  assign _1399_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15494" *) mux_303_nl;
  assign _1400_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15506" *) mux_305_nl;
  assign _1401_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15534" *) mux_314_nl;
  assign _1402_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15566" *) _1872_;
  assign _1403_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15568" *) FpAdd_8U_23U_is_inf_1_lpi_1_dfm_8;
  assign _1404_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15572" *) IsNaN_8U_23U_land_1_lpi_1_dfm_11;
  assign nor_406_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15582" *) _1873_;
  assign _1405_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15586" *) _1874_;
  assign _1406_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15588" *) FpAdd_8U_23U_is_inf_2_lpi_1_dfm_8;
  assign _1407_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15592" *) IsNaN_8U_23U_land_2_lpi_1_dfm_11;
  assign nor_407_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15602" *) _1875_;
  assign _0013_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15603" *) mux_tmp_2;
  assign _0014_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15609" *) mux_tmp_10;
  assign _1408_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15616" *) or_tmp_23;
  assign nand_18_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15616" *) _0892_;
  assign _0015_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15618" *) alu_loop_op_2_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_1_svs_2;
  assign _1409_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15625" *) _1876_;
  assign nor_354_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15628" *) _1880_;
  assign nor_355_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15630" *) _1883_;
  assign nor_356_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15633" *) _1885_;
  assign nor_351_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15636" *) _1888_;
  assign nor_352_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15638" *) _1891_;
  assign nor_353_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15641" *) _1892_;
  assign nor_348_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15644" *) _1895_;
  assign nor_349_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15646" *) _1898_;
  assign nor_350_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15649" *) _1899_;
  assign nor_345_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15652" *) _1902_;
  assign nor_346_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15654" *) _1905_;
  assign nor_347_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15657" *) _1906_;
  assign nor_344_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15660" *) _1908_;
  assign _0016_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15661" *) or_tmp_103;
  assign nor_336_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15665" *) _1914_;
  assign nor_337_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15668" *) _1920_;
  assign nor_338_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15674" *) _1925_;
  assign _1410_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15677" *) _1926_;
  assign nor_334_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15677" *) _1927_;
  assign _1411_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15678" *) alu_loop_op_1_FpMantRNE_49U_24U_else_and_svs_st_2;
  assign _1412_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15679" *) alu_loop_op_1_FpAdd_8U_23U_if_4_if_slc_FpAdd_8U_23U_if_4_if_acc_1_7_svs_st_3;
  assign _1413_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15682" *) _1935_;
  assign nor_340_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15682" *) _1936_;
  assign _1414_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15685" *) _1942_;
  assign nor_342_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15686" *) _1943_;
  assign nor_339_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15688" *) _1944_;
  assign nor_326_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15692" *) _1950_;
  assign nor_327_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15695" *) _1956_;
  assign nor_328_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15701" *) _1959_;
  assign _1415_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15704" *) _1960_;
  assign nor_324_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15704" *) _1961_;
  assign _1416_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15705" *) alu_loop_op_2_FpMantRNE_49U_24U_else_and_2_svs_st_2;
  assign _1417_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15706" *) alu_loop_op_2_FpAdd_8U_23U_if_4_if_slc_FpAdd_8U_23U_if_4_if_acc_1_7_2_svs_st_3;
  assign _1418_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15709" *) _1969_;
  assign nor_330_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15709" *) _1970_;
  assign _1419_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15712" *) _1976_;
  assign nor_332_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15713" *) _1977_;
  assign nor_329_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15715" *) _1978_;
  assign nor_316_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15719" *) _1984_;
  assign nor_317_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15722" *) _1990_;
  assign nor_318_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15728" *) _1993_;
  assign _1420_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15731" *) _1994_;
  assign nor_314_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15731" *) _1995_;
  assign _1421_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15732" *) alu_loop_op_3_FpMantRNE_49U_24U_else_and_1_svs_st_2;
  assign _1422_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15733" *) alu_loop_op_3_FpAdd_8U_23U_if_4_if_slc_FpAdd_8U_23U_if_4_if_acc_1_7_1_svs_st_3;
  assign _1423_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15736" *) _2003_;
  assign nor_320_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15736" *) _2004_;
  assign _1424_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15739" *) _2010_;
  assign nor_322_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15740" *) _2011_;
  assign nor_319_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15742" *) _2012_;
  assign nor_310_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15747" *) _2021_;
  assign nor_311_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15751" *) _2030_;
  assign nor_312_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15758" *) _2037_;
  assign _1425_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15760" *) alu_loop_op_4_FpMantRNE_49U_24U_else_and_3_svs_st_2;
  assign _1426_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15761" *) alu_loop_op_4_FpAdd_8U_23U_if_4_if_slc_FpAdd_8U_23U_if_4_if_acc_1_7_3_svs_st_3;
  assign nor_313_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15767" *) _2045_;
  assign nor_307_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15770" *) _2048_;
  assign _1427_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15771" *) alu_loop_op_1_FpMantRNE_49U_24U_else_and_svs_st;
  assign nor_308_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15772" *) _2051_;
  assign _1428_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15775" *) _0893_;
  assign nor_309_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15775" *) _2053_;
  assign nor_304_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15778" *) _2056_;
  assign _1429_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15779" *) alu_loop_op_2_FpMantRNE_49U_24U_else_and_2_svs_st;
  assign nor_305_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15780" *) _2059_;
  assign _1430_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15783" *) _0894_;
  assign nor_306_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15783" *) _2060_;
  assign nor_301_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15786" *) _2063_;
  assign _1431_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15787" *) alu_loop_op_3_FpMantRNE_49U_24U_else_and_1_svs_st;
  assign nor_302_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15788" *) _2066_;
  assign _1432_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15791" *) _0895_;
  assign nor_303_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15791" *) _2067_;
  assign nor_298_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15794" *) _2070_;
  assign _1433_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15795" *) alu_loop_op_4_FpMantRNE_49U_24U_else_and_3_svs_st;
  assign nor_299_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15796" *) _2073_;
  assign _1434_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15799" *) _0896_;
  assign nor_300_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15799" *) _2074_;
  assign _1435_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15803" *) _2076_;
  assign nor_274_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15811" *) _2084_;
  assign _1436_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15814" *) IsNaN_8U_23U_1_land_3_lpi_1_dfm_9;
  assign nor_275_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15814" *) _2086_;
  assign nor_272_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15818" *) _2088_;
  assign _1437_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15821" *) IsNaN_8U_23U_1_land_2_lpi_1_dfm_9;
  assign nor_273_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15821" *) _2090_;
  assign nor_270_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15825" *) _2092_;
  assign _1438_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15828" *) IsNaN_8U_23U_1_land_1_lpi_1_dfm_9;
  assign nor_271_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15828" *) _2094_;
  assign _1439_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15845" *) FpAlu_8U_23U_equal_tmp_35;
  assign nor_267_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15851" *) _2114_;
  assign _1440_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15854" *) IsNaN_8U_23U_1_land_lpi_1_dfm_9;
  assign nor_268_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15854" *) _2116_;
  assign _1441_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15858" *) nor_tmp_144;
  assign _1442_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15868" *) or_tmp_315;
  assign nor_263_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15882" *) _2127_;
  assign nor_265_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15887" *) _2131_;
  assign nor_260_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15892" *) _2138_;
  assign nor_262_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15897" *) _2142_;
  assign nor_257_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15902" *) _2149_;
  assign nor_259_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15907" *) _2153_;
  assign nor_254_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15912" *) _2160_;
  assign nor_256_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15917" *) _2164_;
  assign nor_252_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15920" *) _2167_;
  assign _1443_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15921" *) acc_12_nl[50];
  assign nor_251_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15925" *) _2172_;
  assign _1444_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15926" *) acc_13_nl[50];
  assign nor_250_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15930" *) _2177_;
  assign _1445_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15931" *) acc_14_nl[50];
  assign nor_249_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15935" *) _2182_;
  assign _1446_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15936" *) acc_15_nl[50];
  assign _1447_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15943" *) alu_loop_op_1_IntSaturation_33U_32U_else_if_acc_nl[2];
  assign _1448_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15946" *) FpAlu_8U_23U_equal_tmp_21;
  assign _1449_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15950" *) alu_loop_op_4_IntSaturation_33U_32U_else_if_acc_1_nl[2];
  assign _1450_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15952" *) alu_loop_op_3_IntSaturation_33U_32U_else_if_acc_nl[2];
  assign _1451_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15954" *) alu_loop_op_2_IntSaturation_33U_32U_else_if_acc_1_nl[2];
  assign _1452_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15966" *) FpAlu_8U_23U_equal_tmp_33;
  assign _1453_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15967" *) FpAlu_8U_23U_equal_tmp_30;
  assign _1454_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15977" *) IsNaN_8U_23U_1_land_3_lpi_1_dfm_7;
  assign nor_237_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15978" *) _2206_;
  assign _1455_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15982" *) _2210_;
  assign _1456_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15982" *) _2211_;
  assign nor_238_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15982" *) _2212_;
  assign _1457_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15985" *) IsNaN_8U_23U_1_land_lpi_1_dfm_7;
  assign nor_232_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15986" *) _2216_;
  assign _1458_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15990" *) _2218_;
  assign _1459_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15990" *) _2219_;
  assign nor_233_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15990" *) _2220_;
  assign _1460_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15993" *) IsNaN_8U_23U_1_land_2_lpi_1_dfm_7;
  assign nor_227_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15994" *) _2224_;
  assign _1461_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15998" *) _2226_;
  assign _1462_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15998" *) _2227_;
  assign nor_228_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15998" *) _2228_;
  assign _1463_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16001" *) IsNaN_8U_23U_1_land_1_lpi_1_dfm_7;
  assign nor_222_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16002" *) _2232_;
  assign _1464_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16006" *) _2234_;
  assign _1465_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16006" *) _2235_;
  assign nor_223_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16006" *) _2236_;
  assign nor_219_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16013" *) _2242_;
  assign nor_220_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16017" *) _2248_;
  assign nor_217_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16022" *) _2254_;
  assign nor_218_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16026" *) _2260_;
  assign nor_215_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16031" *) _2266_;
  assign nor_216_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16035" *) _2272_;
  assign nor_213_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16040" *) _2278_;
  assign nor_214_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16044" *) _2284_;
  assign _1466_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16046" *) FpAdd_8U_23U_is_a_greater_lor_1_lpi_1_dfm_1_mx0w0;
  assign _1467_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16054" *) FpAdd_8U_23U_is_a_greater_lor_2_lpi_1_dfm_1_mx0w0;
  assign nor_207_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16063" *) _2285_;
  assign nor_206_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16066" *) _2286_;
  assign nor_203_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16089" *) _2287_;
  assign nor_195_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16095" *) _2293_;
  assign nor_192_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16101" *) _2299_;
  assign _1468_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16114" *) FpAdd_8U_23U_is_a_greater_lor_lpi_1_dfm_1_mx0w0;
  assign _1469_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16128" *) FpAdd_8U_23U_is_a_greater_lor_3_lpi_1_dfm_1_mx0w0;
  assign _1470_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16141" *) nor_tmp_74;
  assign nand_30_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16141" *) _0927_;
  assign _1471_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16145" *) _2305_;
  assign nor_178_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16157" *) _2307_;
  assign nand_35_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16159" *) _0928_;
  assign _1472_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16163" *) mux_289_nl;
  assign nand_36_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16163" *) _0929_;
  assign nor_176_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16168" *) _2308_;
  assign nand_37_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16170" *) _0930_;
  assign _1473_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16174" *) mux_302_nl;
  assign nand_38_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16174" *) _0931_;
  assign _0025_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16212" *) FpAdd_8U_23U_addend_smaller_qr_1_lpi_1_dfm_mx0;
  assign _1474_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16216" *) FpAdd_8U_23U_if_2_and_tmp;
  assign _0026_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16221" *) FpAdd_8U_23U_addend_smaller_qr_2_lpi_1_dfm_mx0;
  assign _1475_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16225" *) FpAdd_8U_23U_if_2_and_tmp_1;
  assign _0027_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16230" *) FpAdd_8U_23U_addend_smaller_qr_3_lpi_1_dfm_mx0;
  assign _1476_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16234" *) FpAdd_8U_23U_if_2_and_tmp_2;
  assign _0028_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16239" *) FpAdd_8U_23U_addend_smaller_qr_lpi_1_dfm_mx0;
  assign _1477_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16243" *) FpAdd_8U_23U_if_2_and_tmp_3;
  assign chn_alu_out_or_cse = _0480_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12265" *) and_dcpl_40;
  assign _1478_ = asn_267 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12268" *) or_dcpl;
  assign or_1087_cse = _1183_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12269" *) chn_alu_out_rsci_bawt;
  assign _1479_ = or_dcpl_272 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12270" *) FpAlu_8U_23U_nor_dfs_6;
  assign _1480_ = _1479_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12271" *) FpAlu_8U_23U_equal_tmp_23;
  assign _1481_ = _1480_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12271" *) io_read_cfg_alu_bypass_rsc_svs_8;
  assign _1482_ = _1481_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12271" *) alu_loop_op_unequal_tmp_8;
  assign _1483_ = nor_269_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12275" *) chn_alu_in_rsci_bawt;
  assign _1484_ = _1483_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12275" *) _1185_;
  assign or_tmp_386 = cfg_alu_bypass_rsci_d | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12280" *) _1188_;
  assign or_28_cse = _1147_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12281" *) cfg_alu_algo_1_sva_st[1];
  assign cfg_alu_algo_cfg_alu_algo_or_3_cse = _0485_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12282" *) and_dcpl_81;
  assign or_963_cse = _1189_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12285" *) chn_alu_op_rsci_bawt;
  assign or_16_cse = or_963_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12285" *) io_read_cfg_alu_bypass_rsc_svs_st_1;
  assign FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_or_7_cse = and_dcpl_78 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12293" *) and_dcpl_99;
  assign _1485_ = _1192_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12297" *) io_read_cfg_alu_bypass_rsc_svs_st_1;
  assign _1486_ = _1485_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12298" *) _1193_;
  assign _1487_ = _1194_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12299" *) io_read_cfg_alu_bypass_rsc_svs_st_5;
  assign FpAdd_8U_23U_int_mant_p1_or_3_cse = or_dcpl_86 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12307" *) and_dcpl_99;
  assign _1488_ = alu_loop_op_1_FpAdd_8U_23U_if_3_if_acc_1_nl[7] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12311" *) _1195_;
  assign FpAdd_8U_23U_o_expo_FpAdd_8U_23U_o_expo_or_2_cse = _0494_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12313" *) and_dcpl_108;
  assign _1489_ = alu_loop_op_2_FpAdd_8U_23U_if_3_if_acc_4_nl[7] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12314" *) _1197_;
  assign _1490_ = alu_loop_op_3_FpAdd_8U_23U_if_3_if_acc_2_nl[7] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12315" *) _1198_;
  assign _1491_ = alu_loop_op_4_FpAdd_8U_23U_if_3_if_acc_6_nl[7] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12316" *) _1199_;
  assign _1492_ = IsNaN_8U_23U_land_lpi_1_dfm_11 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12328" *) _1183_;
  assign _1493_ = _1492_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12328" *) chn_alu_out_rsci_bawt;
  assign or_735_nl = _1493_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12328" *) io_read_cfg_alu_bypass_rsc_svs_8;
  assign _1494_ = alu_loop_op_unequal_tmp_7 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12334" *) io_read_cfg_alu_bypass_rsc_svs_st_6;
  assign _1495_ = _1148_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12337" *) _1202_;
  assign _1496_ = _1495_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12337" *) _1203_;
  assign _1497_ = _1496_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12337" *) io_read_cfg_alu_bypass_rsc_svs_st_6;
  assign _1498_ = _1497_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12338" *) io_read_cfg_alu_bypass_rsc_svs_7;
  assign _1499_ = _1498_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12338" *) alu_loop_op_unequal_tmp_7;
  assign or_tmp_103 = _1203_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12340" *) io_read_cfg_alu_bypass_rsc_svs_st_6;
  assign _1500_ = or_tmp_103 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12340" *) io_read_cfg_alu_bypass_rsc_svs_7;
  assign _1501_ = _1500_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12340" *) alu_loop_op_unequal_tmp_7;
  assign _1502_ = cfg_alu_algo_1_sva_st_25[1] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12342" *) _1204_;
  assign or_225_nl = _1205_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12343" *) cfg_alu_algo_1_sva_st_25[0];
  assign or_323_nl = _1206_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12345" *) io_read_cfg_alu_bypass_rsc_svs_8;
  assign _1503_ = or_323_nl | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12346" *) alu_loop_op_unequal_tmp_8;
  assign _1504_ = _1503_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12346" *) io_read_cfg_alu_bypass_rsc_svs_st_7;
  assign _1505_ = _1504_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12346" *) mux_106_nl;
  assign _1506_ = nor_269_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12350" *) _1148_;
  assign _1507_ = _1506_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12351" *) io_read_cfg_alu_bypass_rsc_svs_st_6;
  assign or_239_nl = _1507_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12351" *) _1203_;
  assign _1508_ = IsNaN_8U_23U_land_3_lpi_1_dfm_11 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12368" *) _1183_;
  assign _1509_ = _1508_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12368" *) chn_alu_out_rsci_bawt;
  assign or_741_nl = _1509_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12368" *) io_read_cfg_alu_bypass_rsc_svs_8;
  assign _1510_ = IsNaN_8U_23U_land_2_lpi_1_dfm_11 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12384" *) _1183_;
  assign _1511_ = _1510_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12384" *) chn_alu_out_rsci_bawt;
  assign or_744_nl = _1511_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12384" *) io_read_cfg_alu_bypass_rsc_svs_8;
  assign _1512_ = IsNaN_8U_23U_land_1_lpi_1_dfm_11 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12400" *) _1183_;
  assign _1513_ = _1512_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12400" *) chn_alu_out_rsci_bawt;
  assign or_747_nl = _1513_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12400" *) io_read_cfg_alu_bypass_rsc_svs_8;
  assign _1514_ = alu_loop_op_unequal_tmp_8 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12406" *) io_read_cfg_alu_bypass_rsc_svs_8;
  assign or_270_nl = _1514_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12406" *) _1206_;
  assign _1515_ = _1213_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12409" *) alu_loop_op_unequal_tmp_8;
  assign _1516_ = _1515_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12410" *) io_read_cfg_alu_bypass_rsc_svs_8;
  assign or_273_nl = _1516_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12410" *) _1206_;
  assign _1517_ = or_1087_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12413" *) _1213_;
  assign _1518_ = _1517_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12413" *) alu_loop_op_unequal_tmp_8;
  assign _1519_ = _1518_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12414" *) io_read_cfg_alu_bypass_rsc_svs_8;
  assign or_275_nl = _1519_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12414" *) _1206_;
  assign _1520_ = _1216_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12418" *) alu_loop_op_unequal_tmp_8;
  assign _1521_ = _1520_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12419" *) io_read_cfg_alu_bypass_rsc_svs_8;
  assign or_288_nl = _1521_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12419" *) _1206_;
  assign or_dcpl_272 = FpAlu_8U_23U_equal_tmp_29 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12426" *) FpAlu_8U_23U_equal_tmp_26;
  assign _1522_ = _1487_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12437" *) io_read_cfg_alu_bypass_rsc_svs_6;
  assign _1523_ = _1522_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12437" *) alu_loop_op_unequal_tmp_6;
  assign or_dcpl_127 = or_dcpl_91 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12439" *) and_dcpl_32;
  assign _1524_ = or_dcpl_127 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12439" *) io_read_cfg_alu_bypass_rsc_svs_st_5;
  assign _1525_ = nor_269_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12453" *) or_1050_cse;
  assign _1526_ = _1525_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12454" *) cfg_alu_bypass_rsci_d;
  assign _1527_ = _1526_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12454" *) _1188_;
  assign _1528_ = or_dcpl_86 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12466" *) _1235_;
  assign _1529_ = _1528_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12466" *) _1194_;
  assign _1530_ = _1529_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12466" *) io_read_cfg_alu_bypass_rsc_svs_st_5;
  assign _1531_ = _1530_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12467" *) io_read_cfg_alu_bypass_rsc_svs_6;
  assign _1532_ = _1531_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12467" *) alu_loop_op_unequal_tmp_6;
  assign _1533_ = cfg_alu_algo_1_sva_st_24[0] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12471" *) _1236_;
  assign _1534_ = _1501_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12471" *) _0510_;
  assign FpAlu_8U_23U_o_FpAlu_8U_23U_o_or_cse = _0511_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12475" *) and_dcpl_165;
  assign or_426_nl = or_1087_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12478" *) or_tmp_305;
  assign or_441_nl = alu_loop_op_unequal_tmp_6 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12483" *) or_tmp_416;
  assign _1535_ = _1240_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12486" *) _1183_;
  assign _1536_ = _1535_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12486" *) chn_alu_out_rsci_bawt;
  assign _1537_ = _1536_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12486" *) alu_loop_op_unequal_tmp_7;
  assign _1538_ = _1537_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12487" *) io_read_cfg_alu_bypass_rsc_svs_7;
  assign or_443_nl = _1538_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12487" *) _1203_;
  assign _1539_ = or_1087_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12492" *) _1242_;
  assign _1540_ = _1539_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12492" *) alu_loop_op_unequal_tmp_7;
  assign _1541_ = _1540_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12493" *) io_read_cfg_alu_bypass_rsc_svs_7;
  assign or_453_nl = _1541_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12493" *) _1203_;
  assign _1542_ = alu_loop_op_unequal_tmp_6 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12494" *) _1243_;
  assign or_tmp_395 = _1194_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12497" *) io_read_cfg_alu_bypass_rsc_svs_6;
  assign _1543_ = and_dcpl_165 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12499" *) and_dcpl_168;
  assign IntSaturation_33U_32U_IntSaturation_33U_32U_or_7_cse = _1543_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12499" *) and_dcpl_169;
  assign _1544_ = or_1087_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12502" *) _1196_;
  assign _1545_ = _1544_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12502" *) io_read_cfg_alu_bypass_rsc_svs_7;
  assign or_463_nl = _1545_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12502" *) _1203_;
  assign _1546_ = and_dcpl_170 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12508" *) alu_loop_bypass_if_and_6_cse;
  assign _1547_ = _1546_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12508" *) alu_loop_bypass_if_and_7_cse;
  assign _1548_ = or_1050_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12518" *) _1192_;
  assign _1549_ = _1548_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12519" *) io_read_cfg_alu_bypass_rsc_svs_st_1;
  assign _1550_ = _1549_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12519" *) _1248_;
  assign _1551_ = _1550_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12520" *) _1249_;
  assign _1552_ = _1551_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12520" *) _1250_;
  assign _1553_ = _1552_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12521" *) _1251_;
  assign _1554_ = _1553_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12521" *) io_read_cfg_alu_bypass_rsc_svs_5;
  assign _1555_ = _1554_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12521" *) FpAlu_8U_23U_equal_tmp_1_mx0w0;
  assign _1556_ = _1555_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12521" *) nor_202_cse;
  assign _1557_ = cfg_alu_algo_1_sva_st_23[0] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12524" *) _1252_;
  assign _1558_ = _1523_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12524" *) _0522_;
  assign _1559_ = cfg_precision[1] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12532" *) nor_202_cse;
  assign _1560_ = FpAlu_8U_23U_equal_tmp_1_mx0w0 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12533" *) cfg_precision[0];
  assign _1561_ = _1253_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12534" *) io_read_cfg_alu_bypass_rsc_svs_st_1;
  assign _1562_ = _1254_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12539" *) _1194_;
  assign _1563_ = _1562_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12539" *) io_read_cfg_alu_bypass_rsc_svs_6;
  assign _1564_ = nor_202_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12543" *) or_1050_cse;
  assign _1565_ = _1564_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12544" *) _1192_;
  assign _1566_ = _1565_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12544" *) io_read_cfg_alu_bypass_rsc_svs_st_1;
  assign _1567_ = _1566_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12545" *) _1248_;
  assign _1568_ = _1567_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12545" *) _1249_;
  assign _1569_ = _1568_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12546" *) _1250_;
  assign _1570_ = _1569_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12546" *) _1251_;
  assign _1571_ = _1570_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12546" *) _1149_;
  assign _1572_ = _1571_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12546" *) io_read_cfg_alu_bypass_rsc_svs_5;
  assign _1573_ = or_tmp_395 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12548" *) alu_loop_op_unequal_tmp_6;
  assign _1574_ = _1573_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12548" *) _1255_;
  assign FpAlu_8U_23U_or_cse = _0533_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12572" *) _0534_;
  assign _1575_ = and_dcpl_219 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12576" *) and_dcpl_81;
  assign _1576_ = _1575_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12577" *) and_dcpl_222;
  assign IsNaN_8U_23U_2_IsNaN_8U_23U_2_or_5_cse = _1576_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12577" *) and_dcpl_225;
  assign _1577_ = and_486_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12590" *) io_read_cfg_alu_bypass_rsc_svs_5;
  assign _1578_ = and_dcpl_222 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12591" *) and_dcpl_227;
  assign _1579_ = _1578_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12592" *) and_dcpl_229;
  assign IsNaN_8U_23U_2_IsNaN_8U_23U_4_or_2_cse = _1579_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12592" *) and_dcpl_231;
  assign _1580_ = and_dcpl_236 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12596" *) and_dcpl_239;
  assign IsNaN_8U_23U_2_IsNaN_8U_23U_2_or_3_cse = _1580_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12596" *) and_dcpl_243;
  assign _1581_ = FpAdd_8U_23U_and_2_tmp_3 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12622" *) FpAdd_8U_23U_is_inf_3_lpi_1_dfm_8;
  assign _1582_ = asn_267 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12639" *) or_998_tmp;
  assign FpAdd_8U_23U_is_a_greater_lor_lpi_1_dfm_1_mx0w0 = _0543_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12659" *) FpCmp_8U_23U_true_if_acc_10_nl[8];
  assign FpAdd_8U_23U_is_a_greater_lor_3_lpi_1_dfm_1_mx0w0 = _0544_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12669" *) FpCmp_8U_23U_true_if_acc_8_nl[8];
  assign alu_loop_op_3_FpAdd_8U_23U_IsZero_8U_23U_1_or_itm_mx0w0 = _1150_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12671" *) _1151_;
  assign FpAdd_8U_23U_is_a_greater_lor_2_lpi_1_dfm_1_mx0w0 = _0545_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12680" *) FpCmp_8U_23U_true_if_acc_6_nl[8];
  assign alu_loop_op_2_FpAdd_8U_23U_IsZero_8U_23U_1_or_itm_mx0w0 = _1152_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12682" *) _1153_;
  assign FpAdd_8U_23U_is_a_greater_lor_1_lpi_1_dfm_1_mx0w0 = _0546_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12691" *) FpCmp_8U_23U_true_if_acc_4_nl[8];
  assign alu_loop_op_1_FpAdd_8U_23U_IsZero_8U_23U_1_or_itm_mx0w0 = _1154_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12693" *) _1155_;
  assign _1583_ = FpAdd_8U_23U_and_4_tmp | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12711" *) mux_tmp;
  assign _1584_ = FpAdd_8U_23U_and_10_tmp | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12723" *) mux_tmp_348;
  assign _1585_ = FpAdd_8U_23U_and_16_tmp | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12735" *) mux_tmp_349;
  assign _1586_ = FpAdd_8U_23U_and_22_tmp | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12747" *) mux_tmp_350;
  assign FpAdd_8U_23U_is_inf_3_lpi_1_dfm_2_mx0w0 = nor_41_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12751" *) _1271_;
  assign FpAdd_8U_23U_is_inf_2_lpi_1_dfm_2_mx0w0 = nor_37_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12752" *) _1272_;
  assign FpAdd_8U_23U_is_inf_1_lpi_1_dfm_2_mx0w0 = nor_33_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12753" *) _1273_;
  assign FpAdd_8U_23U_is_inf_lpi_1_dfm_2_mx0w0 = nor_45_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12754" *) _1274_;
  assign _1310_ = IsNaN_8U_23U_3_nor_10_tmp | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12759" *) _1156_;
  assign _1304_ = IsNaN_8U_23U_3_nor_8_tmp | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12760" *) _1157_;
  assign _1308_ = IsNaN_8U_23U_3_nor_6_tmp | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12761" *) _1158_;
  assign _1306_ = IsNaN_8U_23U_3_nor_4_tmp | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12762" *) _1159_;
  assign _1587_ = FpAlu_8U_23U_equal_tmp_mx0w0 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12767" *) FpAlu_8U_23U_equal_tmp_1_mx0w0;
  assign _1588_ = _1587_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12767" *) FpAlu_8U_23U_equal_tmp_2_mx0w0;
  assign _1589_ = IsNaN_8U_23U_2_nor_2_mx0w0 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12810" *) IsNaN_8U_23U_4_IsNaN_8U_23U_4_nand_2_itm_mx0w2;
  assign _1590_ = _1275_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12812" *) _1161_;
  assign _1591_ = _1276_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12814" *) _1163_;
  assign _1592_ = IsNaN_8U_23U_2_nor_3_mx0w0 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12816" *) IsNaN_8U_23U_4_IsNaN_8U_23U_4_nand_3_itm_mx0w2;
  assign _1593_ = FpAlu_8U_23U_equal_tmp_2_mx0w0 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12818" *) FpAlu_8U_23U_equal_tmp_1_mx0w0;
  assign _1594_ = _1593_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12818" *) alu_loop_op_else_equal_tmp_2;
  assign FpCmp_8U_23U_false_is_abs_a_greater_2_lpi_1_dfm_1_mx0w0 = _0547_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12823" *) FpCmp_8U_23U_true_if_acc_6_nl[8];
  assign _1595_ = FpAdd_8U_23U_int_mant_1_lpi_1_dfm_2_mx0[0] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12883" *) FpAdd_8U_23U_int_mant_1_lpi_1_dfm_2_mx0[1];
  assign _1596_ = _1595_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12883" *) FpAdd_8U_23U_int_mant_1_lpi_1_dfm_2_mx0[2];
  assign _1597_ = _1596_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12884" *) FpAdd_8U_23U_int_mant_1_lpi_1_dfm_2_mx0[3];
  assign _1598_ = _1597_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12884" *) FpAdd_8U_23U_int_mant_1_lpi_1_dfm_2_mx0[4];
  assign _1599_ = _1598_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12885" *) FpAdd_8U_23U_int_mant_1_lpi_1_dfm_2_mx0[5];
  assign _1600_ = _1599_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12885" *) FpAdd_8U_23U_int_mant_1_lpi_1_dfm_2_mx0[6];
  assign _1601_ = _1600_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12886" *) FpAdd_8U_23U_int_mant_1_lpi_1_dfm_2_mx0[7];
  assign _1602_ = _1601_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12886" *) FpAdd_8U_23U_int_mant_1_lpi_1_dfm_2_mx0[8];
  assign _1603_ = _1602_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12887" *) FpAdd_8U_23U_int_mant_1_lpi_1_dfm_2_mx0[9];
  assign _1604_ = _1603_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12887" *) FpAdd_8U_23U_int_mant_1_lpi_1_dfm_2_mx0[10];
  assign _1605_ = _1604_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12888" *) FpAdd_8U_23U_int_mant_1_lpi_1_dfm_2_mx0[11];
  assign _1606_ = _1605_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12888" *) FpAdd_8U_23U_int_mant_1_lpi_1_dfm_2_mx0[12];
  assign _1607_ = _1606_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12889" *) FpAdd_8U_23U_int_mant_1_lpi_1_dfm_2_mx0[13];
  assign _1608_ = _1607_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12889" *) FpAdd_8U_23U_int_mant_1_lpi_1_dfm_2_mx0[14];
  assign _1609_ = _1608_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12890" *) FpAdd_8U_23U_int_mant_1_lpi_1_dfm_2_mx0[15];
  assign _1610_ = _1609_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12890" *) FpAdd_8U_23U_int_mant_1_lpi_1_dfm_2_mx0[16];
  assign _1611_ = _1610_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12891" *) FpAdd_8U_23U_int_mant_1_lpi_1_dfm_2_mx0[17];
  assign _1612_ = _1611_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12891" *) FpAdd_8U_23U_int_mant_1_lpi_1_dfm_2_mx0[18];
  assign _1613_ = _1612_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12892" *) FpAdd_8U_23U_int_mant_1_lpi_1_dfm_2_mx0[19];
  assign _1614_ = _1613_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12892" *) FpAdd_8U_23U_int_mant_1_lpi_1_dfm_2_mx0[20];
  assign _1615_ = _1614_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12893" *) FpAdd_8U_23U_int_mant_1_lpi_1_dfm_2_mx0[21];
  assign _1616_ = _1615_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12893" *) FpAdd_8U_23U_int_mant_1_lpi_1_dfm_2_mx0[22];
  assign _1617_ = _1616_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12894" *) FpAdd_8U_23U_int_mant_1_lpi_1_dfm_2_mx0[23];
  assign _1618_ = _1617_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12894" *) FpAdd_8U_23U_int_mant_1_lpi_1_dfm_2_mx0[25];
  assign _1619_ = FpAdd_8U_23U_int_mant_4_lpi_1_dfm_2_mx0[0] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12903" *) FpAdd_8U_23U_int_mant_4_lpi_1_dfm_2_mx0[1];
  assign _1620_ = _1619_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12903" *) FpAdd_8U_23U_int_mant_4_lpi_1_dfm_2_mx0[2];
  assign _1621_ = _1620_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12904" *) FpAdd_8U_23U_int_mant_4_lpi_1_dfm_2_mx0[3];
  assign _1622_ = _1621_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12904" *) FpAdd_8U_23U_int_mant_4_lpi_1_dfm_2_mx0[4];
  assign _1623_ = _1622_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12905" *) FpAdd_8U_23U_int_mant_4_lpi_1_dfm_2_mx0[5];
  assign _1624_ = _1623_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12905" *) FpAdd_8U_23U_int_mant_4_lpi_1_dfm_2_mx0[6];
  assign _1625_ = _1624_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12906" *) FpAdd_8U_23U_int_mant_4_lpi_1_dfm_2_mx0[7];
  assign _1626_ = _1625_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12906" *) FpAdd_8U_23U_int_mant_4_lpi_1_dfm_2_mx0[8];
  assign _1627_ = _1626_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12907" *) FpAdd_8U_23U_int_mant_4_lpi_1_dfm_2_mx0[9];
  assign _1628_ = _1627_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12907" *) FpAdd_8U_23U_int_mant_4_lpi_1_dfm_2_mx0[10];
  assign _1629_ = _1628_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12908" *) FpAdd_8U_23U_int_mant_4_lpi_1_dfm_2_mx0[11];
  assign _1630_ = _1629_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12908" *) FpAdd_8U_23U_int_mant_4_lpi_1_dfm_2_mx0[12];
  assign _1631_ = _1630_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12909" *) FpAdd_8U_23U_int_mant_4_lpi_1_dfm_2_mx0[13];
  assign _1632_ = _1631_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12909" *) FpAdd_8U_23U_int_mant_4_lpi_1_dfm_2_mx0[14];
  assign _1633_ = _1632_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12910" *) FpAdd_8U_23U_int_mant_4_lpi_1_dfm_2_mx0[15];
  assign _1634_ = _1633_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12910" *) FpAdd_8U_23U_int_mant_4_lpi_1_dfm_2_mx0[16];
  assign _1635_ = _1634_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12911" *) FpAdd_8U_23U_int_mant_4_lpi_1_dfm_2_mx0[17];
  assign _1636_ = _1635_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12911" *) FpAdd_8U_23U_int_mant_4_lpi_1_dfm_2_mx0[18];
  assign _1637_ = _1636_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12912" *) FpAdd_8U_23U_int_mant_4_lpi_1_dfm_2_mx0[19];
  assign _1638_ = _1637_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12912" *) FpAdd_8U_23U_int_mant_4_lpi_1_dfm_2_mx0[20];
  assign _1639_ = _1638_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12913" *) FpAdd_8U_23U_int_mant_4_lpi_1_dfm_2_mx0[21];
  assign _1640_ = _1639_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12913" *) FpAdd_8U_23U_int_mant_4_lpi_1_dfm_2_mx0[22];
  assign _1641_ = _1640_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12914" *) FpAdd_8U_23U_int_mant_4_lpi_1_dfm_2_mx0[23];
  assign _1642_ = _1641_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12914" *) FpAdd_8U_23U_int_mant_4_lpi_1_dfm_2_mx0[25];
  assign _1643_ = FpAdd_8U_23U_int_mant_3_lpi_1_dfm_2_mx0[0] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12923" *) FpAdd_8U_23U_int_mant_3_lpi_1_dfm_2_mx0[1];
  assign _1644_ = _1643_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12923" *) FpAdd_8U_23U_int_mant_3_lpi_1_dfm_2_mx0[2];
  assign _1645_ = _1644_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12924" *) FpAdd_8U_23U_int_mant_3_lpi_1_dfm_2_mx0[3];
  assign _1646_ = _1645_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12924" *) FpAdd_8U_23U_int_mant_3_lpi_1_dfm_2_mx0[4];
  assign _1647_ = _1646_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12925" *) FpAdd_8U_23U_int_mant_3_lpi_1_dfm_2_mx0[5];
  assign _1648_ = _1647_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12925" *) FpAdd_8U_23U_int_mant_3_lpi_1_dfm_2_mx0[6];
  assign _1649_ = _1648_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12926" *) FpAdd_8U_23U_int_mant_3_lpi_1_dfm_2_mx0[7];
  assign _1650_ = _1649_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12926" *) FpAdd_8U_23U_int_mant_3_lpi_1_dfm_2_mx0[8];
  assign _1651_ = _1650_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12927" *) FpAdd_8U_23U_int_mant_3_lpi_1_dfm_2_mx0[9];
  assign _1652_ = _1651_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12927" *) FpAdd_8U_23U_int_mant_3_lpi_1_dfm_2_mx0[10];
  assign _1653_ = _1652_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12928" *) FpAdd_8U_23U_int_mant_3_lpi_1_dfm_2_mx0[11];
  assign _1654_ = _1653_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12928" *) FpAdd_8U_23U_int_mant_3_lpi_1_dfm_2_mx0[12];
  assign _1655_ = _1654_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12929" *) FpAdd_8U_23U_int_mant_3_lpi_1_dfm_2_mx0[13];
  assign _1656_ = _1655_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12929" *) FpAdd_8U_23U_int_mant_3_lpi_1_dfm_2_mx0[14];
  assign _1657_ = _1656_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12930" *) FpAdd_8U_23U_int_mant_3_lpi_1_dfm_2_mx0[15];
  assign _1658_ = _1657_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12930" *) FpAdd_8U_23U_int_mant_3_lpi_1_dfm_2_mx0[16];
  assign _1659_ = _1658_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12931" *) FpAdd_8U_23U_int_mant_3_lpi_1_dfm_2_mx0[17];
  assign _1660_ = _1659_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12931" *) FpAdd_8U_23U_int_mant_3_lpi_1_dfm_2_mx0[18];
  assign _1661_ = _1660_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12932" *) FpAdd_8U_23U_int_mant_3_lpi_1_dfm_2_mx0[19];
  assign _1662_ = _1661_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12932" *) FpAdd_8U_23U_int_mant_3_lpi_1_dfm_2_mx0[20];
  assign _1663_ = _1662_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12933" *) FpAdd_8U_23U_int_mant_3_lpi_1_dfm_2_mx0[21];
  assign _1664_ = _1663_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12933" *) FpAdd_8U_23U_int_mant_3_lpi_1_dfm_2_mx0[22];
  assign _1665_ = _1664_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12934" *) FpAdd_8U_23U_int_mant_3_lpi_1_dfm_2_mx0[23];
  assign _1666_ = _1665_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12934" *) FpAdd_8U_23U_int_mant_3_lpi_1_dfm_2_mx0[25];
  assign _1667_ = FpAdd_8U_23U_int_mant_2_lpi_1_dfm_2_mx0[0] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12943" *) FpAdd_8U_23U_int_mant_2_lpi_1_dfm_2_mx0[1];
  assign _1668_ = _1667_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12943" *) FpAdd_8U_23U_int_mant_2_lpi_1_dfm_2_mx0[2];
  assign _1669_ = _1668_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12944" *) FpAdd_8U_23U_int_mant_2_lpi_1_dfm_2_mx0[3];
  assign _1670_ = _1669_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12944" *) FpAdd_8U_23U_int_mant_2_lpi_1_dfm_2_mx0[4];
  assign _1671_ = _1670_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12945" *) FpAdd_8U_23U_int_mant_2_lpi_1_dfm_2_mx0[5];
  assign _1672_ = _1671_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12945" *) FpAdd_8U_23U_int_mant_2_lpi_1_dfm_2_mx0[6];
  assign _1673_ = _1672_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12946" *) FpAdd_8U_23U_int_mant_2_lpi_1_dfm_2_mx0[7];
  assign _1674_ = _1673_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12946" *) FpAdd_8U_23U_int_mant_2_lpi_1_dfm_2_mx0[8];
  assign _1675_ = _1674_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12947" *) FpAdd_8U_23U_int_mant_2_lpi_1_dfm_2_mx0[9];
  assign _1676_ = _1675_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12947" *) FpAdd_8U_23U_int_mant_2_lpi_1_dfm_2_mx0[10];
  assign _1677_ = _1676_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12948" *) FpAdd_8U_23U_int_mant_2_lpi_1_dfm_2_mx0[11];
  assign _1678_ = _1677_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12948" *) FpAdd_8U_23U_int_mant_2_lpi_1_dfm_2_mx0[12];
  assign _1679_ = _1678_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12949" *) FpAdd_8U_23U_int_mant_2_lpi_1_dfm_2_mx0[13];
  assign _1680_ = _1679_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12949" *) FpAdd_8U_23U_int_mant_2_lpi_1_dfm_2_mx0[14];
  assign _1681_ = _1680_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12950" *) FpAdd_8U_23U_int_mant_2_lpi_1_dfm_2_mx0[15];
  assign _1682_ = _1681_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12950" *) FpAdd_8U_23U_int_mant_2_lpi_1_dfm_2_mx0[16];
  assign _1683_ = _1682_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12951" *) FpAdd_8U_23U_int_mant_2_lpi_1_dfm_2_mx0[17];
  assign _1684_ = _1683_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12951" *) FpAdd_8U_23U_int_mant_2_lpi_1_dfm_2_mx0[18];
  assign _1685_ = _1684_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12952" *) FpAdd_8U_23U_int_mant_2_lpi_1_dfm_2_mx0[19];
  assign _1686_ = _1685_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12952" *) FpAdd_8U_23U_int_mant_2_lpi_1_dfm_2_mx0[20];
  assign _1687_ = _1686_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12953" *) FpAdd_8U_23U_int_mant_2_lpi_1_dfm_2_mx0[21];
  assign _1688_ = _1687_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12953" *) FpAdd_8U_23U_int_mant_2_lpi_1_dfm_2_mx0[22];
  assign _1689_ = _1688_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12954" *) FpAdd_8U_23U_int_mant_2_lpi_1_dfm_2_mx0[23];
  assign _1690_ = _1689_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12954" *) FpAdd_8U_23U_int_mant_2_lpi_1_dfm_2_mx0[25];
  assign _1691_ = FpAdd_8U_23U_and_3_tmp_3 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12973" *) FpAdd_8U_23U_is_inf_lpi_1_dfm_8;
  assign or_962_nl = IsNaN_8U_23U_1_land_lpi_1_dfm_9 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12993" *) IsNaN_8U_23U_land_lpi_1_dfm_11;
  assign _1692_ = IsNaN_8U_23U_1_land_3_lpi_1_dfm_9 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12995" *) IsNaN_8U_23U_land_3_lpi_1_dfm_11;
  assign _1693_ = IsNaN_8U_23U_1_land_2_lpi_1_dfm_9 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12997" *) IsNaN_8U_23U_land_2_lpi_1_dfm_11;
  assign _1694_ = IsNaN_8U_23U_1_land_1_lpi_1_dfm_9 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12999" *) IsNaN_8U_23U_land_1_lpi_1_dfm_11;
  assign _1695_ = chn_alu_op_rsci_bawt | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13006" *) _1283_;
  assign _1696_ = cfg_alu_algo_rsc_triosy_obj_bawt | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13007" *) _1192_;
  assign _1697_ = cfg_alu_op_rsc_triosy_obj_bawt | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13007" *) _1192_;
  assign _1698_ = cfg_alu_src_rsc_triosy_obj_bawt | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13008" *) _1192_;
  assign _1699_ = cfg_alu_bypass_rsc_triosy_obj_bawt | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13009" *) _1192_;
  assign _1700_ = alu_loop_op_2_IntSaturation_33U_32U_else_if_acc_1_nl[2] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13075" *) alu_loop_op_2_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_1_svs_3;
  assign _1701_ = alu_loop_op_4_IntSaturation_33U_32U_else_if_acc_1_nl[2] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13082" *) alu_loop_op_4_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_1_svs_2;
  assign _1702_ = alu_loop_op_3_IntSaturation_33U_32U_else_if_acc_nl[2] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13089" *) alu_loop_op_3_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_svs_2;
  assign _1703_ = alu_loop_op_1_IntSaturation_33U_32U_else_if_acc_nl[2] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13096" *) alu_loop_op_1_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_svs_2;
  assign _1704_ = FpCmp_8U_23U_false_else_if_acc_4_nl[8] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13125" *) _1288_;
  assign or_861_cse = _1289_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13125" *) FpCmp_8U_23U_true_if_acc_4_nl[8];
  assign _1705_ = AluIn_data_sva_127[31] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13126" *) _1290_;
  assign _1706_ = mux_339_nl | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13129" *) IsNaN_8U_23U_2_IsNaN_8U_23U_2_nor_itm_2;
  assign _1707_ = FpCmp_8U_23U_false_else_if_acc_6_nl[8] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13132" *) _1291_;
  assign or_864_nl = _1292_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13133" *) FpCmp_8U_23U_true_if_acc_6_nl[8];
  assign _1708_ = _0560_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13137" *) mux_340_nl;
  assign _1709_ = _1293_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13137" *) IsNaN_8U_23U_2_IsNaN_8U_23U_2_nor_1_itm_1;
  assign _1710_ = _1294_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13147" *) FpCmp_8U_23U_false_else_if_acc_8_nl[8];
  assign or_867_cse = _1295_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13147" *) FpCmp_8U_23U_true_if_acc_8_nl[8];
  assign _1711_ = AluIn_data_sva_127[95] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13148" *) _1296_;
  assign _1712_ = mux_341_nl | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13151" *) IsNaN_8U_23U_2_IsNaN_8U_23U_2_nor_2_itm_1;
  assign _1713_ = _1297_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13161" *) FpCmp_8U_23U_false_else_if_acc_10_nl[8];
  assign or_871_cse = _1298_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13161" *) FpCmp_8U_23U_true_if_acc_10_nl[8];
  assign _1714_ = AluIn_data_sva_127[127] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13162" *) _1299_;
  assign _1715_ = mux_342_nl | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13165" *) IsNaN_8U_23U_2_IsNaN_8U_23U_2_nor_3_itm_2;
  assign _1716_ = else_mux_tmp_31_23[8] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13169" *) _1290_;
  assign or_876_nl = mux_343_nl | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13171" *) IsNaN_8U_23U_2_IsNaN_8U_23U_2_nor_3_itm_2;
  assign _1717_ = else_mux_2_tmp_31_23[8] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13175" *) _1296_;
  assign _1718_ = IsNaN_8U_23U_2_IsNaN_8U_23U_2_nor_1_itm_1 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13178" *) IsNaN_8U_23U_4_nor_2_itm_2;
  assign or_880_nl = mux_344_nl | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13178" *) _1300_;
  assign _1719_ = else_mux_3_tmp_31_23[8] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13182" *) _1299_;
  assign _1720_ = IsNaN_8U_23U_2_IsNaN_8U_23U_2_nor_2_itm_1 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13185" *) IsNaN_8U_23U_4_nor_3_itm_3;
  assign or_884_nl = mux_345_nl | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13185" *) _1301_;
  assign FpCmp_8U_23U_false_if_1_FpCmp_8U_23U_false_if_1_or_1_nl = FpCmp_8U_23U_false_is_abs_a_greater_2_lpi_1_dfm_1_mx0 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13191" *) else_AluOp_data_1_lpi_1_dfm_mx0[31];
  assign _1721_ = FpCmp_8U_23U_false_mux_4_nl | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13194" *) IsNaN_8U_23U_1_land_2_lpi_1_dfm_mx0w0;
  assign _1722_ = _1485_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13271" *) _1167_;
  assign _1723_ = _1722_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13271" *) or_dcpl_154;
  assign or_tmp_9 = _1723_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13271" *) and_tmp;
  assign _1724_ = _1167_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13274" *) or_dcpl_154;
  assign or_967_nl = _1315_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13275" *) and_tmp;
  assign or_tmp_15 = _1722_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13279" *) and_tmp;
  assign or_965_nl = _1316_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13280" *) and_tmp;
  assign or_tmp_20 = _1485_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13283" *) and_tmp;
  assign _1725_ = nor_269_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13291" *) cfg_alu_bypass_rsci_d;
  assign or_tmp_23 = _1725_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13291" *) not_tmp_24;
  assign _1726_ = _1485_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13293" *) cfg_alu_algo_1_sva_st_22[0];
  assign _1727_ = _1726_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13295" *) _1318_;
  assign _1728_ = _1487_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13297" *) or_dcpl_86;
  assign _1729_ = or_1087_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13300" *) _1194_;
  assign _1730_ = _1148_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13302" *) io_read_cfg_alu_bypass_rsc_svs_st_6;
  assign or_tmp_75 = _1730_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13302" *) _1203_;
  assign _1731_ = or_1087_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13304" *) _1148_;
  assign _1732_ = _1731_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13304" *) io_read_cfg_alu_bypass_rsc_svs_st_6;
  assign _1733_ = _1732_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13305" *) _1203_;
  assign or_87_nl = or_dcpl_86 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13307" *) io_read_cfg_alu_bypass_rsc_svs_st_5;
  assign _1734_ = io_read_cfg_alu_bypass_rsc_svs_st_7 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13312" *) alu_loop_op_unequal_tmp_8;
  assign _1735_ = _1734_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13312" *) io_read_cfg_alu_bypass_rsc_svs_8;
  assign or_tmp_218 = _1735_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13312" *) _1206_;
  assign _1736_ = nor_269_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13313" *) FpAlu_8U_23U_equal_tmp_22;
  assign _1737_ = _1736_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13314" *) alu_loop_op_unequal_tmp_7;
  assign _1738_ = _1737_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13314" *) io_read_cfg_alu_bypass_rsc_svs_7;
  assign _1739_ = _1738_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13314" *) io_read_cfg_alu_bypass_rsc_svs_st_6;
  assign or_230_nl = _1739_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13315" *) _1203_;
  assign _1740_ = FpAlu_8U_23U_equal_tmp_22 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13316" *) alu_loop_op_unequal_tmp_7;
  assign _1741_ = _1740_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13317" *) io_read_cfg_alu_bypass_rsc_svs_7;
  assign _1742_ = _1741_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13317" *) io_read_cfg_alu_bypass_rsc_svs_st_6;
  assign or_233_nl = _1742_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13317" *) _1203_;
  assign or_tmp_224 = io_read_cfg_alu_bypass_rsc_svs_st_7 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13320" *) _1206_;
  assign _1743_ = alu_loop_op_unequal_tmp_7 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13322" *) io_read_cfg_alu_bypass_rsc_svs_7;
  assign or_tmp_251 = _1743_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13322" *) _1203_;
  assign _1744_ = _1319_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13324" *) _1242_;
  assign _1745_ = _1744_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13324" *) alu_loop_op_unequal_tmp_7;
  assign _1746_ = _1745_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13324" *) io_read_cfg_alu_bypass_rsc_svs_7;
  assign or_tmp_261 = _1746_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13324" *) _1203_;
  assign _1747_ = _1242_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13325" *) alu_loop_op_unequal_tmp_7;
  assign _1748_ = _1747_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13326" *) io_read_cfg_alu_bypass_rsc_svs_7;
  assign or_tmp_269 = _1748_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13326" *) _1203_;
  assign _1749_ = _1743_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13328" *) io_read_cfg_alu_bypass_rsc_svs_st_6;
  assign or_tmp_280 = _1749_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13328" *) _1203_;
  assign _1750_ = _1320_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13330" *) _1319_;
  assign _1751_ = _1750_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13330" *) _1242_;
  assign _1752_ = _1751_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13330" *) alu_loop_op_unequal_tmp_7;
  assign _1753_ = _1752_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13331" *) io_read_cfg_alu_bypass_rsc_svs_7;
  assign _1754_ = _1753_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13331" *) io_read_cfg_alu_bypass_rsc_svs_st_6;
  assign or_tmp_293 = _1754_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13331" *) _1203_;
  assign _1755_ = _1321_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13333" *) io_read_cfg_alu_bypass_rsc_svs_7;
  assign or_tmp_305 = _1755_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13333" *) _1203_;
  assign _1756_ = _1322_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13335" *) io_read_cfg_alu_bypass_rsc_svs_8;
  assign or_tmp_309 = _1756_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13335" *) _1206_;
  assign _1757_ = _1196_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13341" *) io_read_cfg_alu_bypass_rsc_svs_7;
  assign or_tmp_312 = _1757_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13341" *) _1203_;
  assign or_tmp_315 = or_239_nl | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13343" *) or_1050_cse;
  assign _1758_ = nor_269_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13344" *) _1194_;
  assign or_tmp_347 = _1758_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13344" *) or_1050_cse;
  assign or_386_nl = io_read_cfg_alu_bypass_rsc_svs_st_1 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13346" *) or_632_cse;
  assign _1759_ = io_read_cfg_alu_bypass_rsc_svs_st_1 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13347" *) not_tmp_152;
  assign or_383_nl = or_16_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13350" *) or_632_cse;
  assign _1760_ = or_16_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13354" *) not_tmp_152;
  assign or_417_nl = io_read_cfg_alu_bypass_rsc_svs_7 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13363" *) _1203_;
  assign _1761_ = io_read_cfg_alu_bypass_rsc_svs_7 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13365" *) io_read_cfg_alu_bypass_rsc_svs_st_6;
  assign or_419_nl = _1761_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13365" *) _1203_;
  assign or_tmp_402 = alu_loop_op_unequal_tmp_6 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13369" *) FpAlu_8U_23U_equal_tmp_21;
  assign _1762_ = or_1087_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13371" *) alu_loop_op_unequal_tmp_7;
  assign _1763_ = _1762_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13371" *) io_read_cfg_alu_bypass_rsc_svs_7;
  assign or_428_nl = _1763_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13371" *) _1203_;
  assign or_tmp_409 = alu_loop_op_unequal_tmp_6 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13374" *) io_read_cfg_alu_bypass_rsc_svs_st_5;
  assign _1764_ = _1763_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13377" *) io_read_cfg_alu_bypass_rsc_svs_st_6;
  assign or_432_nl = _1764_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13377" *) _1203_;
  assign _1765_ = nor_269_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13380" *) io_read_cfg_alu_bypass_rsc_svs_6;
  assign or_tmp_416 = _1765_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13380" *) _1194_;
  assign _1766_ = or_tmp_395 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13388" *) _1237_;
  assign _1767_ = or_1087_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13391" *) io_read_cfg_alu_bypass_rsc_svs_6;
  assign or_tmp_577 = _1767_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13391" *) _1194_;
  assign _1768_ = cfg_alu_algo_1_sva_st_22[0] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13394" *) _1183_;
  assign or_tmp_583 = _1768_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13394" *) chn_alu_out_rsci_bawt;
  assign _1769_ = _0008_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13396" *) _1183_;
  assign or_tmp_585 = _1769_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13396" *) chn_alu_out_rsci_bawt;
  assign or_612_nl = io_read_cfg_alu_bypass_rsc_svs_5 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13400" *) cfg_alu_algo_1_sva_2[1];
  assign or_609_nl = or_612_nl | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13400" *) mux_251_nl;
  assign _1770_ = io_read_cfg_alu_bypass_rsc_svs_5 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13403" *) _1183_;
  assign or_601_nl = _1770_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13403" *) chn_alu_out_rsci_bawt;
  assign or_607_nl = or_612_nl | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13408" *) mux_249_nl;
  assign _1771_ = _0009_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13414" *) _1183_;
  assign or_610_nl = _1771_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13414" *) chn_alu_out_rsci_bawt;
  assign _1772_ = nor_71_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13425" *) cfg_alu_algo_1_sva_st[1];
  assign or_tmp_596 = _1772_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13425" *) not_tmp_259;
  assign or_tmp_597 = cfg_alu_algo_1_sva_st[1] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13426" *) not_tmp_259;
  assign _1773_ = or_dcpl_154 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13427" *) _1325_;
  assign _1774_ = _0012_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13429" *) _1147_;
  assign or_629_nl = _1774_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13429" *) or_400_nl;
  assign _1775_ = io_read_cfg_alu_bypass_rsc_svs_5 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13436" *) or_dcpl_154;
  assign _1776_ = _1775_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13436" *) _1168_;
  assign _1777_ = _1776_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13436" *) or_1055_cse;
  assign _1778_ = _1775_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13439" *) or_1055_cse;
  assign _1779_ = chn_alu_op_rsci_bawt | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13449" *) io_read_cfg_alu_bypass_rsc_svs_st_1;
  assign _1780_ = or_dcpl_20 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13456" *) and_dcpl_34;
  assign or_dcpl_23 = and_dcpl_32 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13459" *) _1206_;
  assign or_dcpl_46 = or_1050_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13468" *) and_dcpl_32;
  assign or_dcpl_49 = and_dcpl_35 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13469" *) and_dcpl_32;
  assign or_tmp_657 = nor_269_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13479" *) io_read_cfg_alu_bypass_rsc_svs_7;
  assign _1781_ = or_1050_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13484" *) _1203_;
  assign _1782_ = _1781_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13485" *) io_read_cfg_alu_bypass_rsc_svs_st_6;
  assign _1783_ = _1782_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13485" *) _1148_;
  assign or_dcpl_85 = _1783_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13485" *) and_dcpl_32;
  assign _1784_ = or_dcpl_46 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13487" *) _1194_;
  assign _1785_ = _1784_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13488" *) io_read_cfg_alu_bypass_rsc_svs_st_5;
  assign or_dcpl_89 = _1785_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13488" *) or_dcpl_86;
  assign or_dcpl_91 = or_1050_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13489" *) _1194_;
  assign _1786_ = or_dcpl_20 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13490" *) and_dcpl_32;
  assign _1787_ = _1786_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13490" *) or_1050_cse;
  assign _1788_ = _1787_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13491" *) cfg_alu_algo_1_sva_st_22[0];
  assign _1789_ = _1788_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13491" *) and_dcpl_33;
  assign _1790_ = _1789_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13491" *) _0011_;
  assign _1791_ = _1790_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13492" *) io_read_cfg_alu_bypass_rsc_svs_st_1;
  assign or_dcpl_100 = _1791_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13492" *) _1192_;
  assign _1792_ = and_dcpl_35 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13493" *) or_tmp_386;
  assign _1793_ = _1792_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13493" *) _1332_;
  assign _1794_ = _1793_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13494" *) and_dcpl_32;
  assign or_dcpl_109 = _1794_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13494" *) cfg_precision[0];
  assign or_dcpl_117 = _1333_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13496" *) FpAdd_8U_23U_is_a_greater_oif_aelse_acc_nl[23];
  assign or_dcpl_119 = _1334_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13498" *) FpAdd_8U_23U_is_a_greater_oif_aelse_acc_1_nl[23];
  assign or_dcpl_121 = _1335_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13500" *) FpAdd_8U_23U_is_a_greater_oif_aelse_acc_2_nl[23];
  assign or_dcpl_123 = _1336_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13502" *) FpAdd_8U_23U_is_a_greater_oif_aelse_acc_3_nl[23];
  assign or_dcpl_125 = io_read_cfg_alu_bypass_rsc_svs_st_5 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13509" *) _1339_;
  assign _1795_ = cfg_precision[0] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13512" *) or_632_cse;
  assign _1796_ = _1795_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13512" *) io_read_cfg_alu_bypass_rsc_svs_st_1;
  assign _1797_ = or_1050_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13516" *) io_read_cfg_alu_bypass_rsc_svs_st_1;
  assign _1257_ = io_read_cfg_alu_bypass_rsc_svs_st_1 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13518" *) and_dcpl_77;
  assign or_tmp_668 = IsNaN_8U_23U_3_nor_4_tmp | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13534" *) _1169_;
  assign or_tmp_674 = IsNaN_8U_23U_3_nor_8_tmp | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13535" *) _1170_;
  assign or_tmp_678 = IsNaN_8U_23U_3_nor_10_tmp | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13536" *) _1171_;
  assign chn_alu_in_rsci_ld_core_psct_mx0c0 = main_stage_en_1 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13540" *) fsm_output[0];
  assign _1798_ = or_tmp_386 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13543" *) _1342_;
  assign cfg_alu_src_1_sva_st_1_mx0c1 = _0611_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13547" *) _0613_;
  assign _1799_ = _1780_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13548" *) _1192_;
  assign or_996_tmp = _0626_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13584" *) io_read_cfg_alu_bypass_rsc_svs_8;
  assign or_997_tmp = _0627_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13586" *) io_read_cfg_alu_bypass_rsc_svs_8;
  assign or_998_tmp = _0629_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13588" *) io_read_cfg_alu_bypass_rsc_svs_8;
  assign _1800_ = _1343_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13596" *) FpCmp_8U_23U_true_if_acc_10_nl[8];
  assign _1801_ = _1345_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13598" *) FpCmp_8U_23U_true_if_acc_8_nl[8];
  assign _1802_ = _1347_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13600" *) FpCmp_8U_23U_true_if_acc_6_nl[8];
  assign _1803_ = _1349_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13602" *) FpCmp_8U_23U_true_if_acc_4_nl[8];
  assign or_dcpl = _0625_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13610" *) io_read_cfg_alu_bypass_rsc_svs_8;
  assign _1804_ = and_dcpl_43 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13720" *) and_dcpl_45;
  assign _1805_ = and_357_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13729" *) _0636_;
  assign _1806_ = _1805_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13729" *) chn_alu_op_rsci_ld_core_psct_mx0c1;
  assign _1807_ = or_tmp_695 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13737" *) main_stage_v_1_mx0c1;
  assign _1808_ = and_dcpl_83 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13788" *) and_167_rgt;
  assign _1809_ = _0644_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13799" *) _0635_;
  assign _1810_ = _1809_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13799" *) cfg_alu_src_1_sva_st_1_mx0c1;
  assign _1811_ = or_dcpl_49 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13809" *) _1188_;
  assign _1812_ = _1811_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13809" *) fsm_output[0];
  assign _1813_ = and_dcpl_64 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13817" *) main_stage_v_2_mx0c1;
  assign _1814_ = and_dcpl_96 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13960" *) main_stage_v_3_mx0c1;
  assign _1815_ = _0654_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14088" *) main_stage_v_4_mx0c1;
  assign _1816_ = _0667_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14184" *) io_read_cfg_alu_bypass_rsc_svs_7;
  assign _1817_ = and_564_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14192" *) _0670_;
  assign _1818_ = _0673_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14194" *) io_read_cfg_alu_bypass_rsc_svs_7;
  assign _1819_ = _0680_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14261" *) io_read_cfg_alu_bypass_rsc_svs_7;
  assign _1820_ = and_564_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14269" *) _0683_;
  assign _1821_ = _0686_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14271" *) io_read_cfg_alu_bypass_rsc_svs_7;
  assign _1822_ = _0689_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14280" *) io_read_cfg_alu_bypass_rsc_svs_7;
  assign _1823_ = and_564_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14288" *) _0692_;
  assign _1824_ = _0695_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14290" *) io_read_cfg_alu_bypass_rsc_svs_7;
  assign _1825_ = _0698_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14299" *) io_read_cfg_alu_bypass_rsc_svs_7;
  assign _1826_ = and_564_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14307" *) _0701_;
  assign _1827_ = _0704_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14309" *) io_read_cfg_alu_bypass_rsc_svs_7;
  assign _1828_ = mux_383_nl | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14345" *) io_read_cfg_alu_bypass_rsc_svs_8;
  assign _1829_ = _0707_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14346" *) nor_tmp_144;
  assign _1830_ = _0711_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14364" *) and_211_rgt;
  assign _1831_ = _0715_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14383" *) nor_tmp_144;
  assign _1832_ = _0718_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14403" *) and_213_rgt;
  assign _1833_ = _0722_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14421" *) and_215_rgt;
  assign _1834_ = FpAlu_8U_23U_equal_tmp_29 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14454" *) FpAlu_8U_23U_equal_tmp_23;
  assign _1835_ = _1834_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14455" *) FpAlu_8U_23U_equal_tmp_26;
  assign _1836_ = _1835_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14455" *) FpAlu_8U_23U_nor_dfs_6;
  assign _1837_ = _1369_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14455" *) alu_loop_op_unequal_tmp_8;
  assign _1838_ = _0733_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14483" *) and_217_rgt;
  assign _1839_ = or_dcpl_109 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14796" *) fsm_output[0];
  assign _1840_ = _1792_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14804" *) and_dcpl_32;
  assign _1841_ = _1840_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14804" *) fsm_output[0];
  assign _1842_ = and_231_rgt | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14821" *) and_233_rgt;
  assign _1843_ = _1842_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14821" *) and_dcpl_99;
  assign _1844_ = and_235_rgt | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14832" *) and_237_rgt;
  assign _1845_ = _1844_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14832" *) and_dcpl_99;
  assign _1846_ = and_239_rgt | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14843" *) and_241_rgt;
  assign _1847_ = _1846_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14843" *) and_dcpl_99;
  assign _1848_ = and_243_rgt | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14854" *) and_245_rgt;
  assign _1849_ = _1848_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14854" *) and_dcpl_99;
  assign _1850_ = or_dcpl_127 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15094" *) or_dcpl_125;
  assign _1851_ = _1850_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15095" *) cfg_alu_algo_1_sva_st_23[0];
  assign _1852_ = _1851_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15095" *) IsNaN_8U_23U_land_1_lpi_1_dfm_st_4;
  assign _1853_ = _1851_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15104" *) IsNaN_8U_23U_land_2_lpi_1_dfm_st_4;
  assign _1854_ = _1851_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15113" *) IsNaN_8U_23U_land_3_lpi_1_dfm_st_4;
  assign _1855_ = _1851_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15122" *) IsNaN_8U_23U_land_lpi_1_dfm_st_4;
  assign _1856_ = _0787_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15163" *) FpAdd_8U_23U_qr_2_lpi_1_dfm_mx0c1;
  assign _1857_ = _0790_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15173" *) FpAdd_8U_23U_qr_3_lpi_1_dfm_mx0c1;
  assign _1858_ = _0793_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15183" *) FpAdd_8U_23U_qr_4_lpi_1_dfm_mx0c1;
  assign _1859_ = _0796_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15193" *) FpAdd_8U_23U_qr_lpi_1_dfm_mx0c1;
  assign _1860_ = mux_363_nl | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15305" *) nor_202_cse;
  assign _1861_ = mux_364_nl | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15326" *) nor_202_cse;
  assign _1862_ = _0836_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15338" *) and_293_rgt;
  assign _1863_ = nor_269_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15372" *) alu_loop_op_4_IntSaturation_33U_32U_if_acc_1_nl[2];
  assign _1864_ = mux_366_nl | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15381" *) nor_202_cse;
  assign _1865_ = or_dcpl_20 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15473" *) or_dcpl_46;
  assign _1866_ = _1865_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15474" *) _1167_;
  assign _1867_ = _1866_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15474" *) and_dcpl_33;
  assign _1868_ = _1867_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15474" *) io_read_cfg_alu_bypass_rsc_svs_st_1;
  assign _1869_ = _1868_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15475" *) _1192_;
  assign _1870_ = _1869_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15475" *) or_dcpl_154;
  assign _1871_ = and_dcpl_239 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15534" *) and_328_rgt;
  assign _1872_ = FpAdd_8U_23U_and_tmp_2 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15566" *) FpAdd_8U_23U_is_inf_1_lpi_1_dfm_8;
  assign _1873_ = asn_267 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15582" *) or_996_tmp;
  assign _1874_ = FpAdd_8U_23U_and_1_tmp_3 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15586" *) FpAdd_8U_23U_is_inf_2_lpi_1_dfm_8;
  assign _1875_ = asn_267 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15602" *) or_997_tmp;
  assign or_43_nl = cfg_alu_bypass_rsci_d | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15617" *) not_tmp_24;
  assign _1876_ = io_read_cfg_alu_bypass_rsc_svs_st_1 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15625" *) _0015_;
  assign _1877_ = _1409_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15626" *) and_dcpl_32;
  assign _1878_ = acc_12_nl[50] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15627" *) _1194_;
  assign _1879_ = _1878_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15628" *) io_read_cfg_alu_bypass_rsc_svs_st_5;
  assign _1880_ = _1879_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15628" *) or_dcpl_86;
  assign _1881_ = alu_loop_op_1_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_itm | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15630" *) _1194_;
  assign _1882_ = _1881_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15630" *) io_read_cfg_alu_bypass_rsc_svs_st_5;
  assign _1883_ = _1882_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15630" *) or_dcpl_86;
  assign _1884_ = or_tmp_103 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15633" *) _1148_;
  assign _1885_ = _1884_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15633" *) alu_loop_op_1_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_itm_2;
  assign _1886_ = acc_13_nl[50] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15635" *) _1194_;
  assign _1887_ = _1886_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15636" *) io_read_cfg_alu_bypass_rsc_svs_st_5;
  assign _1888_ = _1887_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15636" *) or_dcpl_86;
  assign _1889_ = alu_loop_op_2_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_2_itm | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15638" *) _1194_;
  assign _1890_ = _1889_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15638" *) io_read_cfg_alu_bypass_rsc_svs_st_5;
  assign _1891_ = _1890_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15638" *) or_dcpl_86;
  assign _1892_ = _1884_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15641" *) alu_loop_op_2_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_2_itm_2;
  assign _1893_ = acc_14_nl[50] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15643" *) _1194_;
  assign _1894_ = _1893_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15644" *) io_read_cfg_alu_bypass_rsc_svs_st_5;
  assign _1895_ = _1894_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15644" *) or_dcpl_86;
  assign _1896_ = alu_loop_op_3_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_1_itm | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15646" *) _1194_;
  assign _1897_ = _1896_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15646" *) io_read_cfg_alu_bypass_rsc_svs_st_5;
  assign _1898_ = _1897_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15646" *) or_dcpl_86;
  assign _1899_ = _1884_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15649" *) alu_loop_op_3_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_1_itm_2;
  assign _1900_ = acc_15_nl[50] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15651" *) _1194_;
  assign _1901_ = _1900_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15652" *) io_read_cfg_alu_bypass_rsc_svs_st_5;
  assign _1902_ = _1901_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15652" *) or_dcpl_86;
  assign _1903_ = alu_loop_op_4_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_3_itm | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15654" *) _1194_;
  assign _1904_ = _1903_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15654" *) io_read_cfg_alu_bypass_rsc_svs_st_5;
  assign _1905_ = _1904_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15654" *) or_dcpl_86;
  assign _1906_ = _1884_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15657" *) alu_loop_op_4_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_3_itm_2;
  assign _1907_ = or_1087_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15660" *) io_read_cfg_alu_bypass_rsc_svs_st_6;
  assign _1908_ = _1907_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15660" *) _1203_;
  assign _1909_ = nor_33_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15663" *) io_read_cfg_alu_bypass_rsc_svs_st_6;
  assign _1910_ = _1909_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15664" *) _1148_;
  assign _1911_ = _1910_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15664" *) _1202_;
  assign _1912_ = _1911_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15664" *) FpAlu_8U_23U_equal_tmp_22;
  assign _1913_ = _1912_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15665" *) IsNaN_8U_23U_1_land_1_lpi_1_dfm_8;
  assign _1914_ = _1913_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15665" *) IsNaN_8U_23U_land_1_lpi_1_dfm_10;
  assign _1915_ = FpAdd_8U_23U_int_mant_p1_1_lpi_1_dfm_5[49] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15667" *) io_read_cfg_alu_bypass_rsc_svs_st_6;
  assign _1916_ = _1915_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15667" *) _1148_;
  assign _1917_ = _1916_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15667" *) _1202_;
  assign _1918_ = _1917_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15668" *) FpAlu_8U_23U_equal_tmp_22;
  assign _1919_ = _1918_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15668" *) IsNaN_8U_23U_1_land_1_lpi_1_dfm_8;
  assign _1920_ = _1919_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15668" *) IsNaN_8U_23U_land_1_lpi_1_dfm_10;
  assign _1921_ = _1219_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15670" *) alu_loop_op_1_FpAdd_8U_23U_if_4_if_acc_1_nl[7];
  assign _1922_ = _1730_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15673" *) _1202_;
  assign _1923_ = _1922_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15673" *) FpAlu_8U_23U_equal_tmp_22;
  assign _1924_ = _1923_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15674" *) IsNaN_8U_23U_1_land_1_lpi_1_dfm_8;
  assign _1925_ = _1924_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15674" *) IsNaN_8U_23U_land_1_lpi_1_dfm_10;
  assign _1926_ = alu_loop_op_unequal_tmp_7 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15677" *) mux_70_nl;
  assign _1927_ = or_417_nl | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15677" *) _1410_;
  assign _1928_ = _1411_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15680" *) _1412_;
  assign _1929_ = _1928_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15680" *) or_236_nl;
  assign _1930_ = _1929_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15680" *) IsNaN_8U_23U_1_land_1_lpi_1_dfm_9;
  assign _1931_ = _1930_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15681" *) IsNaN_8U_23U_land_1_lpi_1_dfm_11;
  assign _1932_ = _1931_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15681" *) _1205_;
  assign _1933_ = _1932_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15681" *) FpAlu_8U_23U_equal_tmp_23;
  assign _1934_ = _1933_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15682" *) io_read_cfg_alu_bypass_rsc_svs_st_7;
  assign _1935_ = _1934_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15682" *) FpAdd_8U_23U_is_inf_1_lpi_1_dfm_8;
  assign _1936_ = _1413_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15682" *) alu_loop_op_unequal_tmp_8;
  assign _1937_ = or_236_nl | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15684" *) IsNaN_8U_23U_1_land_1_lpi_1_dfm_9;
  assign _1938_ = _1937_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15684" *) IsNaN_8U_23U_land_1_lpi_1_dfm_11;
  assign _1939_ = _1938_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15684" *) _1205_;
  assign _1940_ = _1939_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15685" *) FpAlu_8U_23U_equal_tmp_23;
  assign _1941_ = _1940_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15685" *) io_read_cfg_alu_bypass_rsc_svs_st_7;
  assign _1942_ = _1941_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15685" *) FpAdd_8U_23U_is_inf_1_lpi_1_dfm_8;
  assign _1943_ = _1414_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15686" *) alu_loop_op_unequal_tmp_8;
  assign _1944_ = or_323_nl | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15688" *) mux_73_nl;
  assign _1945_ = nor_37_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15690" *) io_read_cfg_alu_bypass_rsc_svs_st_6;
  assign _1946_ = _1945_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15691" *) _1148_;
  assign _1947_ = _1946_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15691" *) _1202_;
  assign _1948_ = _1947_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15691" *) FpAlu_8U_23U_equal_tmp_22;
  assign _1949_ = _1948_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15692" *) IsNaN_8U_23U_1_land_2_lpi_1_dfm_8;
  assign _1950_ = _1949_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15692" *) IsNaN_8U_23U_land_2_lpi_1_dfm_10;
  assign _1951_ = FpAdd_8U_23U_int_mant_p1_2_lpi_1_dfm_5[49] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15694" *) io_read_cfg_alu_bypass_rsc_svs_st_6;
  assign _1952_ = _1951_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15694" *) _1148_;
  assign _1953_ = _1952_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15694" *) _1202_;
  assign _1954_ = _1953_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15695" *) FpAlu_8U_23U_equal_tmp_22;
  assign _1955_ = _1954_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15695" *) IsNaN_8U_23U_1_land_2_lpi_1_dfm_8;
  assign _1956_ = _1955_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15695" *) IsNaN_8U_23U_land_2_lpi_1_dfm_10;
  assign _1957_ = _1218_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15697" *) alu_loop_op_2_FpAdd_8U_23U_if_4_if_acc_4_nl[7];
  assign _1958_ = _1923_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15701" *) IsNaN_8U_23U_1_land_2_lpi_1_dfm_8;
  assign _1959_ = _1958_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15701" *) IsNaN_8U_23U_land_2_lpi_1_dfm_10;
  assign _1960_ = alu_loop_op_unequal_tmp_7 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15704" *) mux_76_nl;
  assign _1961_ = or_417_nl | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15704" *) _1415_;
  assign _1962_ = _1416_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15707" *) _1417_;
  assign _1963_ = _1962_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15707" *) or_236_nl;
  assign _1964_ = _1963_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15707" *) IsNaN_8U_23U_1_land_2_lpi_1_dfm_9;
  assign _1965_ = _1964_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15708" *) IsNaN_8U_23U_land_2_lpi_1_dfm_11;
  assign _1966_ = _1965_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15708" *) _1205_;
  assign _1967_ = _1966_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15708" *) FpAlu_8U_23U_equal_tmp_23;
  assign _1968_ = _1967_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15709" *) io_read_cfg_alu_bypass_rsc_svs_st_7;
  assign _1969_ = _1968_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15709" *) FpAdd_8U_23U_is_inf_2_lpi_1_dfm_8;
  assign _1970_ = _1418_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15709" *) alu_loop_op_unequal_tmp_8;
  assign _1971_ = or_236_nl | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15711" *) IsNaN_8U_23U_1_land_2_lpi_1_dfm_9;
  assign _1972_ = _1971_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15711" *) IsNaN_8U_23U_land_2_lpi_1_dfm_11;
  assign _1973_ = _1972_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15711" *) _1205_;
  assign _1974_ = _1973_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15712" *) FpAlu_8U_23U_equal_tmp_23;
  assign _1975_ = _1974_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15712" *) io_read_cfg_alu_bypass_rsc_svs_st_7;
  assign _1976_ = _1975_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15712" *) FpAdd_8U_23U_is_inf_2_lpi_1_dfm_8;
  assign _1977_ = _1419_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15713" *) alu_loop_op_unequal_tmp_8;
  assign _1978_ = or_323_nl | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15715" *) mux_79_nl;
  assign _1979_ = nor_41_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15717" *) io_read_cfg_alu_bypass_rsc_svs_st_6;
  assign _1980_ = _1979_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15718" *) _1148_;
  assign _1981_ = _1980_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15718" *) _1202_;
  assign _1982_ = _1981_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15718" *) FpAlu_8U_23U_equal_tmp_22;
  assign _1983_ = _1982_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15719" *) IsNaN_8U_23U_1_land_3_lpi_1_dfm_8;
  assign _1984_ = _1983_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15719" *) IsNaN_8U_23U_land_3_lpi_1_dfm_10;
  assign _1985_ = FpAdd_8U_23U_int_mant_p1_3_lpi_1_dfm_5[49] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15721" *) io_read_cfg_alu_bypass_rsc_svs_st_6;
  assign _1986_ = _1985_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15721" *) _1148_;
  assign _1987_ = _1986_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15721" *) _1202_;
  assign _1988_ = _1987_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15722" *) FpAlu_8U_23U_equal_tmp_22;
  assign _1989_ = _1988_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15722" *) IsNaN_8U_23U_1_land_3_lpi_1_dfm_8;
  assign _1990_ = _1989_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15722" *) IsNaN_8U_23U_land_3_lpi_1_dfm_10;
  assign _1991_ = _1215_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15724" *) alu_loop_op_3_FpAdd_8U_23U_if_4_if_acc_2_nl[7];
  assign _1992_ = _1923_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15728" *) IsNaN_8U_23U_1_land_3_lpi_1_dfm_8;
  assign _1993_ = _1992_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15728" *) IsNaN_8U_23U_land_3_lpi_1_dfm_10;
  assign _1994_ = alu_loop_op_unequal_tmp_7 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15731" *) mux_82_nl;
  assign _1995_ = or_417_nl | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15731" *) _1420_;
  assign _1996_ = _1421_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15734" *) _1422_;
  assign _1997_ = _1996_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15734" *) or_236_nl;
  assign _1998_ = _1997_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15734" *) IsNaN_8U_23U_1_land_3_lpi_1_dfm_9;
  assign _1999_ = _1998_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15735" *) IsNaN_8U_23U_land_3_lpi_1_dfm_11;
  assign _2000_ = _1999_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15735" *) _1205_;
  assign _2001_ = _2000_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15735" *) FpAlu_8U_23U_equal_tmp_23;
  assign _2002_ = _2001_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15736" *) io_read_cfg_alu_bypass_rsc_svs_st_7;
  assign _2003_ = _2002_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15736" *) FpAdd_8U_23U_is_inf_3_lpi_1_dfm_8;
  assign _2004_ = _1423_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15736" *) alu_loop_op_unequal_tmp_8;
  assign _2005_ = or_236_nl | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15738" *) IsNaN_8U_23U_1_land_3_lpi_1_dfm_9;
  assign _2006_ = _2005_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15738" *) IsNaN_8U_23U_land_3_lpi_1_dfm_11;
  assign _2007_ = _2006_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15738" *) _1205_;
  assign _2008_ = _2007_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15739" *) FpAlu_8U_23U_equal_tmp_23;
  assign _2009_ = _2008_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15739" *) io_read_cfg_alu_bypass_rsc_svs_st_7;
  assign _2010_ = _2009_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15739" *) FpAdd_8U_23U_is_inf_3_lpi_1_dfm_8;
  assign _2011_ = _1424_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15740" *) alu_loop_op_unequal_tmp_8;
  assign _2012_ = or_323_nl | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15742" *) mux_85_nl;
  assign _2013_ = nor_45_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15744" *) _1203_;
  assign _2014_ = _2013_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15745" *) io_read_cfg_alu_bypass_rsc_svs_st_6;
  assign _2015_ = _2014_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15745" *) _1148_;
  assign _2016_ = _2015_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15745" *) io_read_cfg_alu_bypass_rsc_svs_7;
  assign _2017_ = _2016_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15746" *) alu_loop_op_unequal_tmp_7;
  assign _2018_ = _2017_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15746" *) _1202_;
  assign _2019_ = _2018_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15746" *) FpAlu_8U_23U_equal_tmp_22;
  assign _2020_ = _2019_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15747" *) IsNaN_8U_23U_1_land_lpi_1_dfm_8;
  assign _2021_ = _2020_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15747" *) IsNaN_8U_23U_land_lpi_1_dfm_10;
  assign _2022_ = FpAdd_8U_23U_int_mant_p1_lpi_1_dfm_5[49] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15749" *) _1203_;
  assign _2023_ = _2022_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15749" *) io_read_cfg_alu_bypass_rsc_svs_st_6;
  assign _2024_ = _2023_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15749" *) _1148_;
  assign _2025_ = _2024_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15750" *) io_read_cfg_alu_bypass_rsc_svs_7;
  assign _2026_ = _2025_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15750" *) alu_loop_op_unequal_tmp_7;
  assign _2027_ = _2026_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15751" *) _1202_;
  assign _2028_ = _2027_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15751" *) FpAlu_8U_23U_equal_tmp_22;
  assign _2029_ = _2028_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15751" *) IsNaN_8U_23U_1_land_lpi_1_dfm_8;
  assign _2030_ = _2029_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15751" *) IsNaN_8U_23U_land_lpi_1_dfm_10;
  assign _2031_ = _1220_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15753" *) alu_loop_op_4_FpAdd_8U_23U_if_4_if_acc_6_nl[7];
  assign _2032_ = _1884_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15756" *) io_read_cfg_alu_bypass_rsc_svs_7;
  assign _2033_ = _2032_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15757" *) alu_loop_op_unequal_tmp_7;
  assign _2034_ = _2033_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15757" *) _1202_;
  assign _2035_ = _2034_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15757" *) FpAlu_8U_23U_equal_tmp_22;
  assign _2036_ = _2035_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15758" *) IsNaN_8U_23U_1_land_lpi_1_dfm_8;
  assign _2037_ = _2036_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15758" *) IsNaN_8U_23U_land_lpi_1_dfm_10;
  assign _2038_ = _1425_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15762" *) _1426_;
  assign _2039_ = _2038_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15762" *) or_236_nl;
  assign _2040_ = _2039_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15762" *) IsNaN_8U_23U_1_land_lpi_1_dfm_9;
  assign or_182_nl = _2040_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15762" *) IsNaN_8U_23U_land_lpi_1_dfm_11;
  assign _2041_ = _1503_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15766" *) _1205_;
  assign _2042_ = _2041_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15766" *) FpAlu_8U_23U_equal_tmp_23;
  assign _2043_ = _2042_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15767" *) io_read_cfg_alu_bypass_rsc_svs_st_7;
  assign _2044_ = _2043_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15767" *) FpAdd_8U_23U_is_inf_lpi_1_dfm_8;
  assign _2045_ = _2044_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15767" *) mux_91_nl;
  assign _2046_ = _1219_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15770" *) _1203_;
  assign _2047_ = _2046_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15770" *) io_read_cfg_alu_bypass_rsc_svs_st_6;
  assign _2048_ = _2047_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15770" *) _1148_;
  assign _2049_ = _1427_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15772" *) _1203_;
  assign _2050_ = _2049_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15772" *) io_read_cfg_alu_bypass_rsc_svs_st_6;
  assign _2051_ = _2050_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15772" *) _1148_;
  assign _2052_ = or_tmp_224 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15775" *) cfg_alu_algo_1_sva_st_25[0];
  assign _2053_ = _2052_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15775" *) _1428_;
  assign _2054_ = _1218_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15778" *) _1203_;
  assign _2055_ = _2054_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15778" *) io_read_cfg_alu_bypass_rsc_svs_st_6;
  assign _2056_ = _2055_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15778" *) _1148_;
  assign _2057_ = _1429_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15780" *) _1203_;
  assign _2058_ = _2057_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15780" *) io_read_cfg_alu_bypass_rsc_svs_st_6;
  assign _2059_ = _2058_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15780" *) _1148_;
  assign _2060_ = _2052_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15783" *) _1430_;
  assign _2061_ = _1215_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15786" *) _1203_;
  assign _2062_ = _2061_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15786" *) io_read_cfg_alu_bypass_rsc_svs_st_6;
  assign _2063_ = _2062_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15786" *) _1148_;
  assign _2064_ = _1431_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15788" *) _1203_;
  assign _2065_ = _2064_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15788" *) io_read_cfg_alu_bypass_rsc_svs_st_6;
  assign _2066_ = _2065_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15788" *) _1148_;
  assign _2067_ = _2052_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15791" *) _1432_;
  assign _2068_ = _1220_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15794" *) _1203_;
  assign _2069_ = _2068_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15794" *) io_read_cfg_alu_bypass_rsc_svs_st_6;
  assign _2070_ = _2069_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15794" *) _1148_;
  assign _2071_ = _1433_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15796" *) _1203_;
  assign _2072_ = _2071_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15796" *) io_read_cfg_alu_bypass_rsc_svs_st_6;
  assign _2073_ = _2072_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15796" *) _1148_;
  assign _2074_ = _2052_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15799" *) _1434_;
  assign _2075_ = _1835_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15802" *) alu_loop_op_unequal_tmp_8;
  assign or_1100_nl = _2075_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15802" *) FpAlu_8U_23U_nor_dfs_6;
  assign _2076_ = alu_loop_op_unequal_tmp_8 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15803" *) _1205_;
  assign _2077_ = _1435_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15804" *) or_dcpl_272;
  assign or_1106_nl = _2077_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15804" *) FpAlu_8U_23U_equal_tmp_23;
  assign _2078_ = _1281_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15807" *) _1216_;
  assign _2079_ = _2078_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15807" *) alu_loop_op_unequal_tmp_8;
  assign _2080_ = _2079_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15807" *) io_read_cfg_alu_bypass_rsc_svs_8;
  assign or_280_nl = _2080_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15807" *) _1206_;
  assign _2081_ = _1501_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15811" *) _1202_;
  assign _2082_ = _2081_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15811" *) FpAlu_8U_23U_equal_tmp_22;
  assign _2083_ = _2082_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15811" *) _1209_;
  assign _2084_ = _2083_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15811" *) IsNaN_8U_23U_land_3_lpi_1_dfm_10;
  assign _2085_ = _2043_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15814" *) _1436_;
  assign _2086_ = _2085_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15814" *) IsNaN_8U_23U_land_3_lpi_1_dfm_11;
  assign _2087_ = _2082_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15818" *) _1210_;
  assign _2088_ = _2087_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15818" *) IsNaN_8U_23U_land_2_lpi_1_dfm_10;
  assign _2089_ = _2043_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15821" *) _1437_;
  assign _2090_ = _2089_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15821" *) IsNaN_8U_23U_land_2_lpi_1_dfm_11;
  assign _2091_ = _2082_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15825" *) _1211_;
  assign _2092_ = _2091_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15825" *) IsNaN_8U_23U_land_1_lpi_1_dfm_10;
  assign _2093_ = _2043_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15828" *) _1438_;
  assign _2094_ = _2093_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15828" *) IsNaN_8U_23U_land_1_lpi_1_dfm_11;
  assign _2095_ = _1213_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15831" *) io_read_cfg_alu_bypass_rsc_svs_st_7;
  assign _2096_ = _2095_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15831" *) alu_loop_op_unequal_tmp_8;
  assign _2097_ = _2096_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15831" *) io_read_cfg_alu_bypass_rsc_svs_8;
  assign or_299_nl = _2097_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15831" *) _1206_;
  assign _2098_ = _1517_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15834" *) io_read_cfg_alu_bypass_rsc_svs_st_7;
  assign _2099_ = _2098_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15835" *) alu_loop_op_unequal_tmp_8;
  assign _2100_ = _2099_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15835" *) io_read_cfg_alu_bypass_rsc_svs_8;
  assign or_301_nl = _2100_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15835" *) _1206_;
  assign _2101_ = _1364_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15837" *) alu_loop_op_unequal_tmp_7;
  assign _2102_ = _2101_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15838" *) io_read_cfg_alu_bypass_rsc_svs_7;
  assign _2103_ = _2102_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15838" *) io_read_cfg_alu_bypass_rsc_svs_st_6;
  assign or_304_nl = _2103_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15839" *) _1203_;
  assign _2104_ = nor_269_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15841" *) _1364_;
  assign _2105_ = _2104_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15842" *) alu_loop_op_unequal_tmp_7;
  assign _2106_ = _2105_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15842" *) io_read_cfg_alu_bypass_rsc_svs_7;
  assign _2107_ = _2106_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15842" *) io_read_cfg_alu_bypass_rsc_svs_st_6;
  assign or_307_nl = _2107_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15843" *) _1203_;
  assign _2108_ = _1439_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15846" *) _1281_;
  assign _2109_ = _2108_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15846" *) _1216_;
  assign _2110_ = _2109_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15846" *) io_read_cfg_alu_bypass_rsc_svs_st_7;
  assign _2111_ = _2110_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15847" *) alu_loop_op_unequal_tmp_8;
  assign _2112_ = _2111_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15847" *) io_read_cfg_alu_bypass_rsc_svs_8;
  assign or_312_nl = _2112_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15847" *) _1206_;
  assign _2113_ = _2082_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15851" *) _1200_;
  assign _2114_ = _2113_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15851" *) IsNaN_8U_23U_land_lpi_1_dfm_10;
  assign _2115_ = _2043_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15854" *) _1440_;
  assign _2116_ = _2115_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15854" *) IsNaN_8U_23U_land_lpi_1_dfm_11;
  assign or_1046_nl = main_stage_v_4 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15860" *) nor_tmp_144;
  assign _2117_ = alu_loop_op_unequal_tmp_8 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15861" *) FpAlu_8U_23U_equal_tmp_23;
  assign _2118_ = _2117_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15862" *) FpAlu_8U_23U_nor_dfs_6;
  assign _2119_ = _2118_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15862" *) FpAlu_8U_23U_equal_tmp_26;
  assign _2120_ = _2119_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15862" *) FpAlu_8U_23U_equal_tmp_29;
  assign or_1048_nl = _2120_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15862" *) nor_tmp_144;
  assign or_333_nl = alu_loop_op_1_FpMantRNE_49U_24U_else_and_tmp | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15867" *) or_tmp_315;
  assign or_334_nl = alu_loop_op_2_FpMantRNE_49U_24U_else_and_2_tmp | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15870" *) or_tmp_315;
  assign or_335_nl = alu_loop_op_3_FpMantRNE_49U_24U_else_and_1_tmp | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15873" *) or_tmp_315;
  assign or_336_nl = alu_loop_op_4_FpMantRNE_49U_24U_else_and_3_tmp | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15876" *) or_tmp_315;
  assign _2121_ = or_dcpl_86 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15880" *) IsNaN_8U_23U_land_1_lpi_1_dfm_st_4;
  assign _2122_ = _2121_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15880" *) _1235_;
  assign _2123_ = _2122_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15880" *) IsNaN_8U_23U_land_1_lpi_1_dfm_9;
  assign _2124_ = _2123_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15881" *) _1194_;
  assign _2125_ = _2124_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15881" *) io_read_cfg_alu_bypass_rsc_svs_st_5;
  assign _2126_ = _2125_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15881" *) io_read_cfg_alu_bypass_rsc_svs_6;
  assign _2127_ = _2126_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15882" *) alu_loop_op_unequal_tmp_6;
  assign _2128_ = _1148_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15886" *) IsNaN_8U_23U_land_1_lpi_1_dfm_st_5;
  assign _2129_ = _2128_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15887" *) _1202_;
  assign _2130_ = _2129_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15887" *) IsNaN_8U_23U_land_1_lpi_1_dfm_10;
  assign _2131_ = _1501_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15887" *) _0899_;
  assign _2132_ = or_dcpl_86 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15890" *) IsNaN_8U_23U_land_2_lpi_1_dfm_st_4;
  assign _2133_ = _2132_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15890" *) _1235_;
  assign _2134_ = _2133_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15890" *) IsNaN_8U_23U_land_2_lpi_1_dfm_9;
  assign _2135_ = _2134_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15891" *) _1194_;
  assign _2136_ = _2135_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15891" *) io_read_cfg_alu_bypass_rsc_svs_st_5;
  assign _2137_ = _2136_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15891" *) io_read_cfg_alu_bypass_rsc_svs_6;
  assign _2138_ = _2137_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15892" *) alu_loop_op_unequal_tmp_6;
  assign _2139_ = _1148_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15896" *) IsNaN_8U_23U_land_2_lpi_1_dfm_st_5;
  assign _2140_ = _2139_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15897" *) _1202_;
  assign _2141_ = _2140_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15897" *) IsNaN_8U_23U_land_2_lpi_1_dfm_10;
  assign _2142_ = _1501_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15897" *) _0900_;
  assign _2143_ = or_dcpl_86 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15900" *) IsNaN_8U_23U_land_3_lpi_1_dfm_st_4;
  assign _2144_ = _2143_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15900" *) _1235_;
  assign _2145_ = _2144_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15900" *) IsNaN_8U_23U_land_3_lpi_1_dfm_9;
  assign _2146_ = _2145_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15901" *) _1194_;
  assign _2147_ = _2146_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15901" *) io_read_cfg_alu_bypass_rsc_svs_st_5;
  assign _2148_ = _2147_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15901" *) io_read_cfg_alu_bypass_rsc_svs_6;
  assign _2149_ = _2148_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15902" *) alu_loop_op_unequal_tmp_6;
  assign _2150_ = _1148_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15906" *) IsNaN_8U_23U_land_3_lpi_1_dfm_st_5;
  assign _2151_ = _2150_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15907" *) _1202_;
  assign _2152_ = _2151_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15907" *) IsNaN_8U_23U_land_3_lpi_1_dfm_10;
  assign _2153_ = _1501_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15907" *) _0901_;
  assign _2154_ = or_dcpl_86 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15910" *) IsNaN_8U_23U_land_lpi_1_dfm_st_4;
  assign _2155_ = _2154_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15910" *) _1235_;
  assign _2156_ = _2155_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15910" *) IsNaN_8U_23U_land_lpi_1_dfm_9;
  assign _2157_ = _2156_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15911" *) _1194_;
  assign _2158_ = _2157_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15911" *) io_read_cfg_alu_bypass_rsc_svs_st_5;
  assign _2159_ = _2158_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15911" *) io_read_cfg_alu_bypass_rsc_svs_6;
  assign _2160_ = _2159_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15912" *) alu_loop_op_unequal_tmp_6;
  assign _2161_ = _1148_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15916" *) IsNaN_8U_23U_land_lpi_1_dfm_st_5;
  assign _2162_ = _2161_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15917" *) _1202_;
  assign _2163_ = _2162_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15917" *) IsNaN_8U_23U_land_lpi_1_dfm_10;
  assign _2164_ = _1501_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15917" *) _0902_;
  assign _2165_ = acc_12_nl[50] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15919" *) or_dcpl_86;
  assign _2166_ = _2165_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15920" *) io_read_cfg_alu_bypass_rsc_svs_st_5;
  assign _2167_ = _2166_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15920" *) or_tmp_347;
  assign _2168_ = _1443_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15921" *) or_dcpl_86;
  assign _2169_ = _2168_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15922" *) io_read_cfg_alu_bypass_rsc_svs_st_5;
  assign or_961_nl = _2169_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15922" *) or_tmp_347;
  assign _2170_ = acc_13_nl[50] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15924" *) or_dcpl_86;
  assign _2171_ = _2170_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15925" *) io_read_cfg_alu_bypass_rsc_svs_st_5;
  assign _2172_ = _2171_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15925" *) or_tmp_347;
  assign _2173_ = _1444_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15926" *) or_dcpl_86;
  assign _2174_ = _2173_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15927" *) io_read_cfg_alu_bypass_rsc_svs_st_5;
  assign or_960_nl = _2174_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15927" *) or_tmp_347;
  assign _2175_ = acc_14_nl[50] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15929" *) or_dcpl_86;
  assign _2176_ = _2175_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15930" *) io_read_cfg_alu_bypass_rsc_svs_st_5;
  assign _2177_ = _2176_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15930" *) or_tmp_347;
  assign _2178_ = _1445_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15931" *) or_dcpl_86;
  assign _2179_ = _2178_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15932" *) io_read_cfg_alu_bypass_rsc_svs_st_5;
  assign or_959_nl = _2179_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15932" *) or_tmp_347;
  assign _2180_ = acc_15_nl[50] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15934" *) or_dcpl_86;
  assign _2181_ = _2180_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15935" *) io_read_cfg_alu_bypass_rsc_svs_st_5;
  assign _2182_ = _2181_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15935" *) or_tmp_347;
  assign _2183_ = _1446_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15936" *) or_dcpl_86;
  assign _2184_ = _2183_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15937" *) io_read_cfg_alu_bypass_rsc_svs_st_5;
  assign or_958_nl = _2184_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15937" *) or_tmp_347;
  assign IntSaturation_33U_32U_IntSaturation_33U_32U_or_nl = _0903_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15943" *) alu_loop_op_1_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_svs_2;
  assign or_422_nl = or_1087_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15945" *) mux_tmp_164;
  assign or_420_nl = _1448_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15946" *) io_read_cfg_alu_bypass_rsc_svs_st_5;
  assign IntSaturation_33U_32U_IntSaturation_33U_32U_or_3_nl = _0904_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15950" *) alu_loop_op_4_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_1_svs_2;
  assign IntSaturation_33U_32U_IntSaturation_33U_32U_or_2_nl = _0905_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15952" *) alu_loop_op_3_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_svs_2;
  assign IntSaturation_33U_32U_IntSaturation_33U_32U_or_1_nl = _0906_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15954" *) alu_loop_op_2_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_1_svs_3;
  assign or_438_nl = or_tmp_409 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15955" *) or_tmp_416;
  assign _2185_ = _1538_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15959" *) io_read_cfg_alu_bypass_rsc_svs_st_6;
  assign or_440_nl = _2185_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15959" *) _1203_;
  assign _2186_ = or_1087_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15962" *) _1320_;
  assign _2187_ = _2186_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15962" *) _1319_;
  assign _2188_ = _2187_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15963" *) _1242_;
  assign _2189_ = _2188_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15963" *) alu_loop_op_unequal_tmp_7;
  assign _2190_ = _2189_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15963" *) io_read_cfg_alu_bypass_rsc_svs_7;
  assign _2191_ = _2190_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15964" *) io_read_cfg_alu_bypass_rsc_svs_st_6;
  assign or_446_nl = _2191_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15964" *) _1203_;
  assign _2192_ = alu_loop_op_unequal_tmp_6 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15966" *) _1452_;
  assign _2193_ = _2192_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15967" *) _1453_;
  assign _2194_ = _2193_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15967" *) _1243_;
  assign or_444_nl = _2194_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15967" *) io_read_cfg_alu_bypass_rsc_svs_st_5;
  assign _2195_ = or_1087_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15971" *) _1319_;
  assign _2196_ = _2195_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15971" *) _1242_;
  assign _2197_ = _2196_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15972" *) alu_loop_op_unequal_tmp_7;
  assign _2198_ = _2197_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15972" *) io_read_cfg_alu_bypass_rsc_svs_7;
  assign or_450_nl = _2198_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15972" *) _1203_;
  assign _2199_ = alu_loop_op_unequal_tmp_6 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15974" *) _1453_;
  assign _2200_ = _2199_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15974" *) _1243_;
  assign _2201_ = io_read_cfg_alu_bypass_rsc_svs_st_5 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15977" *) _1235_;
  assign _2202_ = _2201_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15977" *) FpAlu_8U_23U_equal_tmp_21;
  assign _2203_ = _2202_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15977" *) _1454_;
  assign _2204_ = _2203_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15978" *) IsNaN_8U_23U_land_3_lpi_1_dfm_9;
  assign _2205_ = _2204_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15978" *) _1194_;
  assign _2206_ = _2205_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15978" *) io_read_cfg_alu_bypass_rsc_svs_6;
  assign _2207_ = io_read_cfg_alu_bypass_rsc_svs_st_6 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15981" *) _1202_;
  assign _2208_ = _2207_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15982" *) FpAlu_8U_23U_equal_tmp_22;
  assign _2209_ = _2208_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15982" *) _1209_;
  assign _2210_ = _2209_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15982" *) IsNaN_8U_23U_land_3_lpi_1_dfm_10;
  assign _2211_ = alu_loop_op_unequal_tmp_7 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15982" *) _1455_;
  assign _2212_ = or_417_nl | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15982" *) _1456_;
  assign _2213_ = _2202_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15985" *) _1457_;
  assign _2214_ = _2213_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15986" *) IsNaN_8U_23U_land_lpi_1_dfm_9;
  assign _2215_ = _2214_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15986" *) _1194_;
  assign _2216_ = _2215_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15986" *) io_read_cfg_alu_bypass_rsc_svs_6;
  assign _2217_ = _2208_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15990" *) _1200_;
  assign _2218_ = _2217_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15990" *) IsNaN_8U_23U_land_lpi_1_dfm_10;
  assign _2219_ = alu_loop_op_unequal_tmp_7 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15990" *) _1458_;
  assign _2220_ = or_417_nl | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15990" *) _1459_;
  assign _2221_ = _2202_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15993" *) _1460_;
  assign _2222_ = _2221_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15994" *) IsNaN_8U_23U_land_2_lpi_1_dfm_9;
  assign _2223_ = _2222_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15994" *) _1194_;
  assign _2224_ = _2223_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15994" *) io_read_cfg_alu_bypass_rsc_svs_6;
  assign _2225_ = _2208_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15998" *) _1210_;
  assign _2226_ = _2225_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15998" *) IsNaN_8U_23U_land_2_lpi_1_dfm_10;
  assign _2227_ = alu_loop_op_unequal_tmp_7 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15998" *) _1461_;
  assign _2228_ = or_417_nl | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15998" *) _1462_;
  assign _2229_ = _2202_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16001" *) _1463_;
  assign _2230_ = _2229_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16002" *) IsNaN_8U_23U_land_1_lpi_1_dfm_9;
  assign _2231_ = _2230_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16002" *) _1194_;
  assign _2232_ = _2231_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16002" *) io_read_cfg_alu_bypass_rsc_svs_6;
  assign _2233_ = _2208_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16006" *) _1211_;
  assign _2234_ = _2233_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16006" *) IsNaN_8U_23U_land_1_lpi_1_dfm_10;
  assign _2235_ = alu_loop_op_unequal_tmp_7 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16006" *) _1464_;
  assign _2236_ = or_417_nl | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16006" *) _1465_;
  assign _2237_ = _1728_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16011" *) IsNaN_8U_23U_land_1_lpi_1_dfm_st_4;
  assign _2238_ = _2237_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16012" *) io_read_cfg_alu_bypass_rsc_svs_6;
  assign _2239_ = _2238_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16012" *) alu_loop_op_unequal_tmp_6;
  assign _2240_ = _2239_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16013" *) _1235_;
  assign _2241_ = _2240_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16013" *) _1463_;
  assign _2242_ = _2241_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16013" *) IsNaN_8U_23U_land_1_lpi_1_dfm_9;
  assign _2243_ = _1884_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16015" *) IsNaN_8U_23U_land_1_lpi_1_dfm_st_5;
  assign _2244_ = _2243_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16016" *) io_read_cfg_alu_bypass_rsc_svs_7;
  assign _2245_ = _2244_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16016" *) alu_loop_op_unequal_tmp_7;
  assign _2246_ = _2245_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16017" *) _1202_;
  assign _2247_ = _2246_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16017" *) _1211_;
  assign _2248_ = _2247_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16017" *) IsNaN_8U_23U_land_1_lpi_1_dfm_10;
  assign _2249_ = _1728_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16020" *) IsNaN_8U_23U_land_2_lpi_1_dfm_st_4;
  assign _2250_ = _2249_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16021" *) io_read_cfg_alu_bypass_rsc_svs_6;
  assign _2251_ = _2250_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16021" *) alu_loop_op_unequal_tmp_6;
  assign _2252_ = _2251_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16022" *) _1235_;
  assign _2253_ = _2252_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16022" *) _1460_;
  assign _2254_ = _2253_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16022" *) IsNaN_8U_23U_land_2_lpi_1_dfm_9;
  assign _2255_ = _1884_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16024" *) IsNaN_8U_23U_land_2_lpi_1_dfm_st_5;
  assign _2256_ = _2255_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16025" *) io_read_cfg_alu_bypass_rsc_svs_7;
  assign _2257_ = _2256_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16025" *) alu_loop_op_unequal_tmp_7;
  assign _2258_ = _2257_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16026" *) _1202_;
  assign _2259_ = _2258_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16026" *) _1210_;
  assign _2260_ = _2259_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16026" *) IsNaN_8U_23U_land_2_lpi_1_dfm_10;
  assign _2261_ = _1728_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16029" *) IsNaN_8U_23U_land_3_lpi_1_dfm_st_4;
  assign _2262_ = _2261_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16030" *) io_read_cfg_alu_bypass_rsc_svs_6;
  assign _2263_ = _2262_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16030" *) alu_loop_op_unequal_tmp_6;
  assign _2264_ = _2263_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16031" *) _1235_;
  assign _2265_ = _2264_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16031" *) _1454_;
  assign _2266_ = _2265_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16031" *) IsNaN_8U_23U_land_3_lpi_1_dfm_9;
  assign _2267_ = _1884_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16033" *) IsNaN_8U_23U_land_3_lpi_1_dfm_st_5;
  assign _2268_ = _2267_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16034" *) io_read_cfg_alu_bypass_rsc_svs_7;
  assign _2269_ = _2268_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16034" *) alu_loop_op_unequal_tmp_7;
  assign _2270_ = _2269_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16035" *) _1202_;
  assign _2271_ = _2270_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16035" *) _1209_;
  assign _2272_ = _2271_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16035" *) IsNaN_8U_23U_land_3_lpi_1_dfm_10;
  assign _2273_ = _1728_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16038" *) IsNaN_8U_23U_land_lpi_1_dfm_st_4;
  assign _2274_ = _2273_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16039" *) io_read_cfg_alu_bypass_rsc_svs_6;
  assign _2275_ = _2274_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16039" *) alu_loop_op_unequal_tmp_6;
  assign _2276_ = _2275_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16039" *) _1235_;
  assign _2277_ = _2276_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16040" *) _1457_;
  assign _2278_ = _2277_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16040" *) IsNaN_8U_23U_land_lpi_1_dfm_9;
  assign _2279_ = _1884_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16042" *) IsNaN_8U_23U_land_lpi_1_dfm_st_5;
  assign _2280_ = _2279_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16043" *) io_read_cfg_alu_bypass_rsc_svs_7;
  assign _2281_ = _2280_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16043" *) alu_loop_op_unequal_tmp_7;
  assign _2282_ = _2281_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16043" *) _1202_;
  assign _2283_ = _2282_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16044" *) _1200_;
  assign _2284_ = _2283_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16044" *) IsNaN_8U_23U_land_lpi_1_dfm_10;
  assign FpAlu_8U_23U_or_145_nl = _0907_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16047" *) _0908_;
  assign FpAlu_8U_23U_or_146_nl = _0909_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16049" *) _0910_;
  assign FpAlu_8U_23U_or_147_nl = _0911_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16055" *) _0912_;
  assign FpAlu_8U_23U_or_148_nl = _0913_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16057" *) _0914_;
  assign _2285_ = _1523_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16063" *) _1448_;
  assign _2286_ = _1573_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16066" *) _1448_;
  assign AluOut_data_or_1_nl = and_dcpl_207 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16070" *) _0915_;
  assign AluOut_data_or_2_nl = AluOut_data_and_5_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16074" *) _0916_;
  assign AluOut_data_or_nl = and_dcpl_207 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16080" *) _0917_;
  assign AluOut_data_or_3_nl = AluOut_data_and_5_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16084" *) _0918_;
  assign _2287_ = _1523_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16089" *) _1255_;
  assign _2288_ = _1566_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16092" *) _1167_;
  assign _2289_ = _2288_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16093" *) _1248_;
  assign _2290_ = _2289_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16094" *) _1249_;
  assign _2291_ = _2290_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16094" *) _1250_;
  assign _2292_ = _2291_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16095" *) _1251_;
  assign _2293_ = _2292_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16095" *) io_read_cfg_alu_bypass_rsc_svs_5;
  assign _2294_ = _2288_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16099" *) or_dcpl_154;
  assign _2295_ = _2294_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16100" *) _1248_;
  assign _2296_ = _2295_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16100" *) _1249_;
  assign _2297_ = _2296_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16101" *) _1250_;
  assign _2298_ = _2297_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16101" *) _1251_;
  assign _2299_ = _2298_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16101" *) io_read_cfg_alu_bypass_rsc_svs_5;
  assign or_1069_nl = or_1055_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16107" *) _1167_;
  assign or_1076_nl = or_1069_nl | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16111" *) or_dcpl_154;
  assign _2300_ = _0919_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16115" *) _0920_;
  assign _2301_ = _0921_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16118" *) _0922_;
  assign _2302_ = _0923_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16129" *) _0924_;
  assign _2303_ = _0925_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16132" *) _0926_;
  assign _2304_ = or_1050_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16145" *) cfg_alu_bypass_rsci_d;
  assign _2305_ = _2304_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16145" *) _1188_;
  assign _2306_ = _1471_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16146" *) cfg_alu_algo_1_sva_st[1];
  assign or_624_nl = _2306_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16146" *) not_tmp_259;
  assign or_619_nl = or_1069_nl | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16150" *) io_read_cfg_alu_bypass_rsc_svs_5;
  assign _2307_ = and_501_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16157" *) mux_tmp_268;
  assign _2308_ = and_501_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16168" *) mux_tmp_281;
  assign _2309_ = _0932_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16265" *) _0943_;
  assign _2310_ = _0933_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16265" *) _0944_;
  assign _2311_ = _0934_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16265" *) _0945_;
  assign _2312_ = _0935_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16265" *) _0946_;
  assign _2313_ = _0936_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16265" *) _0947_;
  assign _2314_ = _0937_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16265" *) _0948_;
  assign _2315_ = _0938_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16265" *) _0949_;
  assign _2316_ = _0939_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16265" *) _0950_;
  assign _2317_ = _0940_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16265" *) _0951_;
  assign _2318_ = _0941_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16265" *) _0952_;
  assign _2319_ = _0942_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16265" *) _0953_;
  assign _2320_ = _2309_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16266" *) _0954_;
  assign _2321_ = _2310_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16266" *) _0955_;
  assign _2322_ = _2311_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16266" *) _0956_;
  assign _2323_ = _2312_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16266" *) _0957_;
  assign _2324_ = _2313_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16266" *) _0958_;
  assign _2325_ = _2314_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16266" *) _0959_;
  assign _2326_ = _2315_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16266" *) _0960_;
  assign _2327_ = _2316_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16266" *) _0961_;
  assign _2328_ = _2317_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16266" *) _0962_;
  assign _2329_ = _2318_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16266" *) _0963_;
  assign _2330_ = _2319_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16266" *) _0964_;
  assign _2331_ = _0965_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16279" *) _0975_;
  assign _2332_ = _0966_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16279" *) _0976_;
  assign _2333_ = _0967_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16279" *) _0977_;
  assign _2334_ = _0968_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16279" *) _0978_;
  assign _2335_ = _0969_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16279" *) _0979_;
  assign _2336_ = _0970_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16279" *) _0980_;
  assign _2337_ = _0971_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16279" *) _0981_;
  assign _2338_ = _0972_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16279" *) _0982_;
  assign _2339_ = _0973_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16279" *) _0983_;
  assign _2340_ = _0974_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16279" *) _0984_;
  assign _2341_ = _2331_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16280" *) _0985_;
  assign _2342_ = _2332_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16280" *) _0986_;
  assign _2343_ = _2333_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16280" *) _0987_;
  assign _2344_ = _2334_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16280" *) _0988_;
  assign _2345_ = _2335_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16280" *) _0989_;
  assign _2346_ = _2336_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16280" *) _0990_;
  assign _2347_ = _2337_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16280" *) _0991_;
  assign _2348_ = _2338_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16280" *) _0992_;
  assign _2349_ = _2339_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16280" *) _0993_;
  assign _2350_ = _2340_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16280" *) _0994_;
  assign _2351_ = _2341_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16281" *) _0995_;
  assign _2352_ = _2342_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16281" *) _0996_;
  assign _2353_ = _2343_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16281" *) _0997_;
  assign _2354_ = _2344_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16281" *) _0998_;
  assign _2355_ = _2345_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16281" *) _0999_;
  assign _2356_ = _2346_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16281" *) _1000_;
  assign FpAlu_8U_23U_mux1h_147_nl = _2347_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16281" *) _1001_;
  assign FpAlu_8U_23U_mux1h_151_nl = _2348_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16281" *) _1002_;
  assign FpAlu_8U_23U_mux1h_144_nl = _2349_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16281" *) _1003_;
  assign FpAlu_8U_23U_mux1h_148_nl = _2350_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16281" *) _1004_;
  assign _2357_ = _1005_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16295" *) _1007_;
  assign _2358_ = _1006_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16295" *) _1008_;
  assign _2359_ = _2357_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16296" *) _1009_;
  assign _2360_ = _2358_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16296" *) _1010_;
  assign _2361_ = _2359_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16297" *) _1011_;
  assign _2362_ = _2360_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16297" *) _1012_;
  assign FpAlu_8U_23U_mux1h_155_nl = _2361_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16298" *) _1013_;
  assign FpAlu_8U_23U_o_0_lpi_1_dfm_2 = _2362_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16298" *) _1014_;
  assign _2363_ = _1015_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16314" *) _1017_;
  assign _2364_ = _1016_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16314" *) _1018_;
  assign _2365_ = _2363_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16315" *) _1019_;
  assign _2366_ = _2364_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16315" *) _1020_;
  assign _2367_ = _2365_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16316" *) _1021_;
  assign _2368_ = _2366_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16316" *) _1022_;
  assign _2369_ = _2367_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16317" *) _1023_;
  assign _2370_ = _2368_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16317" *) _1024_;
  assign _2371_ = _2369_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16318" *) _1025_;
  assign _2372_ = _2370_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16318" *) _1026_;
  assign _2373_ = _2371_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16319" *) _1027_;
  assign _2374_ = _2372_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16319" *) _1028_;
  assign _2375_ = _1029_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16331" *) _1034_;
  assign _2376_ = _1030_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16331" *) _1035_;
  assign _2377_ = _1031_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16331" *) _1036_;
  assign _2378_ = _1032_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16331" *) _1037_;
  assign _2379_ = _1033_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16331" *) _1038_;
  assign _2380_ = _2375_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16332" *) _1039_;
  assign _2381_ = _2376_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16332" *) _1040_;
  assign _2382_ = _2377_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16332" *) _1041_;
  assign FpAlu_8U_23U_mux1h_154_nl = _2378_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16332" *) _1042_;
  assign AluOut_data_2_22_1_lpi_1_dfm_3_mx1w0 = _2379_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16332" *) _1043_;
  assign _2383_ = _1044_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16345" *) _1045_;
  assign _2384_ = _2383_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16346" *) _1046_;
  assign FpAlu_8U_23U_mux1h_35_nl = _2384_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16347" *) _1047_;
  assign _2385_ = _1048_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16359" *) _1052_;
  assign _2386_ = _1049_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16359" *) _1053_;
  assign _2387_ = _1050_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16359" *) _1054_;
  assign _2388_ = _1051_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16359" *) _1055_;
  assign IntSaturation_33U_32U_o_31_1_2_lpi_1_dfm_1 = _2385_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16360" *) _1056_;
  assign IntSaturation_33U_32U_o_31_1_lpi_1_dfm_1 = _2386_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16360" *) _1057_;
  assign IntSaturation_33U_32U_o_31_1_3_lpi_1_dfm_1 = _2387_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16360" *) _1058_;
  assign IntSaturation_33U_32U_o_31_1_1_lpi_1_dfm_1 = _2388_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16360" *) { _1135_[30:7], _1059_ };
  assign _2389_ = _1060_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16372" *) _1076_;
  assign _2390_ = _1061_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16372" *) _1077_;
  assign _2391_ = _1062_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16372" *) _1078_;
  assign _2392_ = _1063_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16372" *) _1079_;
  assign _2393_ = _1064_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16372" *) _1080_;
  assign _2394_ = _1065_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16372" *) _1081_;
  assign _2395_ = _1066_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16372" *) _1082_;
  assign _2396_ = _1067_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16372" *) _1083_;
  assign _2397_ = _1068_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16372" *) _1084_;
  assign _2398_ = _1069_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16372" *) _1085_;
  assign _2399_ = _1070_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16372" *) _1086_;
  assign _2400_ = _1071_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16372" *) _1087_;
  assign _2401_ = _1072_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16372" *) _1088_;
  assign _2402_ = _1073_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16372" *) _1089_;
  assign _2403_ = _1074_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16372" *) _1090_;
  assign _2404_ = _1075_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16372" *) _1091_;
  assign _2405_ = _2389_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16373" *) _1092_;
  assign _2406_ = _2390_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16373" *) _1093_;
  assign _2407_ = _2391_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16373" *) _1094_;
  assign _2408_ = _2392_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16373" *) _1095_;
  assign _2409_ = _2393_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16373" *) _1096_;
  assign _2410_ = _2394_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16373" *) _1097_;
  assign _2411_ = _2395_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16373" *) _1098_;
  assign _2412_ = _2396_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16373" *) _1099_;
  assign _2413_ = _2397_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16373" *) _1100_;
  assign _2414_ = _2398_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16373" *) _1101_;
  assign _2415_ = _2399_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16373" *) _1102_;
  assign AluOut_data_2_30_23_lpi_1_dfm_3_mx1w0 = _2400_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16373" *) _1103_;
  assign FpAdd_8U_23U_o_expo_1_lpi_1_dfm_2_mx0w0 = _2401_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16373" *) _1104_;
  assign FpAdd_8U_23U_o_expo_2_lpi_1_dfm_2_mx0w0 = _2402_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16373" *) _1105_;
  assign FpAdd_8U_23U_o_expo_3_lpi_1_dfm_2_mx0w0 = _2403_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16373" *) _1106_;
  assign FpAdd_8U_23U_o_expo_lpi_1_dfm_2_mx0w0 = _2404_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16373" *) _1107_;
  assign _2416_ = _1108_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16388" *) _1110_;
  assign _2417_ = _1109_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16388" *) _1111_;
  assign _2418_ = _2416_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16389" *) _1112_;
  assign _2419_ = _2417_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16389" *) _1113_;
  assign _2420_ = _2418_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16390" *) _1114_;
  assign _2421_ = _2419_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16390" *) _1115_;
  assign _2422_ = _2420_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16391" *) _1116_;
  assign _2423_ = _2421_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16391" *) _1117_;
  assign FpAlu_8U_23U_mux1h_145_nl = _2422_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16392" *) _1118_;
  assign FpAlu_8U_23U_mux1h_149_nl = _2423_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16392" *) _1119_;
  assign _2424_ = _1120_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16408" *) _1121_;
  assign _2425_ = _2424_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16409" *) _1122_;
  assign _2426_ = _2425_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16410" *) _1123_;
  assign _2427_ = _2426_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16411" *) _1124_;
  assign _2428_ = _2427_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16412" *) _1125_;
  assign FpAlu_8U_23U_mux1h_153_nl = _2428_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16413" *) _1126_;
  assign _2429_ = _1127_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16430" *) _1128_;
  assign _2430_ = _2429_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16431" *) _1129_;
  assign _2431_ = _2430_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16432" *) _1130_;
  assign _2432_ = _2431_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16433" *) _1131_;
  assign _2433_ = _2432_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16434" *) _1132_;
  assign _2434_ = _2433_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16435" *) _1133_;
  assign FpAlu_8U_23U_mux1h_34_nl = _2434_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16436" *) _1134_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_8U_23U_4_nor_3_itm_2 <= 1'b0;
    else
      IsNaN_8U_23U_4_nor_3_itm_2 <= _0218_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_8U_23U_2_IsNaN_8U_23U_2_nor_itm <= 1'b0;
    else
      IsNaN_8U_23U_2_IsNaN_8U_23U_2_nor_itm <= _0215_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_8U_23U_2_IsNaN_8U_23U_2_nor_1_itm <= 1'b0;
    else
      IsNaN_8U_23U_2_IsNaN_8U_23U_2_nor_1_itm <= _0209_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_8U_23U_2_IsNaN_8U_23U_2_nor_2_itm <= 1'b0;
    else
      IsNaN_8U_23U_2_IsNaN_8U_23U_2_nor_2_itm <= _0211_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_8U_23U_2_IsNaN_8U_23U_2_nor_3_itm <= 1'b0;
    else
      IsNaN_8U_23U_2_IsNaN_8U_23U_2_nor_3_itm <= _0213_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_8U_23U_4_nor_2_itm_2 <= 1'b0;
    else
      IsNaN_8U_23U_4_nor_2_itm_2 <= _0217_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_8U_23U_4_nor_3_itm_3 <= 1'b0;
    else
      IsNaN_8U_23U_4_nor_3_itm_3 <= _0219_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpCmp_8U_23U_false_is_abs_a_greater_2_lpi_1_dfm_2 <= 1'b0;
    else
      FpCmp_8U_23U_false_is_abs_a_greater_2_lpi_1_dfm_2 <= _0157_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_8U_23U_2_IsNaN_8U_23U_2_nor_1_itm_1 <= 1'b0;
    else
      IsNaN_8U_23U_2_IsNaN_8U_23U_2_nor_1_itm_1 <= _0210_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_8U_23U_2_IsNaN_8U_23U_2_nor_2_itm_1 <= 1'b0;
    else
      IsNaN_8U_23U_2_IsNaN_8U_23U_2_nor_2_itm_1 <= _0212_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_8U_23U_2_IsNaN_8U_23U_2_nor_itm_2 <= 1'b0;
    else
      IsNaN_8U_23U_2_IsNaN_8U_23U_2_nor_itm_2 <= _0216_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_8U_23U_2_IsNaN_8U_23U_2_nor_3_itm_2 <= 1'b0;
    else
      IsNaN_8U_23U_2_IsNaN_8U_23U_2_nor_3_itm_2 <= _0214_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      alu_loop_op_2_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_1_svs_2 <= 1'b0;
    else
      alu_loop_op_2_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_1_svs_2 <= _0266_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpAlu_8U_23U_mux1h_33_itm_2 <= 1'b0;
    else
      FpAlu_8U_23U_mux1h_33_itm_2 <= _0147_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpAlu_8U_23U_mux1h_152_itm_2 <= 1'b0;
    else
      FpAlu_8U_23U_mux1h_152_itm_2 <= _0146_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      alu_loop_op_3_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_svs_2 <= 1'b0;
    else
      alu_loop_op_3_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_svs_2 <= _0280_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      alu_loop_op_1_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_svs_2 <= 1'b0;
    else
      alu_loop_op_1_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_svs_2 <= _0254_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      alu_loop_op_4_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_1_svs_2 <= 1'b0;
    else
      alu_loop_op_4_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_1_svs_2 <= _0293_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      reg_alu_loop_op_else_o_32_1_lpi_1_dfm_4_1_itm <= 31'b0000000000000000000000000000000;
    else
      reg_alu_loop_op_else_o_32_1_lpi_1_dfm_4_1_itm <= _0385_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      reg_alu_loop_op_else_o_32_1_lpi_1_dfm_4_itm <= 1'b0;
    else
      reg_alu_loop_op_else_o_32_1_lpi_1_dfm_4_itm <= _0386_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      reg_alu_loop_op_else_o_32_1_3_lpi_1_dfm_3_1_itm <= 31'b0000000000000000000000000000000;
    else
      reg_alu_loop_op_else_o_32_1_3_lpi_1_dfm_3_1_itm <= _0383_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      reg_alu_loop_op_else_o_32_1_3_lpi_1_dfm_3_itm <= 1'b0;
    else
      reg_alu_loop_op_else_o_32_1_3_lpi_1_dfm_3_itm <= _0384_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      alu_loop_op_2_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_1_svs_3 <= 1'b0;
    else
      alu_loop_op_2_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_1_svs_3 <= _0267_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      reg_alu_loop_op_else_o_32_1_2_lpi_1_dfm_4_1_itm <= 31'b0000000000000000000000000000000;
    else
      reg_alu_loop_op_else_o_32_1_2_lpi_1_dfm_4_1_itm <= _0381_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      reg_alu_loop_op_else_o_32_1_2_lpi_1_dfm_4_itm <= 1'b0;
    else
      reg_alu_loop_op_else_o_32_1_2_lpi_1_dfm_4_itm <= _0382_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      reg_alu_loop_op_else_o_32_1_1_lpi_1_dfm_3_1_itm <= 31'b0000000000000000000000000000000;
    else
      reg_alu_loop_op_else_o_32_1_1_lpi_1_dfm_3_1_itm <= _0379_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      reg_alu_loop_op_else_o_32_1_1_lpi_1_dfm_3_itm <= 1'b0;
    else
      reg_alu_loop_op_else_o_32_1_1_lpi_1_dfm_3_itm <= _0380_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpAlu_8U_23U_equal_tmp_33 <= 1'b0;
    else
      FpAlu_8U_23U_equal_tmp_33 <= _0143_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpAlu_8U_23U_equal_tmp_30 <= 1'b0;
    else
      FpAlu_8U_23U_equal_tmp_30 <= _0140_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpCmp_8U_23U_true_o_3_lpi_1_dfm_5_30_0_1 <= 31'b0000000000000000000000000000000;
    else
      FpCmp_8U_23U_true_o_3_lpi_1_dfm_5_30_0_1 <= _0172_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpCmp_8U_23U_true_o_2_lpi_1_dfm_5_30_0_1 <= 31'b0000000000000000000000000000000;
    else
      FpCmp_8U_23U_true_o_2_lpi_1_dfm_5_30_0_1 <= _0169_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpCmp_8U_23U_true_o_1_lpi_1_dfm_5_30_0_1 <= 31'b0000000000000000000000000000000;
    else
      FpCmp_8U_23U_true_o_1_lpi_1_dfm_5_30_0_1 <= _0166_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpCmp_8U_23U_true_o_lpi_1_dfm_5_30_0_1 <= 31'b0000000000000000000000000000000;
    else
      FpCmp_8U_23U_true_o_lpi_1_dfm_5_30_0_1 <= _0175_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      AluOut_data_1_0_sva_10 <= 1'b0;
    else
      AluOut_data_1_0_sva_10 <= _0066_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      AluOut_data_0_0_sva_9 <= 1'b0;
    else
      AluOut_data_0_0_sva_9 <= _0065_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      AluOut_data_2_0_sva_9 <= 1'b0;
    else
      AluOut_data_2_0_sva_9 <= _0072_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpAlu_8U_23U_o_0_sva_7 <= 1'b0;
    else
      FpAlu_8U_23U_o_0_sva_7 <= _0152_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_8U_23U_land_lpi_1_dfm_9 <= 1'b0;
    else
      IsNaN_8U_23U_land_lpi_1_dfm_9 <= _0241_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_8U_23U_land_3_lpi_1_dfm_9 <= 1'b0;
    else
      IsNaN_8U_23U_land_3_lpi_1_dfm_9 <= _0235_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_8U_23U_land_2_lpi_1_dfm_9 <= 1'b0;
    else
      IsNaN_8U_23U_land_2_lpi_1_dfm_9 <= _0229_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_8U_23U_land_1_lpi_1_dfm_9 <= 1'b0;
    else
      IsNaN_8U_23U_land_1_lpi_1_dfm_9 <= _0223_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      alu_loop_op_2_FpAdd_8U_23U_IsZero_8U_23U_or_itm_3 <= 1'b0;
    else
      alu_loop_op_2_FpAdd_8U_23U_IsZero_8U_23U_or_itm_3 <= _0257_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      alu_loop_op_3_FpAdd_8U_23U_IsZero_8U_23U_or_itm_3 <= 1'b0;
    else
      alu_loop_op_3_FpAdd_8U_23U_IsZero_8U_23U_or_itm_3 <= _0270_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      alu_loop_op_4_FpAdd_8U_23U_IsZero_8U_23U_or_itm_3 <= 1'b0;
    else
      alu_loop_op_4_FpAdd_8U_23U_IsZero_8U_23U_or_itm_3 <= _0283_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpAdd_8U_23U_qr_lpi_1_dfm <= 8'b00000000;
    else
      FpAdd_8U_23U_qr_lpi_1_dfm <= _0126_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpAdd_8U_23U_qr_4_lpi_1_dfm <= 8'b00000000;
    else
      FpAdd_8U_23U_qr_4_lpi_1_dfm <= _0123_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpAdd_8U_23U_qr_3_lpi_1_dfm <= 8'b00000000;
    else
      FpAdd_8U_23U_qr_3_lpi_1_dfm <= _0120_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpAdd_8U_23U_qr_2_lpi_1_dfm <= 8'b00000000;
    else
      FpAdd_8U_23U_qr_2_lpi_1_dfm <= _0117_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpAlu_8U_23U_equal_tmp_21 <= 1'b0;
    else
      FpAlu_8U_23U_equal_tmp_21 <= _0131_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpAlu_8U_23U_equal_tmp_24 <= 1'b0;
    else
      FpAlu_8U_23U_equal_tmp_24 <= _0134_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpAlu_8U_23U_nor_dfs_4 <= 1'b0;
    else
      FpAlu_8U_23U_nor_dfs_4 <= _0148_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpAlu_8U_23U_equal_tmp_27 <= 1'b0;
    else
      FpAlu_8U_23U_equal_tmp_27 <= _0137_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpAlu_8U_23U_and_6_itm_2 <= 1'b0;
    else
      FpAlu_8U_23U_and_6_itm_2 <= _0130_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpAlu_8U_23U_and_3_itm_2 <= 1'b0;
    else
      FpAlu_8U_23U_and_3_itm_2 <= _0129_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      else_AluOp_data_slc_else_AluOp_data_3_30_23_35_itm <= 8'b00000000;
    else
      else_AluOp_data_slc_else_AluOp_data_3_30_23_35_itm <= _0347_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      else_AluOp_data_slc_else_AluOp_data_0_30_23_7_itm <= 8'b00000000;
    else
      else_AluOp_data_slc_else_AluOp_data_0_30_23_7_itm <= _0335_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      else_AluOp_data_slc_else_AluOp_data_1_30_23_21_itm <= 8'b00000000;
    else
      else_AluOp_data_slc_else_AluOp_data_1_30_23_21_itm <= _0339_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      else_AluOp_data_slc_else_AluOp_data_2_30_23_21_itm <= 8'b00000000;
    else
      else_AluOp_data_slc_else_AluOp_data_2_30_23_21_itm <= _0343_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      else_AluOp_data_slc_else_AluOp_data_3_22_0_12_itm <= 23'b00000000000000000000000;
    else
      else_AluOp_data_slc_else_AluOp_data_3_22_0_12_itm <= _0345_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      else_AluOp_data_slc_else_AluOp_data_2_22_0_7_itm <= 23'b00000000000000000000000;
    else
      else_AluOp_data_slc_else_AluOp_data_2_22_0_7_itm <= _0341_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      else_AluOp_data_slc_else_AluOp_data_1_22_0_7_itm <= 23'b00000000000000000000000;
    else
      else_AluOp_data_slc_else_AluOp_data_1_22_0_7_itm <= _0337_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      else_AluOp_data_slc_else_AluOp_data_0_22_0_2_itm <= 23'b00000000000000000000000;
    else
      else_AluOp_data_slc_else_AluOp_data_0_22_0_2_itm <= _0333_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      else_AluOp_data_slc_else_AluOp_data_3_22_0_12_itm_2 <= 23'b00000000000000000000000;
    else
      else_AluOp_data_slc_else_AluOp_data_3_22_0_12_itm_2 <= _0346_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      else_AluOp_data_slc_else_AluOp_data_2_22_0_7_itm_2 <= 23'b00000000000000000000000;
    else
      else_AluOp_data_slc_else_AluOp_data_2_22_0_7_itm_2 <= _0342_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      else_AluOp_data_slc_else_AluOp_data_1_22_0_7_itm_2 <= 23'b00000000000000000000000;
    else
      else_AluOp_data_slc_else_AluOp_data_1_22_0_7_itm_2 <= _0338_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      else_AluOp_data_slc_else_AluOp_data_0_22_0_2_itm_2 <= 23'b00000000000000000000000;
    else
      else_AluOp_data_slc_else_AluOp_data_0_22_0_2_itm_2 <= _0334_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      AluOut_data_2_31_lpi_1_dfm_6 <= 1'b0;
    else
      AluOut_data_2_31_lpi_1_dfm_6 <= _0075_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      mux_189_itm_3 <= 1'b0;
    else
      mux_189_itm_3 <= _0365_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      mux_181_itm_3 <= 1'b0;
    else
      mux_181_itm_3 <= _0363_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      mux_177_itm_3 <= 1'b0;
    else
      mux_177_itm_3 <= _0361_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntSaturation_33U_32U_slc_IntSaturation_33U_32U_o_31_1_1_29_22_itm_2 <= 8'b00000000;
    else
      IntSaturation_33U_32U_slc_IntSaturation_33U_32U_o_31_1_1_29_22_itm_2 <= _0187_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntSaturation_33U_32U_slc_IntSaturation_33U_32U_o_31_1_2_29_22_itm_3 <= 8'b00000000;
    else
      IntSaturation_33U_32U_slc_IntSaturation_33U_32U_o_31_1_2_29_22_itm_3 <= _0193_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntSaturation_33U_32U_slc_IntSaturation_33U_32U_o_31_1_29_22_itm_3 <= 8'b00000000;
    else
      IntSaturation_33U_32U_slc_IntSaturation_33U_32U_o_31_1_29_22_itm_3 <= _0190_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntSaturation_33U_32U_slc_IntSaturation_33U_32U_o_31_1_3_21_0_itm_3 <= 22'b0000000000000000000000;
    else
      IntSaturation_33U_32U_slc_IntSaturation_33U_32U_o_31_1_3_21_0_itm_3 <= _0194_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntSaturation_33U_32U_slc_IntSaturation_33U_32U_o_31_1_21_0_itm_3 <= 22'b0000000000000000000000;
    else
      IntSaturation_33U_32U_slc_IntSaturation_33U_32U_o_31_1_21_0_itm_3 <= _0188_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntSaturation_33U_32U_slc_IntSaturation_33U_32U_o_31_1_2_21_0_itm_3 <= 22'b0000000000000000000000;
    else
      IntSaturation_33U_32U_slc_IntSaturation_33U_32U_o_31_1_2_21_0_itm_3 <= _0191_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntSaturation_33U_32U_slc_IntSaturation_33U_32U_o_31_1_1_21_0_itm_2 <= 22'b0000000000000000000000;
    else
      IntSaturation_33U_32U_slc_IntSaturation_33U_32U_o_31_1_1_21_0_itm_2 <= _0186_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntSaturation_33U_32U_slc_IntSaturation_33U_32U_o_31_1_3_29_22_itm_3 <= 8'b00000000;
    else
      IntSaturation_33U_32U_slc_IntSaturation_33U_32U_o_31_1_3_29_22_itm_3 <= _0196_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpAlu_8U_23U_equal_tmp_34 <= 1'b0;
    else
      FpAlu_8U_23U_equal_tmp_34 <= _0144_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpCmp_8U_23U_false_o_2_lpi_1_dfm_7_30_0_1 <= 31'b0000000000000000000000000000000;
    else
      FpCmp_8U_23U_false_o_2_lpi_1_dfm_7_30_0_1 <= _0160_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpCmp_8U_23U_false_o_1_lpi_1_dfm_6_30_0_1 <= 31'b0000000000000000000000000000000;
    else
      FpCmp_8U_23U_false_o_1_lpi_1_dfm_6_30_0_1 <= _0158_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpCmp_8U_23U_false_o_3_lpi_1_dfm_7_30_0_1 <= 31'b0000000000000000000000000000000;
    else
      FpCmp_8U_23U_false_o_3_lpi_1_dfm_7_30_0_1 <= _0162_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpCmp_8U_23U_false_o_lpi_1_dfm_8_30_0_1 <= 31'b0000000000000000000000000000000;
    else
      FpCmp_8U_23U_false_o_lpi_1_dfm_8_30_0_1 <= _0164_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpCmp_8U_23U_true_o_3_lpi_1_dfm_6_30_0_1 <= 31'b0000000000000000000000000000000;
    else
      FpCmp_8U_23U_true_o_3_lpi_1_dfm_6_30_0_1 <= _0173_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpCmp_8U_23U_true_o_2_lpi_1_dfm_6_30_0_1 <= 31'b0000000000000000000000000000000;
    else
      FpCmp_8U_23U_true_o_2_lpi_1_dfm_6_30_0_1 <= _0170_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpCmp_8U_23U_true_o_1_lpi_1_dfm_6_30_0_1 <= 31'b0000000000000000000000000000000;
    else
      FpCmp_8U_23U_true_o_1_lpi_1_dfm_6_30_0_1 <= _0167_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpCmp_8U_23U_true_o_lpi_1_dfm_6_30_0_1 <= 31'b0000000000000000000000000000000;
    else
      FpCmp_8U_23U_true_o_lpi_1_dfm_6_30_0_1 <= _0176_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpAlu_8U_23U_equal_tmp_22 <= 1'b0;
    else
      FpAlu_8U_23U_equal_tmp_22 <= _0132_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpAlu_8U_23U_equal_tmp_25 <= 1'b0;
    else
      FpAlu_8U_23U_equal_tmp_25 <= _0135_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpAlu_8U_23U_nor_dfs_5 <= 1'b0;
    else
      FpAlu_8U_23U_nor_dfs_5 <= _0149_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpAlu_8U_23U_equal_tmp_28 <= 1'b0;
    else
      FpAlu_8U_23U_equal_tmp_28 <= _0138_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpAlu_8U_23U_equal_tmp_31 <= 1'b0;
    else
      FpAlu_8U_23U_equal_tmp_31 <= _0141_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      AluOut_data_2_0_sva_10 <= 1'b0;
    else
      AluOut_data_2_0_sva_10 <= _0070_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      AluOut_data_1_0_sva_11 <= 1'b0;
    else
      AluOut_data_1_0_sva_11 <= _0067_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      AluOut_data_0_0_sva_10 <= 1'b0;
    else
      AluOut_data_0_0_sva_10 <= _0063_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpAlu_8U_23U_o_0_sva_8 <= 1'b0;
    else
      FpAlu_8U_23U_o_0_sva_8 <= _0153_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_8U_23U_land_lpi_1_dfm_10 <= 1'b0;
    else
      IsNaN_8U_23U_land_lpi_1_dfm_10 <= _0238_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_8U_23U_land_3_lpi_1_dfm_10 <= 1'b0;
    else
      IsNaN_8U_23U_land_3_lpi_1_dfm_10 <= _0232_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_8U_23U_land_2_lpi_1_dfm_10 <= 1'b0;
    else
      IsNaN_8U_23U_land_2_lpi_1_dfm_10 <= _0226_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_8U_23U_land_1_lpi_1_dfm_10 <= 1'b0;
    else
      IsNaN_8U_23U_land_1_lpi_1_dfm_10 <= _0220_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpAdd_8U_23U_qr_lpi_1_dfm_6 <= 8'b00000000;
    else
      FpAdd_8U_23U_qr_lpi_1_dfm_6 <= _0127_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpAdd_8U_23U_qr_4_lpi_1_dfm_6 <= 8'b00000000;
    else
      FpAdd_8U_23U_qr_4_lpi_1_dfm_6 <= _0124_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpAdd_8U_23U_qr_3_lpi_1_dfm_6 <= 8'b00000000;
    else
      FpAdd_8U_23U_qr_3_lpi_1_dfm_6 <= _0121_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpAdd_8U_23U_qr_2_lpi_1_dfm_6 <= 8'b00000000;
    else
      FpAdd_8U_23U_qr_2_lpi_1_dfm_6 <= _0118_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cfg_alu_algo_1_sva_2 <= 2'b00;
    else
      cfg_alu_algo_1_sva_2 <= _0297_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cfg_alu_src_1_sva_st <= 1'b0;
    else
      cfg_alu_src_1_sva_st <= _0306_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cfg_alu_algo_1_sva_st <= 2'b00;
    else
      cfg_alu_algo_1_sva_st <= _0298_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cfg_alu_algo_1_sva_st_20 <= 2'b00;
    else
      cfg_alu_algo_1_sva_st_20 <= _0299_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      alu_loop_op_1_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_st <= 1'b0;
    else
      alu_loop_op_1_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_st <= _0249_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      alu_loop_op_2_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_2_svs_st <= 1'b0;
    else
      alu_loop_op_2_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_2_svs_st <= _0261_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      alu_loop_op_3_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_1_svs_st <= 1'b0;
    else
      alu_loop_op_3_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_1_svs_st <= _0275_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      alu_loop_op_4_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_3_svs_st <= 1'b0;
    else
      alu_loop_op_4_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_3_svs_st <= _0288_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpAdd_8U_23U_b_right_shift_qr_lpi_1_dfm <= 8'b00000000;
    else
      FpAdd_8U_23U_b_right_shift_qr_lpi_1_dfm <= _0095_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpAdd_8U_23U_a_right_shift_qr_lpi_1_dfm <= 8'b00000000;
    else
      FpAdd_8U_23U_a_right_shift_qr_lpi_1_dfm <= _0083_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpAdd_8U_23U_b_right_shift_qr_1_lpi_1_dfm <= 8'b00000000;
    else
      FpAdd_8U_23U_b_right_shift_qr_1_lpi_1_dfm <= _0089_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpAdd_8U_23U_a_right_shift_qr_1_lpi_1_dfm <= 8'b00000000;
    else
      FpAdd_8U_23U_a_right_shift_qr_1_lpi_1_dfm <= _0077_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpAdd_8U_23U_b_right_shift_qr_2_lpi_1_dfm <= 8'b00000000;
    else
      FpAdd_8U_23U_b_right_shift_qr_2_lpi_1_dfm <= _0091_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpAdd_8U_23U_a_right_shift_qr_2_lpi_1_dfm <= 8'b00000000;
    else
      FpAdd_8U_23U_a_right_shift_qr_2_lpi_1_dfm <= _0079_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpAdd_8U_23U_b_right_shift_qr_3_lpi_1_dfm <= 8'b00000000;
    else
      FpAdd_8U_23U_b_right_shift_qr_3_lpi_1_dfm <= _0093_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpAdd_8U_23U_a_right_shift_qr_3_lpi_1_dfm <= 8'b00000000;
    else
      FpAdd_8U_23U_a_right_shift_qr_3_lpi_1_dfm <= _0081_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      alu_loop_op_1_FpAdd_8U_23U_IsZero_8U_23U_1_or_itm <= 1'b0;
    else
      alu_loop_op_1_FpAdd_8U_23U_IsZero_8U_23U_1_or_itm <= _0244_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      alu_loop_op_2_FpAdd_8U_23U_IsZero_8U_23U_1_or_itm <= 1'b0;
    else
      alu_loop_op_2_FpAdd_8U_23U_IsZero_8U_23U_1_or_itm <= _0255_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      alu_loop_op_3_FpAdd_8U_23U_IsZero_8U_23U_1_or_itm <= 1'b0;
    else
      alu_loop_op_3_FpAdd_8U_23U_IsZero_8U_23U_1_or_itm <= _0268_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      alu_loop_op_4_FpAdd_8U_23U_IsZero_8U_23U_1_or_itm <= 1'b0;
    else
      alu_loop_op_4_FpAdd_8U_23U_IsZero_8U_23U_1_or_itm <= _0281_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      alu_loop_op_3_FpAdd_8U_23U_IsZero_8U_23U_or_itm_4 <= 1'b0;
    else
      alu_loop_op_3_FpAdd_8U_23U_IsZero_8U_23U_or_itm_4 <= _0271_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      alu_loop_op_4_FpAdd_8U_23U_IsZero_8U_23U_or_itm_4 <= 1'b0;
    else
      alu_loop_op_4_FpAdd_8U_23U_IsZero_8U_23U_or_itm_4 <= _0284_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      alu_loop_op_1_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_itm <= 1'b0;
    else
      alu_loop_op_1_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_itm <= _0250_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      alu_loop_op_2_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_2_itm <= 1'b0;
    else
      alu_loop_op_2_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_2_itm <= _0262_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      alu_loop_op_3_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_1_itm <= 1'b0;
    else
      alu_loop_op_3_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_1_itm <= _0276_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      alu_loop_op_4_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_3_itm <= 1'b0;
    else
      alu_loop_op_4_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_3_itm <= _0289_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpNormalize_8U_49U_if_or_3_itm <= 1'b0;
    else
      FpNormalize_8U_49U_if_or_3_itm <= _0182_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpNormalize_8U_49U_if_or_2_itm <= 1'b0;
    else
      FpNormalize_8U_49U_if_or_2_itm <= _0180_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpNormalize_8U_49U_if_or_1_itm <= 1'b0;
    else
      FpNormalize_8U_49U_if_or_1_itm <= _0178_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpAdd_8U_23U_int_mant_p1_1_lpi_1_dfm <= 50'b00000000000000000000000000000000000000000000000000;
    else
      FpAdd_8U_23U_int_mant_p1_1_lpi_1_dfm <= _0097_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpAdd_8U_23U_int_mant_p1_2_lpi_1_dfm <= 50'b00000000000000000000000000000000000000000000000000;
    else
      FpAdd_8U_23U_int_mant_p1_2_lpi_1_dfm <= _0099_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpAdd_8U_23U_int_mant_p1_3_lpi_1_dfm <= 50'b00000000000000000000000000000000000000000000000000;
    else
      FpAdd_8U_23U_int_mant_p1_3_lpi_1_dfm <= _0101_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpAdd_8U_23U_int_mant_p1_lpi_1_dfm <= 50'b00000000000000000000000000000000000000000000000000;
    else
      FpAdd_8U_23U_int_mant_p1_lpi_1_dfm <= _0103_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpNormalize_8U_49U_if_or_itm <= 1'b0;
    else
      FpNormalize_8U_49U_if_or_itm <= _0184_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_8U_23U_1_land_lpi_1_dfm_8 <= 1'b0;
    else
      IsNaN_8U_23U_1_land_lpi_1_dfm_8 <= _0207_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_8U_23U_1_land_3_lpi_1_dfm_8 <= 1'b0;
    else
      IsNaN_8U_23U_1_land_3_lpi_1_dfm_8 <= _0204_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_8U_23U_1_land_2_lpi_1_dfm_8 <= 1'b0;
    else
      IsNaN_8U_23U_1_land_2_lpi_1_dfm_8 <= _0201_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_8U_23U_1_land_1_lpi_1_dfm_8 <= 1'b0;
    else
      IsNaN_8U_23U_1_land_1_lpi_1_dfm_8 <= _0198_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      alu_loop_op_1_FpMantRNE_49U_24U_else_and_svs_st <= 1'b0;
    else
      alu_loop_op_1_FpMantRNE_49U_24U_else_and_svs_st <= _0252_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      alu_loop_op_2_FpMantRNE_49U_24U_else_and_2_svs_st <= 1'b0;
    else
      alu_loop_op_2_FpMantRNE_49U_24U_else_and_2_svs_st <= _0264_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      alu_loop_op_3_FpMantRNE_49U_24U_else_and_1_svs_st <= 1'b0;
    else
      alu_loop_op_3_FpMantRNE_49U_24U_else_and_1_svs_st <= _0278_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      alu_loop_op_4_FpMantRNE_49U_24U_else_and_3_svs_st <= 1'b0;
    else
      alu_loop_op_4_FpMantRNE_49U_24U_else_and_3_svs_st <= _0291_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      alu_loop_op_4_FpAdd_8U_23U_if_4_if_slc_FpAdd_8U_23U_if_4_if_acc_1_7_3_svs_st_2 <= 1'b0;
    else
      alu_loop_op_4_FpAdd_8U_23U_if_4_if_slc_FpAdd_8U_23U_if_4_if_acc_1_7_3_svs_st_2 <= _0286_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      alu_loop_op_3_FpAdd_8U_23U_if_4_if_slc_FpAdd_8U_23U_if_4_if_acc_1_7_1_svs_st_2 <= 1'b0;
    else
      alu_loop_op_3_FpAdd_8U_23U_if_4_if_slc_FpAdd_8U_23U_if_4_if_acc_1_7_1_svs_st_2 <= _0273_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      alu_loop_op_2_FpAdd_8U_23U_if_4_if_slc_FpAdd_8U_23U_if_4_if_acc_1_7_2_svs_st_2 <= 1'b0;
    else
      alu_loop_op_2_FpAdd_8U_23U_if_4_if_slc_FpAdd_8U_23U_if_4_if_acc_1_7_2_svs_st_2 <= _0259_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      alu_loop_op_1_FpAdd_8U_23U_if_4_if_slc_FpAdd_8U_23U_if_4_if_acc_1_7_svs_st_2 <= 1'b0;
    else
      alu_loop_op_1_FpAdd_8U_23U_if_4_if_slc_FpAdd_8U_23U_if_4_if_acc_1_7_svs_st_2 <= _0247_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      AluOut_data_2_0_sva_11 <= 1'b0;
    else
      AluOut_data_2_0_sva_11 <= _0071_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      AluOut_data_2_0_lpi_1_dfm_3 <= 1'b0;
    else
      AluOut_data_2_0_lpi_1_dfm_3 <= _0069_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntSaturation_33U_32U_slc_IntSaturation_33U_32U_o_31_1_3_21_0_itm_4 <= 22'b0000000000000000000000;
    else
      IntSaturation_33U_32U_slc_IntSaturation_33U_32U_o_31_1_3_21_0_itm_4 <= _0195_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntSaturation_33U_32U_slc_IntSaturation_33U_32U_o_31_1_21_0_itm_4 <= 22'b0000000000000000000000;
    else
      IntSaturation_33U_32U_slc_IntSaturation_33U_32U_o_31_1_21_0_itm_4 <= _0189_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntSaturation_33U_32U_slc_IntSaturation_33U_32U_o_31_1_2_21_0_itm_4 <= 22'b0000000000000000000000;
    else
      IntSaturation_33U_32U_slc_IntSaturation_33U_32U_o_31_1_2_21_0_itm_4 <= _0192_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      AluOut_data_1_0_sva_12 <= 1'b0;
    else
      AluOut_data_1_0_sva_12 <= _0068_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      AluOut_data_0_0_sva_11 <= 1'b0;
    else
      AluOut_data_0_0_sva_11 <= _0064_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      alu_loop_op_unequal_tmp_8 <= 1'b0;
    else
      alu_loop_op_unequal_tmp_8 <= _0296_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      io_read_cfg_alu_bypass_rsc_svs_8 <= 1'b0;
    else
      io_read_cfg_alu_bypass_rsc_svs_8 <= _0352_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      AluOut_data_2_31_lpi_1_dfm_7 <= 1'b0;
    else
      AluOut_data_2_31_lpi_1_dfm_7 <= _0076_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      mux_189_itm_4 <= 1'b0;
    else
      mux_189_itm_4 <= _0366_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      mux_181_itm_4 <= 1'b0;
    else
      mux_181_itm_4 <= _0364_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      mux_177_itm_4 <= 1'b0;
    else
      mux_177_itm_4 <= _0362_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      io_read_cfg_alu_bypass_rsc_svs_st_7 <= 1'b0;
    else
      io_read_cfg_alu_bypass_rsc_svs_st_7 <= _0356_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cfg_alu_algo_1_sva_st_25 <= 2'b00;
    else
      cfg_alu_algo_1_sva_st_25 <= _0303_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpAlu_8U_23U_equal_tmp_35 <= 1'b0;
    else
      FpAlu_8U_23U_equal_tmp_35 <= _0145_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      else_AluOp_data_slc_else_AluOp_data_3_30_23_35_itm_3 <= 8'b00000000;
    else
      else_AluOp_data_slc_else_AluOp_data_3_30_23_35_itm_3 <= _0348_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpAdd_8U_23U_is_inf_lpi_1_dfm_8 <= 1'b0;
    else
      FpAdd_8U_23U_is_inf_lpi_1_dfm_8 <= _0112_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpAlu_8U_23U_o_30_23_lpi_1_dfm_4 <= 8'b00000000;
    else
      FpAlu_8U_23U_o_30_23_lpi_1_dfm_4 <= _0156_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpAlu_8U_23U_o_22_1_lpi_1_dfm_4 <= 22'b0000000000000000000000;
    else
      FpAlu_8U_23U_o_22_1_lpi_1_dfm_4 <= _0155_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpCmp_8U_23U_false_o_lpi_1_dfm_9_30_0_1 <= 31'b0000000000000000000000000000000;
    else
      FpCmp_8U_23U_false_o_lpi_1_dfm_9_30_0_1 <= _0165_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpAlu_8U_23U_o_0_lpi_1_dfm_4 <= 1'b0;
    else
      FpAlu_8U_23U_o_0_lpi_1_dfm_4 <= _0151_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpAlu_8U_23U_o_0_sva_9 <= 1'b0;
    else
      FpAlu_8U_23U_o_0_sva_9 <= _0154_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpCmp_8U_23U_true_o_lpi_1_dfm_7_30_0_1 <= 31'b0000000000000000000000000000000;
    else
      FpCmp_8U_23U_true_o_lpi_1_dfm_7_30_0_1 <= _0177_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      else_AluOp_data_slc_else_AluOp_data_0_30_23_7_itm_3 <= 8'b00000000;
    else
      else_AluOp_data_slc_else_AluOp_data_0_30_23_7_itm_3 <= _0336_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpAdd_8U_23U_is_inf_1_lpi_1_dfm_8 <= 1'b0;
    else
      FpAdd_8U_23U_is_inf_1_lpi_1_dfm_8 <= _0109_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      else_AluOp_data_slc_else_AluOp_data_1_30_23_21_itm_3 <= 8'b00000000;
    else
      else_AluOp_data_slc_else_AluOp_data_1_30_23_21_itm_3 <= _0340_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpAdd_8U_23U_is_inf_2_lpi_1_dfm_8 <= 1'b0;
    else
      FpAdd_8U_23U_is_inf_2_lpi_1_dfm_8 <= _0110_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpCmp_8U_23U_false_o_2_lpi_1_dfm_8_30_0_1 <= 31'b0000000000000000000000000000000;
    else
      FpCmp_8U_23U_false_o_2_lpi_1_dfm_8_30_0_1 <= _0161_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpCmp_8U_23U_false_o_1_lpi_1_dfm_7_30_0_1 <= 31'b0000000000000000000000000000000;
    else
      FpCmp_8U_23U_false_o_1_lpi_1_dfm_7_30_0_1 <= _0159_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      AluOut_data_2_30_23_lpi_1_dfm_3 <= 8'b00000000;
    else
      AluOut_data_2_30_23_lpi_1_dfm_3 <= _0074_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      else_AluOp_data_slc_else_AluOp_data_2_30_23_21_itm_3 <= 8'b00000000;
    else
      else_AluOp_data_slc_else_AluOp_data_2_30_23_21_itm_3 <= _0344_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpAdd_8U_23U_is_inf_3_lpi_1_dfm_8 <= 1'b0;
    else
      FpAdd_8U_23U_is_inf_3_lpi_1_dfm_8 <= _0111_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpCmp_8U_23U_false_o_3_lpi_1_dfm_8_30_0_1 <= 31'b0000000000000000000000000000000;
    else
      FpCmp_8U_23U_false_o_3_lpi_1_dfm_8_30_0_1 <= _0163_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      AluOut_data_2_22_1_lpi_1_dfm_3 <= 22'b0000000000000000000000;
    else
      AluOut_data_2_22_1_lpi_1_dfm_3 <= _0073_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpCmp_8U_23U_true_o_3_lpi_1_dfm_7_30_0_1 <= 31'b0000000000000000000000000000000;
    else
      FpCmp_8U_23U_true_o_3_lpi_1_dfm_7_30_0_1 <= _0174_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpCmp_8U_23U_true_o_2_lpi_1_dfm_7_30_0_1 <= 31'b0000000000000000000000000000000;
    else
      FpCmp_8U_23U_true_o_2_lpi_1_dfm_7_30_0_1 <= _0171_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpCmp_8U_23U_true_o_1_lpi_1_dfm_7_30_0_1 <= 31'b0000000000000000000000000000000;
    else
      FpCmp_8U_23U_true_o_1_lpi_1_dfm_7_30_0_1 <= _0168_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpAlu_8U_23U_equal_tmp_23 <= 1'b0;
    else
      FpAlu_8U_23U_equal_tmp_23 <= _0133_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpAlu_8U_23U_equal_tmp_26 <= 1'b0;
    else
      FpAlu_8U_23U_equal_tmp_26 <= _0136_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpAlu_8U_23U_nor_dfs_6 <= 1'b0;
    else
      FpAlu_8U_23U_nor_dfs_6 <= _0150_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpAlu_8U_23U_equal_tmp_29 <= 1'b0;
    else
      FpAlu_8U_23U_equal_tmp_29 <= _0139_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpAlu_8U_23U_equal_tmp_32 <= 1'b0;
    else
      FpAlu_8U_23U_equal_tmp_32 <= _0142_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      reg_AluIn_data_sva_4_30_0_1_itm <= 23'b00000000000000000000000;
    else
      reg_AluIn_data_sva_4_30_0_1_itm <= _0369_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      reg_AluIn_data_sva_4_30_0_itm <= 8'b00000000;
    else
      reg_AluIn_data_sva_4_30_0_itm <= _0370_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      reg_AluIn_data_sva_4_62_32_1_itm <= 23'b00000000000000000000000;
    else
      reg_AluIn_data_sva_4_62_32_1_itm <= _0371_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      reg_AluIn_data_sva_4_62_32_itm <= 8'b00000000;
    else
      reg_AluIn_data_sva_4_62_32_itm <= _0372_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      reg_AluIn_data_sva_4_94_64_1_itm <= 23'b00000000000000000000000;
    else
      reg_AluIn_data_sva_4_94_64_1_itm <= _0373_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      reg_AluIn_data_sva_4_94_64_itm <= 8'b00000000;
    else
      reg_AluIn_data_sva_4_94_64_itm <= _0374_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      alu_loop_op_1_FpMantRNE_49U_24U_else_and_svs_st_2 <= 1'b0;
    else
      alu_loop_op_1_FpMantRNE_49U_24U_else_and_svs_st_2 <= _0253_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      alu_loop_op_2_FpMantRNE_49U_24U_else_and_2_svs_st_2 <= 1'b0;
    else
      alu_loop_op_2_FpMantRNE_49U_24U_else_and_2_svs_st_2 <= _0265_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      alu_loop_op_3_FpMantRNE_49U_24U_else_and_1_svs_st_2 <= 1'b0;
    else
      alu_loop_op_3_FpMantRNE_49U_24U_else_and_1_svs_st_2 <= _0279_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      alu_loop_op_4_FpMantRNE_49U_24U_else_and_3_svs_st_2 <= 1'b0;
    else
      alu_loop_op_4_FpMantRNE_49U_24U_else_and_3_svs_st_2 <= _0292_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_8U_23U_1_land_1_lpi_1_dfm_9 <= 1'b0;
    else
      IsNaN_8U_23U_1_land_1_lpi_1_dfm_9 <= _0199_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_8U_23U_1_land_2_lpi_1_dfm_9 <= 1'b0;
    else
      IsNaN_8U_23U_1_land_2_lpi_1_dfm_9 <= _0202_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_8U_23U_1_land_3_lpi_1_dfm_9 <= 1'b0;
    else
      IsNaN_8U_23U_1_land_3_lpi_1_dfm_9 <= _0205_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_8U_23U_1_land_lpi_1_dfm_9 <= 1'b0;
    else
      IsNaN_8U_23U_1_land_lpi_1_dfm_9 <= _0208_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpAdd_8U_23U_and_2_tmp_3 <= 1'b0;
    else
      FpAdd_8U_23U_and_2_tmp_3 <= _0086_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpAdd_8U_23U_and_1_tmp_3 <= 1'b0;
    else
      FpAdd_8U_23U_and_1_tmp_3 <= _0085_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpAdd_8U_23U_and_tmp_2 <= 1'b0;
    else
      FpAdd_8U_23U_and_tmp_2 <= _0088_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpAdd_8U_23U_and_3_tmp_3 <= 1'b0;
    else
      FpAdd_8U_23U_and_3_tmp_3 <= _0087_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_8U_23U_land_1_lpi_1_dfm_11 <= 1'b0;
    else
      IsNaN_8U_23U_land_1_lpi_1_dfm_11 <= _0221_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_8U_23U_land_2_lpi_1_dfm_11 <= 1'b0;
    else
      IsNaN_8U_23U_land_2_lpi_1_dfm_11 <= _0227_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_8U_23U_land_3_lpi_1_dfm_11 <= 1'b0;
    else
      IsNaN_8U_23U_land_3_lpi_1_dfm_11 <= _0233_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_8U_23U_land_lpi_1_dfm_11 <= 1'b0;
    else
      IsNaN_8U_23U_land_lpi_1_dfm_11 <= _0239_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      reg_AluIn_data_sva_4_126_96_1_itm <= 23'b00000000000000000000000;
    else
      reg_AluIn_data_sva_4_126_96_1_itm <= _0367_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      reg_AluIn_data_sva_4_126_96_itm <= 8'b00000000;
    else
      reg_AluIn_data_sva_4_126_96_itm <= _0368_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      alu_loop_op_4_FpAdd_8U_23U_if_4_if_slc_FpAdd_8U_23U_if_4_if_acc_1_7_3_svs_st_3 <= 1'b0;
    else
      alu_loop_op_4_FpAdd_8U_23U_if_4_if_slc_FpAdd_8U_23U_if_4_if_acc_1_7_3_svs_st_3 <= _0287_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      alu_loop_op_3_FpAdd_8U_23U_if_4_if_slc_FpAdd_8U_23U_if_4_if_acc_1_7_1_svs_st_3 <= 1'b0;
    else
      alu_loop_op_3_FpAdd_8U_23U_if_4_if_slc_FpAdd_8U_23U_if_4_if_acc_1_7_1_svs_st_3 <= _0274_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      alu_loop_op_2_FpAdd_8U_23U_if_4_if_slc_FpAdd_8U_23U_if_4_if_acc_1_7_2_svs_st_3 <= 1'b0;
    else
      alu_loop_op_2_FpAdd_8U_23U_if_4_if_slc_FpAdd_8U_23U_if_4_if_acc_1_7_2_svs_st_3 <= _0260_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      alu_loop_op_1_FpAdd_8U_23U_if_4_if_slc_FpAdd_8U_23U_if_4_if_acc_1_7_svs_st_3 <= 1'b0;
    else
      alu_loop_op_1_FpAdd_8U_23U_if_4_if_slc_FpAdd_8U_23U_if_4_if_acc_1_7_svs_st_3 <= _0248_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpAdd_8U_23U_o_expo_lpi_1_dfm_13 <= 8'b00000000;
    else
      FpAdd_8U_23U_o_expo_lpi_1_dfm_13 <= _0116_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpAdd_8U_23U_o_expo_3_lpi_1_dfm_13 <= 8'b00000000;
    else
      FpAdd_8U_23U_o_expo_3_lpi_1_dfm_13 <= _0115_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpAdd_8U_23U_o_expo_2_lpi_1_dfm_13 <= 8'b00000000;
    else
      FpAdd_8U_23U_o_expo_2_lpi_1_dfm_13 <= _0114_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpAdd_8U_23U_o_expo_1_lpi_1_dfm_13 <= 8'b00000000;
    else
      FpAdd_8U_23U_o_expo_1_lpi_1_dfm_13 <= _0113_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      main_stage_v_4 <= 1'b0;
    else
      main_stage_v_4 <= _0360_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      io_read_cfg_alu_bypass_rsc_svs_7 <= 1'b0;
    else
      io_read_cfg_alu_bypass_rsc_svs_7 <= _0351_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      io_read_cfg_alu_bypass_rsc_svs_st_6 <= 1'b0;
    else
      io_read_cfg_alu_bypass_rsc_svs_st_6 <= _0355_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      alu_loop_op_unequal_tmp_7 <= 1'b0;
    else
      alu_loop_op_unequal_tmp_7 <= _0295_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      AluIn_data_sva_3_126_96_1 <= 31'b0000000000000000000000000000000;
    else
      AluIn_data_sva_3_126_96_1 <= _0059_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      AluIn_data_sva_3_94_64_1 <= 31'b0000000000000000000000000000000;
    else
      AluIn_data_sva_3_94_64_1 <= _0062_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      AluIn_data_sva_3_62_32_1 <= 31'b0000000000000000000000000000000;
    else
      AluIn_data_sva_3_62_32_1 <= _0061_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      AluIn_data_sva_3_30_0_1 <= 31'b0000000000000000000000000000000;
    else
      AluIn_data_sva_3_30_0_1 <= _0060_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cfg_alu_algo_1_sva_st_24 <= 2'b00;
    else
      cfg_alu_algo_1_sva_st_24 <= _0302_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpNormalize_8U_49U_if_or_3_itm_2 <= 1'b0;
    else
      FpNormalize_8U_49U_if_or_3_itm_2 <= _0183_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpNormalize_8U_49U_if_or_2_itm_2 <= 1'b0;
    else
      FpNormalize_8U_49U_if_or_2_itm_2 <= _0181_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpNormalize_8U_49U_if_or_1_itm_2 <= 1'b0;
    else
      FpNormalize_8U_49U_if_or_1_itm_2 <= _0179_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpNormalize_8U_49U_if_or_itm_2 <= 1'b0;
    else
      FpNormalize_8U_49U_if_or_itm_2 <= _0185_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpAdd_8U_23U_int_mant_p1_1_lpi_1_dfm_5 <= 50'b00000000000000000000000000000000000000000000000000;
    else
      FpAdd_8U_23U_int_mant_p1_1_lpi_1_dfm_5 <= _0098_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpAdd_8U_23U_int_mant_p1_2_lpi_1_dfm_5 <= 50'b00000000000000000000000000000000000000000000000000;
    else
      FpAdd_8U_23U_int_mant_p1_2_lpi_1_dfm_5 <= _0100_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpAdd_8U_23U_int_mant_p1_3_lpi_1_dfm_5 <= 50'b00000000000000000000000000000000000000000000000000;
    else
      FpAdd_8U_23U_int_mant_p1_3_lpi_1_dfm_5 <= _0102_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpAdd_8U_23U_int_mant_p1_lpi_1_dfm_5 <= 50'b00000000000000000000000000000000000000000000000000;
    else
      FpAdd_8U_23U_int_mant_p1_lpi_1_dfm_5 <= _0104_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      alu_loop_op_1_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_itm_2 <= 1'b0;
    else
      alu_loop_op_1_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_itm_2 <= _0251_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      alu_loop_op_2_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_2_itm_2 <= 1'b0;
    else
      alu_loop_op_2_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_2_itm_2 <= _0263_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      alu_loop_op_3_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_1_itm_2 <= 1'b0;
    else
      alu_loop_op_3_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_1_itm_2 <= _0277_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      alu_loop_op_4_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_3_itm_2 <= 1'b0;
    else
      alu_loop_op_4_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_3_itm_2 <= _0290_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_8U_23U_land_1_lpi_1_dfm_st_5 <= 1'b0;
    else
      IsNaN_8U_23U_land_1_lpi_1_dfm_st_5 <= _0225_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_8U_23U_land_2_lpi_1_dfm_st_5 <= 1'b0;
    else
      IsNaN_8U_23U_land_2_lpi_1_dfm_st_5 <= _0231_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_8U_23U_land_3_lpi_1_dfm_st_5 <= 1'b0;
    else
      IsNaN_8U_23U_land_3_lpi_1_dfm_st_5 <= _0237_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_8U_23U_land_lpi_1_dfm_st_5 <= 1'b0;
    else
      IsNaN_8U_23U_land_lpi_1_dfm_st_5 <= _0243_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpAdd_8U_23U_qr_2_lpi_1_dfm_7 <= 8'b00000000;
    else
      FpAdd_8U_23U_qr_2_lpi_1_dfm_7 <= _0119_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpAdd_8U_23U_qr_3_lpi_1_dfm_7 <= 8'b00000000;
    else
      FpAdd_8U_23U_qr_3_lpi_1_dfm_7 <= _0122_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpAdd_8U_23U_qr_4_lpi_1_dfm_7 <= 8'b00000000;
    else
      FpAdd_8U_23U_qr_4_lpi_1_dfm_7 <= _0125_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpAdd_8U_23U_qr_lpi_1_dfm_7 <= 8'b00000000;
    else
      FpAdd_8U_23U_qr_lpi_1_dfm_7 <= _0128_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      main_stage_v_3 <= 1'b0;
    else
      main_stage_v_3 <= _0359_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_8U_23U_1_land_lpi_1_dfm_7 <= 1'b0;
    else
      IsNaN_8U_23U_1_land_lpi_1_dfm_7 <= _0206_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_8U_23U_1_land_3_lpi_1_dfm_7 <= 1'b0;
    else
      IsNaN_8U_23U_1_land_3_lpi_1_dfm_7 <= _0203_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_8U_23U_1_land_2_lpi_1_dfm_7 <= 1'b0;
    else
      IsNaN_8U_23U_1_land_2_lpi_1_dfm_7 <= _0200_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_8U_23U_1_land_1_lpi_1_dfm_7 <= 1'b0;
    else
      IsNaN_8U_23U_1_land_1_lpi_1_dfm_7 <= _0197_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      io_read_cfg_alu_bypass_rsc_svs_st_5 <= 1'b0;
    else
      io_read_cfg_alu_bypass_rsc_svs_st_5 <= _0354_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      alu_loop_op_unequal_tmp_6 <= 1'b0;
    else
      alu_loop_op_unequal_tmp_6 <= _0294_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      AluIn_data_sva_128 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    else
      AluIn_data_sva_128 <= _0058_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      io_read_cfg_alu_bypass_rsc_svs_6 <= 1'b0;
    else
      io_read_cfg_alu_bypass_rsc_svs_6 <= _0350_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cfg_alu_algo_1_sva_st_23 <= 2'b00;
    else
      cfg_alu_algo_1_sva_st_23 <= _0301_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      else_AluOp_data_0_lpi_1_dfm_2_30_0_1 <= 31'b0000000000000000000000000000000;
    else
      else_AluOp_data_0_lpi_1_dfm_2_30_0_1 <= _0329_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      else_AluOp_data_2_lpi_1_dfm_2_30_0_1 <= 31'b0000000000000000000000000000000;
    else
      else_AluOp_data_2_lpi_1_dfm_2_30_0_1 <= _0331_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      else_AluOp_data_1_lpi_1_dfm_2_30_0_1 <= 31'b0000000000000000000000000000000;
    else
      else_AluOp_data_1_lpi_1_dfm_2_30_0_1 <= _0330_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      else_AluOp_data_3_lpi_1_dfm_2_30_0_1 <= 31'b0000000000000000000000000000000;
    else
      else_AluOp_data_3_lpi_1_dfm_2_30_0_1 <= _0332_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpAdd_8U_23U_a_right_shift_qr_1_lpi_1_dfm_5 <= 8'b00000000;
    else
      FpAdd_8U_23U_a_right_shift_qr_1_lpi_1_dfm_5 <= _0078_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpAdd_8U_23U_b_right_shift_qr_1_lpi_1_dfm_5 <= 8'b00000000;
    else
      FpAdd_8U_23U_b_right_shift_qr_1_lpi_1_dfm_5 <= _0090_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpAdd_8U_23U_a_right_shift_qr_2_lpi_1_dfm_5 <= 8'b00000000;
    else
      FpAdd_8U_23U_a_right_shift_qr_2_lpi_1_dfm_5 <= _0080_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpAdd_8U_23U_b_right_shift_qr_2_lpi_1_dfm_5 <= 8'b00000000;
    else
      FpAdd_8U_23U_b_right_shift_qr_2_lpi_1_dfm_5 <= _0092_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpAdd_8U_23U_a_right_shift_qr_3_lpi_1_dfm_5 <= 8'b00000000;
    else
      FpAdd_8U_23U_a_right_shift_qr_3_lpi_1_dfm_5 <= _0082_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpAdd_8U_23U_b_right_shift_qr_3_lpi_1_dfm_5 <= 8'b00000000;
    else
      FpAdd_8U_23U_b_right_shift_qr_3_lpi_1_dfm_5 <= _0094_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpAdd_8U_23U_a_right_shift_qr_lpi_1_dfm_5 <= 8'b00000000;
    else
      FpAdd_8U_23U_a_right_shift_qr_lpi_1_dfm_5 <= _0084_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpAdd_8U_23U_b_right_shift_qr_lpi_1_dfm_5 <= 8'b00000000;
    else
      FpAdd_8U_23U_b_right_shift_qr_lpi_1_dfm_5 <= _0096_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      alu_loop_op_1_FpAdd_8U_23U_IsZero_8U_23U_1_or_itm_2 <= 1'b0;
    else
      alu_loop_op_1_FpAdd_8U_23U_IsZero_8U_23U_1_or_itm_2 <= _0245_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      alu_loop_op_2_FpAdd_8U_23U_IsZero_8U_23U_1_or_itm_2 <= 1'b0;
    else
      alu_loop_op_2_FpAdd_8U_23U_IsZero_8U_23U_1_or_itm_2 <= _0256_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      alu_loop_op_3_FpAdd_8U_23U_IsZero_8U_23U_1_or_itm_2 <= 1'b0;
    else
      alu_loop_op_3_FpAdd_8U_23U_IsZero_8U_23U_1_or_itm_2 <= _0269_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      alu_loop_op_4_FpAdd_8U_23U_IsZero_8U_23U_1_or_itm_2 <= 1'b0;
    else
      alu_loop_op_4_FpAdd_8U_23U_IsZero_8U_23U_1_or_itm_2 <= _0282_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      reg_alu_loop_op_4_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_3_svs_1_cse <= 1'b0;
    else
      reg_alu_loop_op_4_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_3_svs_1_cse <= _0378_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      reg_alu_loop_op_3_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_1_svs_1_cse <= 1'b0;
    else
      reg_alu_loop_op_3_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_1_svs_1_cse <= _0377_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      reg_alu_loop_op_2_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_2_svs_1_cse <= 1'b0;
    else
      reg_alu_loop_op_2_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_2_svs_1_cse <= _0376_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      reg_alu_loop_op_1_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_1_cse <= 1'b0;
    else
      reg_alu_loop_op_1_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_1_cse <= _0375_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_8U_23U_land_lpi_1_dfm_st_4 <= 1'b0;
    else
      IsNaN_8U_23U_land_lpi_1_dfm_st_4 <= _0242_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      alu_loop_op_2_FpAdd_8U_23U_IsZero_8U_23U_or_itm_4 <= 1'b0;
    else
      alu_loop_op_2_FpAdd_8U_23U_IsZero_8U_23U_or_itm_4 <= _0258_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      alu_loop_op_3_FpAdd_8U_23U_IsZero_8U_23U_or_itm_5 <= 1'b0;
    else
      alu_loop_op_3_FpAdd_8U_23U_IsZero_8U_23U_or_itm_5 <= _0272_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      alu_loop_op_4_FpAdd_8U_23U_IsZero_8U_23U_or_itm_5 <= 1'b0;
    else
      alu_loop_op_4_FpAdd_8U_23U_IsZero_8U_23U_or_itm_5 <= _0285_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_8U_23U_land_1_lpi_1_dfm_st_4 <= 1'b0;
    else
      IsNaN_8U_23U_land_1_lpi_1_dfm_st_4 <= _0224_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_8U_23U_land_2_lpi_1_dfm_st_4 <= 1'b0;
    else
      IsNaN_8U_23U_land_2_lpi_1_dfm_st_4 <= _0230_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_8U_23U_land_3_lpi_1_dfm_st_4 <= 1'b0;
    else
      IsNaN_8U_23U_land_3_lpi_1_dfm_st_4 <= _0236_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpAdd_8U_23U_is_a_greater_lor_2_lpi_1_dfm_6 <= 1'b0;
    else
      FpAdd_8U_23U_is_a_greater_lor_2_lpi_1_dfm_6 <= _0106_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpAdd_8U_23U_is_a_greater_lor_1_lpi_1_dfm_6 <= 1'b0;
    else
      FpAdd_8U_23U_is_a_greater_lor_1_lpi_1_dfm_6 <= _0105_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpAdd_8U_23U_is_a_greater_lor_3_lpi_1_dfm_6 <= 1'b0;
    else
      FpAdd_8U_23U_is_a_greater_lor_3_lpi_1_dfm_6 <= _0107_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpAdd_8U_23U_is_a_greater_lor_lpi_1_dfm_6 <= 1'b0;
    else
      FpAdd_8U_23U_is_a_greater_lor_lpi_1_dfm_6 <= _0108_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      alu_loop_op_1_FpAdd_8U_23U_IsZero_8U_23U_or_itm_3 <= 1'b0;
    else
      alu_loop_op_1_FpAdd_8U_23U_IsZero_8U_23U_or_itm_3 <= _0246_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      main_stage_v_2 <= 1'b0;
    else
      main_stage_v_2 <= _0358_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      io_read_cfg_alu_bypass_rsc_svs_st_1 <= 1'b0;
    else
      io_read_cfg_alu_bypass_rsc_svs_st_1 <= _0353_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cfg_alu_src_1_sva_st_1 <= 1'b0;
    else
      cfg_alu_src_1_sva_st_1 <= _0307_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cfg_alu_op_1_sva_1 <= 32'd0;
    else
      cfg_alu_op_1_sva_1 <= _0305_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cfg_alu_algo_1_sva_st_22 <= 2'b00;
    else
      cfg_alu_algo_1_sva_st_22 <= _0300_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      reg_cfg_alu_algo_1_sva_st_13_cse <= 2'b00;
    else
      reg_cfg_alu_algo_1_sva_st_13_cse <= _0387_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cfg_alu_algo_1_sva_st_28 <= 2'b00;
    else
      cfg_alu_algo_1_sva_st_28 <= _0304_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_8U_23U_land_lpi_1_dfm_8 <= 1'b0;
    else
      IsNaN_8U_23U_land_lpi_1_dfm_8 <= _0240_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_8U_23U_land_3_lpi_1_dfm_8 <= 1'b0;
    else
      IsNaN_8U_23U_land_3_lpi_1_dfm_8 <= _0234_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_8U_23U_land_2_lpi_1_dfm_8 <= 1'b0;
    else
      IsNaN_8U_23U_land_2_lpi_1_dfm_8 <= _0228_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_8U_23U_land_1_lpi_1_dfm_8 <= 1'b0;
    else
      IsNaN_8U_23U_land_1_lpi_1_dfm_8 <= _0222_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      AluIn_data_sva_127 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    else
      AluIn_data_sva_127 <= _0057_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      io_read_cfg_alu_bypass_rsc_svs_5 <= 1'b0;
    else
      io_read_cfg_alu_bypass_rsc_svs_5 <= _0349_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      main_stage_v_1 <= 1'b0;
    else
      main_stage_v_1 <= _0357_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_alu_op_rsci_ld_core_psct <= 1'b0;
    else
      chn_alu_op_rsci_ld_core_psct <= _0311_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      reg_chn_alu_out_rsci_ld_core_psct_cse <= 1'b0;
    else
      reg_chn_alu_out_rsci_ld_core_psct_cse <= _0389_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_alu_out_rsci_d_94_87 <= 8'b00000000;
    else
      chn_alu_out_rsci_d_94_87 <= _0325_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_alu_out_rsci_d_86_65 <= 22'b0000000000000000000000;
    else
      chn_alu_out_rsci_d_86_65 <= _0324_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_alu_out_rsci_d_64 <= 1'b0;
    else
      chn_alu_out_rsci_d_64 <= _0323_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_alu_out_rsci_d_127 <= 1'b0;
    else
      chn_alu_out_rsci_d_127 <= _0315_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_alu_out_rsci_d_126_119 <= 8'b00000000;
    else
      chn_alu_out_rsci_d_126_119 <= _0314_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_alu_out_rsci_d_118_97 <= 22'b0000000000000000000000;
    else
      chn_alu_out_rsci_d_118_97 <= _0313_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_alu_out_rsci_d_95 <= 1'b0;
    else
      chn_alu_out_rsci_d_95 <= _0326_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_alu_out_rsci_d_63 <= 1'b0;
    else
      chn_alu_out_rsci_d_63 <= _0322_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_alu_out_rsci_d_62_55 <= 8'b00000000;
    else
      chn_alu_out_rsci_d_62_55 <= _0321_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_alu_out_rsci_d_31 <= 1'b0;
    else
      chn_alu_out_rsci_d_31 <= _0318_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_alu_out_rsci_d_30_23 <= 8'b00000000;
    else
      chn_alu_out_rsci_d_30_23 <= _0317_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_alu_out_rsci_d_22_1 <= 22'b0000000000000000000000;
    else
      chn_alu_out_rsci_d_22_1 <= _0316_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_alu_out_rsci_d_54_33 <= 22'b0000000000000000000000;
    else
      chn_alu_out_rsci_d_54_33 <= _0320_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_alu_out_rsci_d_0 <= 1'b0;
    else
      chn_alu_out_rsci_d_0 <= _0312_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_alu_out_rsci_d_96 <= 1'b0;
    else
      chn_alu_out_rsci_d_96 <= _0327_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_alu_out_rsci_d_32 <= 1'b0;
    else
      chn_alu_out_rsci_d_32 <= _0319_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_alu_in_rsci_ld_core_psct <= 1'b0;
    else
      chn_alu_in_rsci_ld_core_psct <= _0309_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_alu_out_rsci_iswt0 <= 1'b0;
    else
      chn_alu_out_rsci_iswt0 <= _0328_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_alu_op_rsci_iswt0 <= 1'b0;
    else
      chn_alu_op_rsci_iswt0 <= _0310_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_alu_in_rsci_iswt0 <= 1'b0;
    else
      chn_alu_in_rsci_iswt0 <= _0308_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      reg_cfg_alu_algo_rsc_triosy_obj_ld_core_psct_cse <= 1'b0;
    else
      reg_cfg_alu_algo_rsc_triosy_obj_ld_core_psct_cse <= _0388_;
  assign FpAdd_8U_23U_else_2_mux_15_nl = FpAdd_8U_23U_if_2_and_tmp_3 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16549|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16548" *) FpAdd_8U_23U_addend_smaller_qr_lpi_1_dfm_mx0 : FpAdd_8U_23U_addend_larger_qr_lpi_1_dfm_mx0;
  assign FpAdd_8U_23U_else_2_mux_14_nl = FpAdd_8U_23U_if_2_and_tmp_3 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16549|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16548" *) FpAdd_8U_23U_addend_larger_qr_lpi_1_dfm_mx0 : _0028_;
  assign FpAdd_8U_23U_else_2_mux_13_nl = FpAdd_8U_23U_if_2_and_tmp_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16549|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16548" *) FpAdd_8U_23U_addend_smaller_qr_3_lpi_1_dfm_mx0 : FpAdd_8U_23U_addend_larger_qr_3_lpi_1_dfm_mx0;
  assign FpAdd_8U_23U_else_2_mux_12_nl = FpAdd_8U_23U_if_2_and_tmp_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16549|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16548" *) FpAdd_8U_23U_addend_larger_qr_3_lpi_1_dfm_mx0 : _0027_;
  assign FpAdd_8U_23U_else_2_mux_11_nl = FpAdd_8U_23U_if_2_and_tmp_1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16549|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16548" *) FpAdd_8U_23U_addend_smaller_qr_2_lpi_1_dfm_mx0 : FpAdd_8U_23U_addend_larger_qr_2_lpi_1_dfm_mx0;
  assign FpAdd_8U_23U_else_2_mux_10_nl = FpAdd_8U_23U_if_2_and_tmp_1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16549|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16548" *) FpAdd_8U_23U_addend_larger_qr_2_lpi_1_dfm_mx0 : _0026_;
  assign FpAdd_8U_23U_else_2_mux_9_nl = FpAdd_8U_23U_if_2_and_tmp ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16549|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16548" *) FpAdd_8U_23U_addend_smaller_qr_1_lpi_1_dfm_mx0 : FpAdd_8U_23U_addend_larger_qr_1_lpi_1_dfm_mx0;
  assign FpAdd_8U_23U_else_2_mux_8_nl = FpAdd_8U_23U_if_2_and_tmp ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16549|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16548" *) FpAdd_8U_23U_addend_larger_qr_1_lpi_1_dfm_mx0 : _0025_;
  assign FpAdd_8U_23U_b_right_shift_qif_mux_22_nl = FpAdd_8U_23U_a_right_shift_qelse_and_tmp_3 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16600|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16599" *) _0040_ : _0039_;
  assign FpAdd_8U_23U_b_right_shift_qif_mux_21_nl = FpAdd_8U_23U_a_right_shift_qelse_and_tmp_3 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16600|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16599" *) else_AluOp_data_0_lpi_1_dfm_mx0[30:23] : AluIn_data_sva_127[30:23];
  assign FpAdd_8U_23U_b_right_shift_qif_mux_20_nl = FpAdd_8U_23U_a_right_shift_qelse_and_tmp_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16600|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16599" *) _0038_ : _0037_;
  assign FpAdd_8U_23U_b_right_shift_qif_mux_19_nl = FpAdd_8U_23U_a_right_shift_qelse_and_tmp_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16600|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16599" *) else_AluOp_data_1_lpi_1_dfm_mx2_30_0[30:23] : AluIn_data_sva_127[62:55];
  assign FpAdd_8U_23U_b_right_shift_qif_mux_18_nl = FpAdd_8U_23U_a_right_shift_qelse_and_tmp_1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16600|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16599" *) _0036_ : _0035_;
  assign FpAdd_8U_23U_b_right_shift_qif_mux_17_nl = FpAdd_8U_23U_a_right_shift_qelse_and_tmp_1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16600|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16599" *) else_AluOp_data_2_lpi_1_dfm_mx0[30:23] : AluIn_data_sva_127[94:87];
  assign FpAdd_8U_23U_b_right_shift_qif_mux_16_nl = FpAdd_8U_23U_a_right_shift_qelse_and_tmp ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16600|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16599" *) _0034_ : _0033_;
  assign FpAdd_8U_23U_b_right_shift_qif_mux_15_nl = FpAdd_8U_23U_a_right_shift_qelse_and_tmp ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16600|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16599" *) else_AluOp_data_3_lpi_1_dfm_mx0[30:23] : AluIn_data_sva_127[126:119];
  assign mux_314_nl = _1527_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) mux_tmp_296 : mux_313_nl;
  assign mux_313_nl = and_489_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) mux_tmp_296 : mux_312_cse;
  assign mux_305_nl = _1527_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) nor_tmp_126 : mux_304_nl;
  assign mux_304_nl = and_489_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) nor_tmp_126 : and_451_cse;
  assign mux_303_nl = or_1087_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) mux_301_nl : nand_38_nl;
  assign mux_302_nl = io_read_cfg_alu_bypass_rsc_svs_st_1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) io_read_cfg_alu_bypass_rsc_svs_5 : mux_tmp_281;
  assign mux_301_nl = or_tmp_386 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) nand_37_nl : mux_299_nl;
  assign mux_300_nl = io_read_cfg_alu_bypass_rsc_svs_st_1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) nor_177_cse : nor_176_nl;
  assign mux_299_nl = main_stage_v_1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) mux_298_nl : mux_tmp_265;
  assign mux_298_nl = io_read_cfg_alu_bypass_rsc_svs_st_1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) mux_281_cse : mux_297_nl;
  assign mux_297_nl = and_501_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) mux_tmp_265 : mux_tmp_281;
  assign mux_290_nl = or_1087_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) mux_288_nl : nand_36_nl;
  assign mux_289_nl = io_read_cfg_alu_bypass_rsc_svs_st_1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) io_read_cfg_alu_bypass_rsc_svs_5 : mux_tmp_268;
  assign mux_288_nl = or_tmp_386 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) nand_35_nl : mux_286_nl;
  assign mux_287_nl = io_read_cfg_alu_bypass_rsc_svs_st_1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) nor_177_cse : nor_178_nl;
  assign mux_286_nl = main_stage_v_1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) mux_285_nl : mux_tmp_265;
  assign mux_285_nl = io_read_cfg_alu_bypass_rsc_svs_st_1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) mux_281_cse : mux_284_nl;
  assign mux_284_nl = and_501_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) mux_tmp_265 : mux_tmp_268;
  assign mux_277_nl = main_stage_v_1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) mux_276_nl : or_tmp_596;
  assign mux_276_nl = io_read_cfg_alu_bypass_rsc_svs_st_1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) mux_271_nl : mux_275_nl;
  assign mux_275_nl = or_619_nl ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) mux_272_nl : mux_274_nl;
  assign mux_274_nl = and_501_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) mux_273_nl : not_tmp_261;
  assign mux_273_nl = or_1087_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) or_624_nl : not_tmp_261;
  assign mux_272_nl = and_501_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) or_tmp_596 : or_tmp_597;
  assign mux_271_nl = and_486_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) or_tmp_596 : or_tmp_597;
  assign mux_175_nl = or_1087_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) mux_174_nl : nand_30_nl;
  assign mux_174_nl = main_stage_v_1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) mux_173_nl : or_tmp_386;
  assign mux_173_nl = and_486_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) and_74_nl : nor_tmp_74;
  assign alu_loop_op_else_mux_4_nl = io_read_cfg_alu_bypass_rsc_svs_st_1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) IsNaN_8U_23U_2_IsNaN_8U_23U_2_nor_itm_2 : alu_loop_op_else_equal_tmp_2;
  assign alu_loop_op_else_mux_5_nl = io_read_cfg_alu_bypass_rsc_svs_st_1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) IsNaN_8U_23U_2_IsNaN_8U_23U_2_nor_3_itm_2 : FpAlu_8U_23U_equal_tmp_1_mx0w0;
  assign mux_366_nl = or_1050_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) alu_loop_op_4_IntSaturation_33U_32U_if_acc_1_nl[2] : or_1076_nl;
  assign mux_365_nl = or_1050_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) alu_loop_op_3_IntSaturation_33U_32U_if_acc_nl[2] : or_1069_nl;
  assign mux_364_nl = or_1050_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) alu_loop_op_2_IntSaturation_33U_32U_if_acc_1_nl[2] : or_1055_cse;
  assign mux_363_nl = or_1050_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) alu_loop_op_1_IntSaturation_33U_32U_if_acc_nl[2] : or_1055_cse;
  assign mux_226_nl = or_1087_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) nor_192_nl : nor_264_cse;
  assign mux_225_nl = or_1087_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) nor_195_nl : nor_197_cse;
  assign mux_223_nl = or_1087_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) nor_201_cse : nor_203_nl;
  assign alu_loop_op_else_mux_3_nl = io_read_cfg_alu_bypass_rsc_svs_st_1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) IsNaN_8U_23U_4_nor_2_itm_2 : alu_loop_op_else_equal_tmp_2;
  assign FpAlu_8U_23U_mux_20_nl = io_read_cfg_alu_bypass_rsc_svs_st_1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) IsNaN_8U_23U_2_IsNaN_8U_23U_2_nor_1_itm_1 : FpAlu_8U_23U_equal_tmp_2_mx0w0;
  assign FpAlu_8U_23U_mux_21_nl = io_read_cfg_alu_bypass_rsc_svs_st_1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) IsNaN_8U_23U_2_IsNaN_8U_23U_2_nor_2_itm_1 : FpAlu_8U_23U_equal_tmp_1_mx0w0;
  assign alu_loop_op_else_mux_nl = io_read_cfg_alu_bypass_rsc_svs_st_1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) alu_loop_op_4_FpAdd_8U_23U_IsZero_8U_23U_or_itm_4 : alu_loop_op_else_equal_tmp_2;
  assign alu_loop_op_else_mux_2_nl = io_read_cfg_alu_bypass_rsc_svs_st_1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) IsNaN_8U_23U_4_nor_3_itm_3 : FpAlu_8U_23U_equal_tmp_2_mx0w0;
  assign alu_loop_op_else_mux_1_nl = io_read_cfg_alu_bypass_rsc_svs_st_1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) alu_loop_op_3_FpAdd_8U_23U_IsZero_8U_23U_or_itm_4 : FpAlu_8U_23U_equal_tmp_1_mx0w0;
  assign mux_219_nl = or_1087_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) and_481_cse : nor_206_nl;
  assign mux_218_nl = or_1087_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) and_481_cse : nor_207_nl;
  assign mux_212_nl = or_1087_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) nor_213_nl : nor_214_nl;
  assign mux_211_nl = or_1087_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) nor_215_nl : nor_216_nl;
  assign mux_210_nl = or_1087_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) nor_217_nl : nor_218_nl;
  assign mux_209_nl = or_1087_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) nor_219_nl : nor_220_nl;
  assign mux_208_nl = or_1087_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) mux_207_nl : nor_223_nl;
  assign mux_207_nl = alu_loop_op_unequal_tmp_6 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) nor_236_cse : nor_222_nl;
  assign mux_206_nl = or_1087_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) mux_205_nl : nor_228_nl;
  assign mux_205_nl = alu_loop_op_unequal_tmp_6 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) nor_236_cse : nor_227_nl;
  assign mux_204_nl = or_1087_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) mux_203_nl : nor_233_nl;
  assign mux_203_nl = alu_loop_op_unequal_tmp_6 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) nor_236_cse : nor_232_nl;
  assign mux_200_nl = or_1087_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) mux_199_nl : nor_238_nl;
  assign mux_199_nl = alu_loop_op_unequal_tmp_6 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) nor_236_cse : nor_237_nl;
  assign mux_196_nl = _2200_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) or_450_nl : mux_195_nl;
  assign mux_195_nl = or_1087_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) or_tmp_395 : or_tmp_261;
  assign mux_194_nl = or_444_nl ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) or_446_nl : mux_193_nl;
  assign mux_193_nl = or_1087_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) or_tmp_395 : or_tmp_293;
  assign mux_190_nl = FpAlu_8U_23U_equal_tmp_24 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) mux_189_nl : or_440_nl;
  assign mux_189_nl = FpAlu_8U_23U_equal_tmp_25 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) mux_tmp_173 : or_438_nl;
  assign mux_182_nl = alu_loop_op_unequal_tmp_6 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) mux_tmp_165 : mux_181_nl;
  assign mux_181_nl = or_420_nl ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) or_422_nl : mux_tmp_165;
  assign mux_172_nl = _1527_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) or_tmp_382 : mux_171_nl;
  assign mux_171_nl = and_489_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) or_tmp_382 : or_400_nl;
  assign mux_160_nl = alu_loop_op_4_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_3_itm ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) nor_249_nl : or_958_nl;
  assign mux_159_nl = alu_loop_op_3_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_1_itm ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) nor_250_nl : or_959_nl;
  assign mux_158_nl = alu_loop_op_2_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_2_itm ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) nor_251_nl : or_960_nl;
  assign mux_157_nl = alu_loop_op_1_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_itm ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) nor_252_nl : or_961_nl;
  assign mux_156_nl = or_1087_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) mux_155_nl : nor_256_nl;
  assign mux_155_nl = FpAlu_8U_23U_equal_tmp_21 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) nor_254_nl : nor_264_cse;
  assign mux_154_nl = or_1087_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) mux_153_nl : nor_259_nl;
  assign mux_153_nl = FpAlu_8U_23U_equal_tmp_21 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) nor_257_nl : nor_264_cse;
  assign mux_152_nl = or_1087_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) mux_151_nl : nor_262_nl;
  assign mux_151_nl = FpAlu_8U_23U_equal_tmp_21 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) nor_260_nl : nor_264_cse;
  assign mux_150_nl = or_1087_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) mux_149_nl : nor_265_nl;
  assign mux_149_nl = FpAlu_8U_23U_equal_tmp_21 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) nor_263_nl : nor_264_cse;
  assign mux_148_nl = alu_loop_op_4_FpMantRNE_49U_24U_else_and_3_svs_st ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) or_336_nl : and_493_nl;
  assign mux_147_nl = alu_loop_op_3_FpMantRNE_49U_24U_else_and_1_svs_st ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) or_335_nl : and_494_nl;
  assign mux_146_nl = alu_loop_op_2_FpMantRNE_49U_24U_else_and_2_svs_st ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) or_334_nl : and_495_nl;
  assign mux_145_nl = alu_loop_op_1_FpMantRNE_49U_24U_else_and_svs_st ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) or_333_nl : and_496_nl;
  assign mux_362_nl = or_1087_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) mux_361_nl : and_218_nl;
  assign mux_361_nl = io_read_cfg_alu_bypass_rsc_svs_8 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) or_1046_nl : mux_nl;
  assign mux_nl = main_stage_v_4 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) or_1048_nl : nor_tmp_144;
  assign mux_139_nl = or_1087_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) or_tmp_103 : or_tmp_224;
  assign mux_138_nl = or_1087_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) or_tmp_280 : or_tmp_218;
  assign mux_137_nl = or_1087_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) nor_267_nl : nor_268_nl;
  assign mux_136_nl = or_1087_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) or_tmp_293 : or_312_nl;
  assign mux_135_nl = FpAlu_8U_23U_equal_tmp_23 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) mux_134_nl : or_307_nl;
  assign mux_134_nl = or_1087_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) or_304_nl : or_tmp_218;
  assign mux_133_nl = FpAlu_8U_23U_equal_tmp_25 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) mux_132_nl : or_301_nl;
  assign mux_132_nl = or_1087_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) or_tmp_280 : or_299_nl;
  assign mux_131_nl = or_1087_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) nor_270_nl : nor_271_nl;
  assign mux_130_nl = or_1087_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) nor_272_nl : nor_273_nl;
  assign mux_128_nl = or_1087_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) nor_274_nl : nor_275_nl;
  assign mux_127_nl = or_1087_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) or_tmp_261 : or_280_nl;
  assign mux_383_nl = asn_267 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) or_1100_nl : or_1106_nl;
  assign mux_100_nl = or_1087_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) mux_99_nl : nor_300_nl;
  assign mux_99_nl = or_1050_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) nor_299_nl : nor_298_nl;
  assign mux_98_nl = or_1087_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) mux_97_nl : nor_303_nl;
  assign mux_97_nl = or_1050_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) nor_302_nl : nor_301_nl;
  assign mux_96_nl = or_1087_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) mux_95_nl : nor_306_nl;
  assign mux_95_nl = or_1050_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) nor_305_nl : nor_304_nl;
  assign mux_94_nl = or_1087_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) mux_93_nl : nor_309_nl;
  assign mux_93_nl = or_1050_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) nor_308_nl : nor_307_nl;
  assign mux_92_nl = or_1087_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) mux_88_nl : nor_313_nl;
  assign mux_91_nl = FpAdd_8U_23U_and_3_tmp_3 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) or_182_nl : or_962_nl;
  assign mux_88_nl = or_1050_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) nor_312_nl : and_497_nl;
  assign mux_87_nl = alu_loop_op_4_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_3_itm_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) nor_310_nl : nor_311_nl;
  assign mux_86_nl = or_1087_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) nor_314_nl : nor_319_nl;
  assign mux_85_nl = FpAdd_8U_23U_and_2_tmp_3 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) nor_320_nl : nor_322_nl;
  assign mux_82_nl = or_1050_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) nor_318_nl : and_498_nl;
  assign mux_81_nl = alu_loop_op_3_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_1_itm_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) nor_316_nl : nor_317_nl;
  assign mux_80_nl = or_1087_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) nor_324_nl : nor_329_nl;
  assign mux_79_nl = FpAdd_8U_23U_and_1_tmp_3 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) nor_330_nl : nor_332_nl;
  assign mux_76_nl = or_1050_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) nor_328_nl : and_499_nl;
  assign mux_75_nl = alu_loop_op_2_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_2_itm_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) nor_326_nl : nor_327_nl;
  assign mux_74_nl = or_1087_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) nor_334_nl : nor_339_nl;
  assign mux_73_nl = FpAdd_8U_23U_and_tmp_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) nor_340_nl : nor_342_nl;
  assign mux_70_nl = or_1050_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) nor_338_nl : and_500_nl;
  assign mux_69_nl = alu_loop_op_1_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_itm_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) nor_336_nl : nor_337_nl;
  assign mux_67_nl = io_read_cfg_alu_bypass_rsc_svs_st_5 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) nor_344_nl : mux_66_nl;
  assign mux_66_nl = or_1087_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) main_stage_v_2 : _0016_;
  assign mux_65_nl = or_1087_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) mux_64_nl : nor_347_nl;
  assign mux_64_nl = or_1050_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) nor_346_nl : nor_345_nl;
  assign mux_63_nl = or_1087_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) mux_62_nl : nor_350_nl;
  assign mux_62_nl = or_1050_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) nor_349_nl : nor_348_nl;
  assign mux_61_nl = or_1087_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) mux_60_nl : nor_353_nl;
  assign mux_60_nl = or_1050_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) nor_352_nl : nor_351_nl;
  assign mux_59_nl = or_1087_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) mux_58_nl : nor_356_nl;
  assign mux_58_nl = or_1050_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) nor_355_nl : nor_354_nl;
  assign mux_38_nl = main_stage_v_1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) mux_37_nl : or_tmp_23;
  assign mux_37_nl = io_read_cfg_alu_bypass_rsc_svs_st_1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) nand_18_nl : mux_36_nl;
  assign mux_36_nl = and_501_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) mux_35_nl : _0015_;
  assign mux_35_nl = or_1087_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) or_43_nl : _0015_;
  assign mux_31_nl = or_tmp_386 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) or_tmp_15 : mux_30_nl;
  assign mux_30_nl = or_1050_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) mux_29_nl : mux_27_nl;
  assign mux_29_nl = cfg_alu_algo_1_sva_st[1] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) or_tmp_15 : mux_28_nl;
  assign mux_28_nl = cfg_alu_algo_1_sva_st[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) _0014_ : or_tmp_15;
  assign mux_27_nl = cfg_alu_algo_rsci_d[1] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) or_tmp_15 : mux_26_nl;
  assign mux_26_nl = cfg_alu_algo_rsci_d[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) _0014_ : or_tmp_15;
  assign mux_23_nl = or_tmp_386 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) or_tmp_9 : mux_22_nl;
  assign mux_22_nl = or_1050_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) mux_21_nl : mux_19_nl;
  assign mux_21_nl = or_28_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) or_tmp_9 : mux_20_nl;
  assign mux_20_nl = cfg_alu_algo_1_sva_st[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) _0013_ : or_tmp_9;
  assign mux_19_nl = cfg_alu_algo_rsci_d[1] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) or_tmp_9 : mux_18_nl;
  assign mux_18_nl = cfg_alu_algo_rsci_d[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) _0013_ : or_tmp_9;
  assign FpAlu_8U_23U_and_7_nl = FpAlu_8U_23U_equal_tmp_23 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16600|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16599" *) 8'b00000000 : FpAlu_8U_23U_mux1h_149_nl;
  assign FpAlu_8U_23U_and_4_nl = FpAlu_8U_23U_equal_tmp_23 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16600|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16599" *) 8'b00000000 : FpAlu_8U_23U_mux1h_145_nl;
  assign FpAlu_8U_23U_and_8_nl = FpAlu_8U_23U_equal_tmp_23 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16464|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16463" *) 22'b0000000000000000000000 : FpAlu_8U_23U_FpAlu_8U_23U_mux_1_nl;
  assign FpAlu_8U_23U_FpAlu_8U_23U_mux_1_nl = FpAlu_8U_23U_equal_tmp_29 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16464|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16463" *) FpCmp_8U_23U_false_o_2_lpi_1_dfm_8_30_0_1[22:1] : FpCmp_8U_23U_true_o_2_lpi_1_dfm_7_30_0_1[22:1];
  assign FpAlu_8U_23U_and_5_nl = FpAlu_8U_23U_equal_tmp_23 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16464|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16463" *) 22'b0000000000000000000000 : FpAlu_8U_23U_FpAlu_8U_23U_mux_nl;
  assign FpAlu_8U_23U_FpAlu_8U_23U_mux_nl = FpAlu_8U_23U_equal_tmp_29 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16464|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16463" *) FpCmp_8U_23U_false_o_1_lpi_1_dfm_7_30_0_1[22:1] : FpCmp_8U_23U_true_o_1_lpi_1_dfm_7_30_0_1[22:1];
  assign alu_loop_op_mux_212_nl = alu_loop_op_unequal_tmp_8 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) AluOut_data_2_0_lpi_1_dfm_3 : FpAlu_8U_23U_o_0_lpi_1_dfm_2;
  assign alu_loop_op_mux_210_nl = alu_loop_op_unequal_tmp_8 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) AluOut_data_0_0_sva_11 : FpAlu_8U_23U_mux1h_151_nl;
  assign alu_loop_op_mux_209_nl = alu_loop_op_unequal_tmp_8 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) AluOut_data_2_0_sva_11 : FpAlu_8U_23U_mux1h_147_nl;
  assign mux_tmp_350 = FpAdd_8U_23U_int_mant_p1_lpi_1_dfm_5[49] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) alu_loop_op_4_FpAdd_8U_23U_if_3_if_acc_6_nl[7] : FpNormalize_8U_49U_oelse_not_15;
  assign mux_tmp_349 = FpAdd_8U_23U_int_mant_p1_3_lpi_1_dfm_5[49] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) alu_loop_op_3_FpAdd_8U_23U_if_3_if_acc_2_nl[7] : FpNormalize_8U_49U_oelse_not_13;
  assign mux_tmp_348 = FpAdd_8U_23U_int_mant_p1_2_lpi_1_dfm_5[49] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) alu_loop_op_2_FpAdd_8U_23U_if_3_if_acc_4_nl[7] : FpNormalize_8U_49U_oelse_not_11;
  assign mux_tmp = FpAdd_8U_23U_int_mant_p1_1_lpi_1_dfm_5[49] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) alu_loop_op_1_FpAdd_8U_23U_if_3_if_acc_1_nl[7] : FpNormalize_8U_49U_oelse_not_9;
  assign mux_337_itm = alu_loop_op_unequal_tmp_6 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) or_dcpl_46 : and_dcpl_99;
  assign mux_tmp_311 = or_1087_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) io_read_cfg_alu_bypass_rsc_svs_7 : io_read_cfg_alu_bypass_rsc_svs_8;
  assign mux_tmp_296 = _1147_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) or_391_cse : mux_310_nl;
  assign mux_310_nl = cfg_alu_algo_1_sva_st[1] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) cfg_alu_algo_1_sva_st[0] : _0012_;
  assign mux_tmp_281 = _1778_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) or_632_cse : mux_282_cse;
  assign mux_tmp_268 = _1777_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) or_632_cse : mux_282_cse;
  assign mux_282_cse = cfg_alu_algo_1_sva_st_22[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) cfg_alu_algo_1_sva_st_22[1] : _0011_;
  assign mux_tmp_265 = or_1050_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) mux_279_nl : mux_312_cse;
  assign mux_279_nl = cfg_alu_algo_1_sva_st[1] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) cfg_alu_algo_1_sva_st[0] : or_629_nl;
  assign mux_tmp_246 = main_stage_v_1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) mux_260_nl : or_1087_cse;
  assign mux_260_nl = io_read_cfg_alu_bypass_rsc_svs_st_1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) mux_255_nl : mux_259_nl;
  assign mux_259_nl = and_501_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) mux_258_nl : _0010_;
  assign mux_258_nl = cfg_alu_algo_1_sva_st_22[1] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) or_tmp_585 : mux_257_nl;
  assign mux_257_nl = or_612_nl ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) or_1087_cse : mux_256_nl;
  assign mux_256_nl = cfg_alu_algo_1_sva_2[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) or_tmp_583 : or_tmp_585;
  assign mux_255_nl = and_486_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) or_610_nl : _0009_;
  assign mux_254_nl = io_read_cfg_alu_bypass_rsc_svs_st_1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) mux_248_nl : mux_253_nl;
  assign mux_253_nl = and_501_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) mux_250_nl : mux_tmp_237;
  assign mux_250_nl = cfg_alu_algo_1_sva_st_22[1] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) or_tmp_583 : or_607_nl;
  assign mux_249_nl = cfg_alu_algo_1_sva_2[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) or_tmp_585 : or_tmp_583;
  assign mux_248_nl = and_486_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) or_601_nl : io_read_cfg_alu_bypass_rsc_svs_5;
  assign mux_tmp_237 = cfg_alu_algo_1_sva_st_22[1] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) cfg_alu_algo_1_sva_st_22[0] : or_609_nl;
  assign mux_251_nl = cfg_alu_algo_1_sva_2[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) _0008_ : cfg_alu_algo_1_sva_st_22[0];
  assign mux_tmp_227 = or_1087_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) and_dcpl_4 : nor_236_cse;
  assign not_tmp_232 = or_1087_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) mux_233_nl : nor_187_nl;
  assign mux_233_nl = io_read_cfg_alu_bypass_rsc_svs_st_1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) and_484_cse : and_474_nl;
  assign mux_tmp_173 = or_tmp_409 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) or_432_nl : mux_187_nl;
  assign mux_187_nl = or_1087_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) or_tmp_395 : or_tmp_280;
  assign mux_tmp_171 = alu_loop_op_unequal_tmp_6 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) or_428_nl : mux_185_nl;
  assign mux_185_nl = or_1087_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) or_tmp_395 : or_tmp_251;
  assign mux_tmp_165 = or_1087_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) or_tmp_395 : mux_tmp_164;
  assign mux_tmp_164 = FpAlu_8U_23U_equal_tmp_22 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) mux_178_nl : or_tmp_312;
  assign mux_178_nl = alu_loop_op_unequal_tmp_7 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) or_417_nl : or_419_nl;
  assign mux_163_nl = and_486_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) nor_379_nl : mux_tmp_146;
  assign mux_162_nl = and_486_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) or_383_nl : mux_tmp_146;
  assign mux_tmp_146 = io_read_cfg_alu_bypass_rsc_svs_5 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) or_386_nl : nor_248_nl;
  assign mux_143_itm = FpAlu_8U_23U_equal_tmp_23 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) mux_141_nl : mux_142_nl;
  assign mux_142_nl = or_1087_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) or_tmp_305 : or_tmp_309;
  assign mux_141_nl = or_1087_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) or_tmp_305 : or_323_nl;
  assign mux_109_itm = FpAlu_8U_23U_equal_tmp_23 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) or_230_nl : mux_108_nl;
  assign mux_108_nl = or_1087_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) or_233_nl : or_tmp_218;
  assign mux_tmp_53 = or_1087_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) main_stage_v_2 : main_stage_v_3;
  assign not_tmp_57 = or_87_nl ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) nor_357_nl : mux_56_nl;
  assign mux_56_nl = or_1087_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) main_stage_v_2 : _0007_;
  assign not_tmp_29 = or_1087_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) nor_371_nl : nor_372_nl;
  assign mux_34_itm = cfg_alu_bypass_rsci_d ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) or_tmp_20 : mux_33_nl;
  assign mux_33_nl = chn_alu_in_rsci_bawt ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) _0006_ : or_tmp_20;
  assign mux_32_nl = main_stage_v_1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) nand_17_nl : or_1087_cse;
  assign mux_tmp_10 = main_stage_v_1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) mux_24_nl : or_1087_cse;
  assign mux_24_nl = io_read_cfg_alu_bypass_rsc_svs_st_1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) and_37_cse : or_965_nl;
  assign mux_tmp_2 = main_stage_v_1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) mux_16_nl : or_1087_cse;
  assign mux_16_nl = io_read_cfg_alu_bypass_rsc_svs_st_1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) and_37_cse : or_967_nl;
  assign else_mux_tmp_31_23 = alu_loop_op_2_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_1_svs_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16617|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16616" *) chn_alu_op_rsci_d_mxwt[31:23] : cfg_alu_op_1_sva_1[31:23];
  assign else_mux_1_tmp_31_23 = alu_loop_op_2_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_1_svs_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16617|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16616" *) chn_alu_op_rsci_d_mxwt[63:55] : cfg_alu_op_1_sva_1[31:23];
  assign else_mux_2_tmp_31_23 = alu_loop_op_2_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_1_svs_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16617|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16616" *) chn_alu_op_rsci_d_mxwt[95:87] : cfg_alu_op_1_sva_1[31:23];
  assign else_mux_3_tmp_31_23 = alu_loop_op_2_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_1_svs_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16617|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16616" *) chn_alu_op_rsci_d_mxwt[127:119] : cfg_alu_op_1_sva_1[31:23];
  assign else_else_mux_13_nl = alu_loop_op_2_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_1_svs_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16481|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16480" *) chn_alu_op_rsci_d_mxwt[54:32] : cfg_alu_op_1_sva_1[22:0];
  assign FpCmp_8U_23U_false_o_2_lpi_1_dfm_2 = FpAlu_8U_23U_and_61_nl ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16532|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16531" *) else_AluOp_data_1_lpi_1_dfm_mx0 : AluIn_data_sva_127[63:32];
  assign FpCmp_8U_23U_false_mux_4_nl = AluIn_data_sva_127[63] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) FpCmp_8U_23U_false_else_1_FpCmp_8U_23U_false_else_1_and_1_nl : FpCmp_8U_23U_false_if_1_FpCmp_8U_23U_false_if_1_or_1_nl;
  assign FpCmp_8U_23U_false_o_lpi_1_dfm_1_mx0 = or_884_nl ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16532|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16531" *) AluIn_data_sva_127[127:96] : else_AluOp_data_3_lpi_1_dfm_mx0;
  assign mux_345_nl = or_871_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) and_340_nl : nor_156_nl;
  assign FpCmp_8U_23U_false_o_3_lpi_1_dfm_1_mx0 = or_880_nl ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16532|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16531" *) AluIn_data_sva_127[95:64] : else_AluOp_data_2_lpi_1_dfm_mx0;
  assign mux_344_nl = or_867_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) and_338_nl : nor_159_nl;
  assign FpCmp_8U_23U_false_o_1_lpi_1_dfm_1_mx0 = or_876_nl ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16532|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16531" *) AluIn_data_sva_127[31:0] : else_AluOp_data_0_lpi_1_dfm_mx0;
  assign mux_343_nl = or_861_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) and_336_nl : nor_162_nl;
  assign FpCmp_8U_23U_true_o_lpi_1_dfm_1_mx0 = _1715_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16532|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16531" *) AluIn_data_sva_127[127:96] : else_AluOp_data_3_lpi_1_dfm_mx0;
  assign mux_342_nl = or_871_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) nor_163_nl : and_443_nl;
  assign FpCmp_8U_23U_true_o_3_lpi_1_dfm_1_mx0 = _1712_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16532|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16531" *) AluIn_data_sva_127[95:64] : else_AluOp_data_2_lpi_1_dfm_mx0;
  assign mux_341_nl = or_867_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) nor_165_nl : and_444_nl;
  assign FpCmp_8U_23U_true_o_2_lpi_1_dfm_1_mx0 = _1709_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16532|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16531" *) AluIn_data_sva_127[63:32] : else_AluOp_data_1_lpi_1_dfm_mx0;
  assign mux_340_nl = or_864_nl ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) AluIn_data_sva_127[63] : _0005_;
  assign FpCmp_8U_23U_true_o_1_lpi_1_dfm_1_mx0 = _1706_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16532|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16531" *) AluIn_data_sva_127[31:0] : else_AluOp_data_0_lpi_1_dfm_mx0;
  assign mux_339_nl = or_861_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) nor_168_nl : and_446_nl;
  assign alu_loop_op_else_if_qr_31_0_lpi_1_dfm_mx0 = acc_9_nl[33] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16532|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16531" *) AluIn_data_sva_127[127:96] : else_AluOp_data_3_lpi_1_dfm_mx0;
  assign alu_loop_op_else_if_mux_11_nl = alu_loop_op_else_else_if_and_1_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16532|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16531" *) _0024_ : _0023_;
  assign alu_loop_op_else_if_mux_10_nl = alu_loop_op_else_else_if_and_1_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16532|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16531" *) AluIn_data_sva_127[127:96] : else_AluOp_data_3_lpi_1_dfm_mx0;
  assign alu_loop_op_else_if_qr_31_0_3_lpi_1_dfm_mx0 = acc_11_nl[33] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16532|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16531" *) AluIn_data_sva_127[95:64] : else_AluOp_data_2_lpi_1_dfm_mx0;
  assign alu_loop_op_else_if_mux_15_nl = alu_loop_op_else_else_if_and_1_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16532|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16531" *) _0022_ : _0021_;
  assign alu_loop_op_else_if_mux_14_nl = alu_loop_op_else_else_if_and_1_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16532|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16531" *) AluIn_data_sva_127[95:64] : else_AluOp_data_2_lpi_1_dfm_mx0;
  assign alu_loop_op_else_if_qr_31_0_2_lpi_1_dfm_mx0 = acc_10_nl[33] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16532|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16531" *) AluIn_data_sva_127[63:32] : else_AluOp_data_1_lpi_1_dfm_mx0;
  assign alu_loop_op_else_if_mux_13_nl = alu_loop_op_else_else_if_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16532|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16531" *) _0020_ : _0019_;
  assign alu_loop_op_else_if_mux_12_nl = alu_loop_op_else_else_if_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16532|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16531" *) AluIn_data_sva_127[63:32] : else_AluOp_data_1_lpi_1_dfm_mx0;
  assign alu_loop_op_else_if_qr_31_0_1_lpi_1_dfm_mx0 = acc_8_nl[33] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16532|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16531" *) AluIn_data_sva_127[31:0] : else_AluOp_data_0_lpi_1_dfm_mx0;
  assign alu_loop_op_else_if_mux_9_nl = alu_loop_op_else_else_if_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16532|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16531" *) _0018_ : _0017_;
  assign alu_loop_op_else_if_mux_8_nl = alu_loop_op_else_else_if_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16532|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16531" *) AluIn_data_sva_127[31:0] : else_AluOp_data_0_lpi_1_dfm_mx0;
  assign FpAlu_8U_23U_o_30_23_lpi_1_dfm_2 = FpAlu_8U_23U_equal_tmp_23 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16600|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16599" *) 8'b00000000 : FpAlu_8U_23U_mux1h_34_nl;
  assign FpAlu_8U_23U_o_22_1_lpi_1_dfm_2 = FpAlu_8U_23U_equal_tmp_23 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16464|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16463" *) 22'b0000000000000000000000 : FpAlu_8U_23U_mux1h_35_nl;
  assign FpAdd_8U_23U_int_mant_2_lpi_1_dfm_2_mx0 = FpAdd_8U_23U_int_mant_p1_1_lpi_1_dfm_5[49] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16549|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16548" *) { 1'b1, FpAdd_8U_23U_int_mant_p1_1_lpi_1_dfm_5[48:1] } : FpNormalize_8U_49U_FpNormalize_8U_49U_and_1_nl;
  assign FpNormalize_8U_49U_FpNormalize_8U_49U_and_1_nl = FpNormalize_8U_49U_oelse_not_9 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16549|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16548" *) alu_loop_op_1_FpNormalize_8U_49U_else_lshift_itm : 49'b0000000000000000000000000000000000000000000000000;
  assign FpAdd_8U_23U_int_mant_3_lpi_1_dfm_2_mx0 = FpAdd_8U_23U_int_mant_p1_2_lpi_1_dfm_5[49] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16549|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16548" *) { 1'b1, FpAdd_8U_23U_int_mant_p1_2_lpi_1_dfm_5[48:1] } : FpNormalize_8U_49U_FpNormalize_8U_49U_and_3_nl;
  assign FpNormalize_8U_49U_FpNormalize_8U_49U_and_3_nl = FpNormalize_8U_49U_oelse_not_11 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16549|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16548" *) alu_loop_op_2_FpNormalize_8U_49U_else_lshift_2_itm : 49'b0000000000000000000000000000000000000000000000000;
  assign FpAdd_8U_23U_int_mant_4_lpi_1_dfm_2_mx0 = FpAdd_8U_23U_int_mant_p1_3_lpi_1_dfm_5[49] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16549|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16548" *) { 1'b1, FpAdd_8U_23U_int_mant_p1_3_lpi_1_dfm_5[48:1] } : FpNormalize_8U_49U_FpNormalize_8U_49U_and_5_nl;
  assign FpNormalize_8U_49U_FpNormalize_8U_49U_and_5_nl = FpNormalize_8U_49U_oelse_not_13 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16549|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16548" *) alu_loop_op_3_FpNormalize_8U_49U_else_lshift_1_itm : 49'b0000000000000000000000000000000000000000000000000;
  assign FpAdd_8U_23U_int_mant_1_lpi_1_dfm_2_mx0 = FpAdd_8U_23U_int_mant_p1_lpi_1_dfm_5[49] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16549|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16548" *) { 1'b1, FpAdd_8U_23U_int_mant_p1_lpi_1_dfm_5[48:1] } : FpNormalize_8U_49U_FpNormalize_8U_49U_and_7_nl;
  assign FpNormalize_8U_49U_FpNormalize_8U_49U_and_7_nl = FpNormalize_8U_49U_oelse_not_15 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16549|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16548" *) alu_loop_op_4_FpNormalize_8U_49U_else_lshift_3_itm : 49'b0000000000000000000000000000000000000000000000000;
  assign FpAdd_8U_23U_addend_smaller_qr_lpi_1_dfm_mx0 = FpAdd_8U_23U_is_a_greater_lor_lpi_1_dfm_6 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16549|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16548" *) FpAdd_8U_23U_addend_larger_asn_1_mx0w1 : FpAdd_8U_23U_a_int_mant_p1_sva;
  assign FpAdd_8U_23U_addend_larger_qr_lpi_1_dfm_mx0 = FpAdd_8U_23U_is_a_greater_lor_lpi_1_dfm_6 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16549|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16548" *) FpAdd_8U_23U_a_int_mant_p1_sva : FpAdd_8U_23U_addend_larger_asn_1_mx0w1;
  assign FpAdd_8U_23U_addend_smaller_qr_3_lpi_1_dfm_mx0 = FpAdd_8U_23U_is_a_greater_lor_3_lpi_1_dfm_6 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16549|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16548" *) FpAdd_8U_23U_addend_larger_asn_7_mx0w1 : FpAdd_8U_23U_a_int_mant_p1_3_sva;
  assign FpAdd_8U_23U_addend_larger_qr_3_lpi_1_dfm_mx0 = FpAdd_8U_23U_is_a_greater_lor_3_lpi_1_dfm_6 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16549|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16548" *) FpAdd_8U_23U_a_int_mant_p1_3_sva : FpAdd_8U_23U_addend_larger_asn_7_mx0w1;
  assign FpAdd_8U_23U_addend_smaller_qr_2_lpi_1_dfm_mx0 = FpAdd_8U_23U_is_a_greater_lor_2_lpi_1_dfm_6 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16549|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16548" *) FpAdd_8U_23U_addend_larger_asn_13_mx0w1 : FpAdd_8U_23U_a_int_mant_p1_2_sva;
  assign FpAdd_8U_23U_addend_larger_qr_2_lpi_1_dfm_mx0 = FpAdd_8U_23U_is_a_greater_lor_2_lpi_1_dfm_6 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16549|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16548" *) FpAdd_8U_23U_a_int_mant_p1_2_sva : FpAdd_8U_23U_addend_larger_asn_13_mx0w1;
  assign FpAdd_8U_23U_addend_smaller_qr_1_lpi_1_dfm_mx0 = FpAdd_8U_23U_is_a_greater_lor_1_lpi_1_dfm_6 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16549|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16548" *) FpAdd_8U_23U_addend_larger_asn_19_mx0w1 : FpAdd_8U_23U_a_int_mant_p1_1_sva;
  assign FpAdd_8U_23U_addend_larger_qr_1_lpi_1_dfm_mx0 = FpAdd_8U_23U_is_a_greater_lor_1_lpi_1_dfm_6 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16549|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16548" *) FpAdd_8U_23U_a_int_mant_p1_1_sva : FpAdd_8U_23U_addend_larger_asn_19_mx0w1;
  assign else_AluOp_data_2_lpi_1_dfm_mx3_30_0 = alu_loop_op_2_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_1_svs_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16515|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16514" *) chn_alu_op_rsci_d_mxwt[94:64] : cfg_alu_op_1_sva_1[30:0];
  assign else_AluOp_data_2_lpi_1_dfm_mx1_tmp_30_23 = alu_loop_op_2_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_1_svs_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16600|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16599" *) chn_alu_op_rsci_d_mxwt[94:87] : cfg_alu_op_1_sva_1[30:23];
  assign else_AluOp_data_2_lpi_1_dfm_mx0 = alu_loop_op_2_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_1_svs_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16532|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16531" *) chn_alu_op_rsci_d_mxwt[95:64] : cfg_alu_op_1_sva_1;
  assign else_AluOp_data_1_lpi_1_dfm_mx2_30_0 = alu_loop_op_2_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_1_svs_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16515|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16514" *) chn_alu_op_rsci_d_mxwt[62:32] : cfg_alu_op_1_sva_1[30:0];
  assign else_AluOp_data_1_lpi_1_dfm_mx1_tmp_30_23 = alu_loop_op_2_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_1_svs_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16600|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16599" *) chn_alu_op_rsci_d_mxwt[62:55] : cfg_alu_op_1_sva_1[30:23];
  assign else_AluOp_data_1_lpi_1_dfm_mx0 = alu_loop_op_2_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_1_svs_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16532|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16531" *) chn_alu_op_rsci_d_mxwt[63:32] : cfg_alu_op_1_sva_1;
  assign else_AluOp_data_0_lpi_1_dfm_mx3_30_0 = alu_loop_op_2_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_1_svs_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16515|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16514" *) chn_alu_op_rsci_d_mxwt[30:0] : cfg_alu_op_1_sva_1[30:0];
  assign else_AluOp_data_0_lpi_1_dfm_mx1_tmp_30_23 = alu_loop_op_2_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_1_svs_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16600|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16599" *) chn_alu_op_rsci_d_mxwt[30:23] : cfg_alu_op_1_sva_1[30:23];
  assign else_AluOp_data_0_lpi_1_dfm_mx0 = alu_loop_op_2_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_1_svs_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16532|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16531" *) chn_alu_op_rsci_d_mxwt[31:0] : cfg_alu_op_1_sva_1;
  assign FpCmp_8U_23U_false_is_abs_a_greater_2_lpi_1_dfm_1_mx0 = or_dcpl_154 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) FpCmp_8U_23U_false_is_abs_a_greater_2_lpi_1_dfm_2 : FpCmp_8U_23U_false_is_abs_a_greater_2_lpi_1_dfm_1_mx0w0;
  assign else_AluOp_data_3_lpi_1_dfm_mx1_tmp_30_23 = alu_loop_op_2_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_1_svs_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16600|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16599" *) chn_alu_op_rsci_d_mxwt[126:119] : cfg_alu_op_1_sva_1[30:23];
  assign else_AluOp_data_3_lpi_1_dfm_mx0 = alu_loop_op_2_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_1_svs_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16532|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16531" *) chn_alu_op_rsci_d_mxwt[127:96] : cfg_alu_op_1_sva_1;
  assign alu_loop_op_else_o_32_1_lpi_1_dfm_mx0w0 = FpAlu_8U_23U_equal_tmp_1_mx0w0 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16532|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16531" *) 32'd0 : alu_loop_op_else_alu_loop_op_else_mux_nl;
  assign alu_loop_op_else_alu_loop_op_else_mux_nl = alu_loop_op_else_equal_tmp_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16532|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16531" *) alu_loop_op_else_else_else_else_ac_int_cctor_sva[32:1] : { alu_loop_op_else_if_qr_31_0_lpi_1_dfm_mx0[31], alu_loop_op_else_if_qr_31_0_lpi_1_dfm_mx0[31:1] };
  assign alu_loop_op_else_o_32_1_3_lpi_1_dfm_mx0w0 = FpAlu_8U_23U_equal_tmp_1_mx0w0 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16532|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16531" *) 32'd0 : alu_loop_op_else_alu_loop_op_else_mux_1_nl;
  assign alu_loop_op_else_alu_loop_op_else_mux_1_nl = alu_loop_op_else_equal_tmp_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16532|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16531" *) alu_loop_op_else_else_else_else_ac_int_cctor_3_sva[32:1] : { alu_loop_op_else_if_qr_31_0_3_lpi_1_dfm_mx0[31], alu_loop_op_else_if_qr_31_0_3_lpi_1_dfm_mx0[31:1] };
  assign alu_loop_op_else_o_32_1_2_lpi_1_dfm_mx0w0 = FpAlu_8U_23U_equal_tmp_1_mx0w0 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16532|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16531" *) 32'd0 : alu_loop_op_else_alu_loop_op_else_mux_2_nl;
  assign alu_loop_op_else_alu_loop_op_else_mux_2_nl = alu_loop_op_else_equal_tmp_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16532|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16531" *) alu_loop_op_else_else_else_else_ac_int_cctor_2_sva[32:1] : { alu_loop_op_else_if_qr_31_0_2_lpi_1_dfm_mx0[31], alu_loop_op_else_if_qr_31_0_2_lpi_1_dfm_mx0[31:1] };
  assign alu_loop_op_else_o_32_1_1_lpi_1_dfm_mx0w0 = FpAlu_8U_23U_equal_tmp_1_mx0w0 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16532|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16531" *) 32'd0 : alu_loop_op_else_alu_loop_op_else_mux_3_nl;
  assign alu_loop_op_else_alu_loop_op_else_mux_3_nl = alu_loop_op_else_equal_tmp_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16532|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16531" *) alu_loop_op_else_else_else_else_ac_int_cctor_1_sva[32:1] : { alu_loop_op_else_if_qr_31_0_1_lpi_1_dfm_mx0[31], alu_loop_op_else_if_qr_31_0_1_lpi_1_dfm_mx0[31:1] };
  assign FpNormalize_8U_49U_else_mux_7_nl = FpAdd_8U_23U_if_3_if_and_tmp_3 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16583|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16582" *) 6'b000001 : _0032_;
  assign FpNormalize_8U_49U_else_mux_6_nl = FpAdd_8U_23U_if_3_if_and_tmp_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16583|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16582" *) 6'b000001 : _0031_;
  assign FpNormalize_8U_49U_else_mux_5_nl = FpAdd_8U_23U_if_3_if_and_tmp_1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16583|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16582" *) 6'b000001 : _0030_;
  assign FpNormalize_8U_49U_else_mux_4_nl = FpAdd_8U_23U_if_3_if_and_tmp ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16583|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16582" *) 6'b000001 : _0029_;
  assign FpAdd_8U_23U_a_right_shift_qr_1_lpi_1_dfm_mx0w0 = FpAdd_8U_23U_is_a_greater_lor_1_lpi_1_dfm_1_mx0w0 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16600|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16599" *) 8'b00000000 : acc_7_nl[8:1];
  assign FpAdd_8U_23U_b_right_shift_qr_1_lpi_1_dfm_mx0w0 = FpAdd_8U_23U_is_a_greater_lor_1_lpi_1_dfm_1_mx0w0 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16600|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16599" *) acc_7_nl[8:1] : 8'b00000000;
  assign FpAdd_8U_23U_a_right_shift_qr_2_lpi_1_dfm_mx0w0 = FpAdd_8U_23U_is_a_greater_lor_2_lpi_1_dfm_1_mx0w0 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16600|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16599" *) 8'b00000000 : acc_6_nl[8:1];
  assign FpAdd_8U_23U_b_right_shift_qr_2_lpi_1_dfm_mx0w0 = FpAdd_8U_23U_is_a_greater_lor_2_lpi_1_dfm_1_mx0w0 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16600|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16599" *) acc_6_nl[8:1] : 8'b00000000;
  assign FpAdd_8U_23U_a_right_shift_qr_3_lpi_1_dfm_mx0w0 = FpAdd_8U_23U_is_a_greater_lor_3_lpi_1_dfm_1_mx0w0 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16600|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16599" *) 8'b00000000 : acc_5_nl[8:1];
  assign FpAdd_8U_23U_b_right_shift_qr_3_lpi_1_dfm_mx0w0 = FpAdd_8U_23U_is_a_greater_lor_3_lpi_1_dfm_1_mx0w0 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16600|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16599" *) acc_5_nl[8:1] : 8'b00000000;
  assign FpAdd_8U_23U_a_right_shift_qr_lpi_1_dfm_mx0w0 = FpAdd_8U_23U_is_a_greater_lor_lpi_1_dfm_1_mx0w0 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16600|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16599" *) 8'b00000000 : acc_4_nl[8:1];
  assign FpAdd_8U_23U_b_right_shift_qr_lpi_1_dfm_mx0w0 = FpAdd_8U_23U_is_a_greater_lor_lpi_1_dfm_1_mx0w0 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16600|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16599" *) acc_4_nl[8:1] : 8'b00000000;
  assign FpAlu_8U_23U_and_10_nl = FpAlu_8U_23U_equal_tmp_23 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16600|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16599" *) 8'b00000000 : FpAlu_8U_23U_mux1h_153_nl;
  assign FpAlu_8U_23U_and_11_nl = FpAlu_8U_23U_equal_tmp_23 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16464|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16463" *) 22'b0000000000000000000000 : FpAlu_8U_23U_mux1h_154_nl;
  assign alu_loop_op_mux_204_mx1w1 = alu_loop_op_unequal_tmp_8 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) AluOut_data_1_0_sva_12 : FpAlu_8U_23U_mux1h_155_nl;
  assign mux_312_cse = cfg_alu_algo_rsci_d[1] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) cfg_alu_algo_rsci_d[0] : _0004_;
  assign mux_307_nl = _1527_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) and_tmp_35 : mux_306_nl;
  assign mux_306_nl = and_489_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) and_tmp_35 : and_451_cse;
  assign mux_281_cse = and_486_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) mux_tmp_265 : io_read_cfg_alu_bypass_rsc_svs_5;
  assign mux_270_nl = or_tmp_386 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) nand_tmp_20 : mux_269_nl;
  assign mux_269_nl = or_1050_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) mux_268_nl : mux_262_nl;
  assign mux_268_nl = cfg_alu_algo_1_sva_st[1] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) mux_263_nl : mux_267_nl;
  assign mux_267_nl = cfg_alu_algo_rsci_d[1] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) nand_tmp_20 : _0003_;
  assign mux_266_nl = cfg_alu_algo_1_sva_st[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) mux_264_nl : mux_265_nl;
  assign mux_265_nl = cfg_alu_algo_rsci_d[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) _0002_ : mux_tmp_246;
  assign mux_264_nl = cfg_alu_algo_rsci_d[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) mux_tmp_246 : _0002_;
  assign mux_263_nl = cfg_alu_algo_1_sva_st[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) nand_tmp_20 : _0001_;
  assign mux_262_nl = and_451_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) nand_tmp_20 : _0001_;
  assign mux_247_nl = main_stage_v_1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) mux_246_nl : or_tmp_577;
  assign mux_246_nl = io_read_cfg_alu_bypass_rsc_svs_st_1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) mux_243_nl : mux_245_nl;
  assign mux_245_nl = io_read_cfg_alu_bypass_rsc_svs_5 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) or_tmp_577 : mux_244_nl;
  assign mux_244_nl = or_963_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) _0000_ : or_tmp_577;
  assign mux_243_nl = io_read_cfg_alu_bypass_rsc_svs_5 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) or_tmp_577 : _0000_;
  assign alu_loop_op_else_o_mux1h_7_itm = mux_337_itm ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16532|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16531" *) alu_loop_op_else_o_32_1_lpi_1_dfm_mx0w0 : { 1'b0, FpCmp_8U_23U_false_o_lpi_1_dfm_1_mx0[30:0] };
  assign alu_loop_op_else_o_mux1h_5_itm = mux_337_itm ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16532|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16531" *) alu_loop_op_else_o_32_1_3_lpi_1_dfm_mx0w0 : { 1'b0, FpCmp_8U_23U_false_o_3_lpi_1_dfm_1_mx0[30:0] };
  assign alu_loop_op_else_o_mux1h_3_itm = mux_337_itm ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16532|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16531" *) alu_loop_op_else_o_32_1_2_lpi_1_dfm_mx0w0 : { 1'b0, FpCmp_8U_23U_false_o_2_lpi_1_dfm_2[30:0] };
  assign alu_loop_op_else_o_mux1h_1_itm = mux_337_itm ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16532|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16531" *) alu_loop_op_else_o_32_1_1_lpi_1_dfm_mx0w0 : { 1'b0, FpCmp_8U_23U_false_o_1_lpi_1_dfm_1_mx0[30:0] };
  assign mux_224_nl = or_1087_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) nor_201_cse : nor_200_nl;
  assign mux_222_nl = or_1087_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) and_478_nl : nor_205_nl;
  assign mux_221_nl = _1561_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) nor_204_nl : or_963_cse;
  assign mux_217_nl = or_1087_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) nor_208_nl : nor_210_nl;
  assign mux_216_nl = _1527_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) or_391_cse : mux_215_nl;
  assign mux_215_nl = and_489_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) or_391_cse : or_381_cse;
  assign mux_214_nl = or_1087_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) mux_213_nl : nor_197_cse;
  assign mux_213_nl = io_read_cfg_alu_bypass_rsc_svs_st_1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) and_484_cse : and_485_nl;
  assign mux_202_nl = alu_loop_op_unequal_tmp_6 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) mux_201_nl : or_463_nl;
  assign mux_201_nl = or_1087_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) or_tmp_395 : or_tmp_312;
  assign mux_198_nl = _1542_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) or_453_nl : mux_197_nl;
  assign mux_197_nl = or_1087_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) or_tmp_395 : or_tmp_269;
  assign mux_192_nl = FpAlu_8U_23U_equal_tmp_24 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) mux_191_nl : or_443_nl;
  assign mux_191_nl = FpAlu_8U_23U_equal_tmp_25 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) mux_tmp_171 : or_441_nl;
  assign mux_184_nl = or_tmp_402 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) mux_183_nl : or_426_nl;
  assign mux_183_nl = or_1087_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) or_tmp_395 : or_tmp_305;
  assign mux_177_nl = or_1087_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) mux_176_nl : nor_243_nl;
  assign mux_176_nl = FpAlu_8U_23U_equal_tmp_21 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) nor_241_nl : nor_264_cse;
  assign mux_168_nl = or_1087_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) mux_167_nl : nand_29_nl;
  assign mux_167_nl = or_tmp_386 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) nand_tmp_13 : mux_166_nl;
  assign mux_166_nl = or_1050_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) mux_165_nl : mux_164_nl;
  assign mux_165_nl = or_391_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) nand_tmp_13 : not_tmp_157;
  assign mux_164_nl = or_381_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) nand_tmp_13 : not_tmp_157;
  assign mux_144_nl = or_1087_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) or_tmp_312 : or_tmp_309;
  assign mux_140_nl = or_1087_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) main_stage_v_3 : main_stage_v_4;
  assign mux_129_nl = or_1087_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) or_tmp_269 : or_288_nl;
  assign mux_126_nl = FpAlu_8U_23U_equal_tmp_25 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) mux_125_nl : or_275_nl;
  assign mux_125_nl = or_1087_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) or_tmp_251 : or_273_nl;
  assign mux_124_nl = or_1087_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) or_tmp_251 : or_270_nl;
  assign AluIn_data_mux1h_13_itm = mux_334_nl ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16515|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16514" *) AluIn_data_sva_3_30_0_1 : { 8'b00000000, else_AluOp_data_else_AluOp_data_mux_4_nl };
  assign mux_334_nl = IsNaN_8U_23U_land_1_lpi_1_dfm_10 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) or_747_nl : mux_333_nl;
  assign mux_333_nl = IsNaN_8U_23U_land_1_lpi_1_dfm_11 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) or_tmp_657 : mux_tmp_311;
  assign else_AluOp_data_else_AluOp_data_mux_4_nl = and_204_nl ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16481|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16480" *) FpAdd_8U_23U_FpAdd_8U_23U_or_7_nl : else_AluOp_data_slc_else_AluOp_data_0_22_0_2_itm_2;
  assign FpAdd_8U_23U_FpAdd_8U_23U_or_7_nl = FpAdd_8U_23U_is_inf_mux_nl ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16481|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16480" *) 23'b11111111111111111111111 : alu_loop_op_1_FpMantRNE_49U_24U_else_acc_nl;
  assign FpAdd_8U_23U_is_inf_mux_nl = alu_loop_op_1_FpMantRNE_49U_24U_else_and_tmp ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) FpAdd_8U_23U_is_inf_1_lpi_1_dfm_2_mx0w0 : nor_33_cse;
  assign AluIn_data_mux1h_11_itm = mux_332_nl ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16515|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16514" *) AluIn_data_sva_3_62_32_1 : { 8'b00000000, else_AluOp_data_else_AluOp_data_mux_5_nl };
  assign mux_332_nl = IsNaN_8U_23U_land_2_lpi_1_dfm_10 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) or_744_nl : mux_331_nl;
  assign mux_331_nl = IsNaN_8U_23U_land_2_lpi_1_dfm_11 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) or_tmp_657 : mux_tmp_311;
  assign else_AluOp_data_else_AluOp_data_mux_5_nl = and_200_nl ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16481|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16480" *) FpAdd_8U_23U_FpAdd_8U_23U_or_6_nl : else_AluOp_data_slc_else_AluOp_data_1_22_0_7_itm_2;
  assign FpAdd_8U_23U_FpAdd_8U_23U_or_6_nl = FpAdd_8U_23U_is_inf_mux_1_nl ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16481|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16480" *) 23'b11111111111111111111111 : alu_loop_op_2_FpMantRNE_49U_24U_else_acc_2_nl;
  assign FpAdd_8U_23U_is_inf_mux_1_nl = alu_loop_op_2_FpMantRNE_49U_24U_else_and_2_tmp ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) FpAdd_8U_23U_is_inf_2_lpi_1_dfm_2_mx0w0 : nor_37_cse;
  assign AluIn_data_mux1h_9_itm = mux_330_nl ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16515|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16514" *) AluIn_data_sva_3_94_64_1 : { 8'b00000000, else_AluOp_data_else_AluOp_data_mux_6_nl };
  assign mux_330_nl = IsNaN_8U_23U_land_3_lpi_1_dfm_10 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) or_741_nl : mux_329_nl;
  assign mux_329_nl = IsNaN_8U_23U_land_3_lpi_1_dfm_11 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) or_tmp_657 : mux_tmp_311;
  assign else_AluOp_data_else_AluOp_data_mux_6_nl = and_196_nl ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16481|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16480" *) FpAdd_8U_23U_FpAdd_8U_23U_or_5_nl : else_AluOp_data_slc_else_AluOp_data_2_22_0_7_itm_2;
  assign FpAdd_8U_23U_FpAdd_8U_23U_or_5_nl = FpAdd_8U_23U_is_inf_mux_2_nl ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16481|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16480" *) 23'b11111111111111111111111 : alu_loop_op_3_FpMantRNE_49U_24U_else_acc_1_nl;
  assign FpAdd_8U_23U_is_inf_mux_2_nl = alu_loop_op_3_FpMantRNE_49U_24U_else_and_1_tmp ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) FpAdd_8U_23U_is_inf_3_lpi_1_dfm_2_mx0w0 : nor_41_cse;
  assign mux_111_nl = or_236_nl ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) or_239_nl : mux_110_nl;
  assign mux_110_nl = or_1087_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) or_tmp_75 : or_tmp_224;
  assign mux_107_nl = or_1087_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) mux_105_nl : nor_292_nl;
  assign mux_106_nl = or_225_nl ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) FpAlu_8U_23U_equal_tmp_23 : nor_293_nl;
  assign mux_105_nl = FpAlu_8U_23U_equal_tmp_22 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) nor_290_nl : nor_291_nl;
  assign AluIn_data_mux1h_7_itm = mux_328_nl ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16515|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16514" *) AluIn_data_sva_3_126_96_1 : { 8'b00000000, else_AluOp_data_else_AluOp_data_mux_7_nl };
  assign mux_328_nl = IsNaN_8U_23U_land_lpi_1_dfm_10 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) or_735_nl : mux_327_nl;
  assign mux_327_nl = IsNaN_8U_23U_land_lpi_1_dfm_11 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) or_tmp_657 : mux_tmp_311;
  assign else_AluOp_data_else_AluOp_data_mux_7_nl = and_192_nl ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16481|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16480" *) FpAdd_8U_23U_FpAdd_8U_23U_or_4_nl : else_AluOp_data_slc_else_AluOp_data_3_22_0_12_itm_2;
  assign FpAdd_8U_23U_FpAdd_8U_23U_or_4_nl = FpAdd_8U_23U_is_inf_mux_3_nl ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16481|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16480" *) 23'b11111111111111111111111 : alu_loop_op_4_FpMantRNE_49U_24U_else_acc_3_nl;
  assign FpAdd_8U_23U_is_inf_mux_3_nl = alu_loop_op_4_FpMantRNE_49U_24U_else_and_3_tmp ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) FpAdd_8U_23U_is_inf_lpi_1_dfm_2_mx0w0 : nor_45_cse;
  assign mux_46_nl = main_stage_v_1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) mux_45_nl : not_tmp_38;
  assign mux_45_nl = or_16_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) mux_44_nl : not_tmp_38;
  assign mux_44_nl = or_1087_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) and_dcpl_4 : main_stage_v_2;
  assign mux_43_nl = or_1087_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) nor_367_nl : nor_368_nl;
  assign cfg_alu_algo_cfg_alu_algo_mux_3_itm = and_dcpl_81 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16498|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16497" *) cfg_alu_algo_1_sva_st_20 : cfg_alu_algo_rsci_d;
  assign mux_15_nl = main_stage_v_1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) nand_nl : and_502_nl;
  assign _0431_ = and_328_rgt ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) alu_loop_op_1_FpAdd_8U_23U_IsZero_8U_23U_or_itm_mx0w2 : IsNaN_8U_23U_2_nor_3_mx0w0;
  assign _0218_ = _0881_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15534" *) _0431_ : IsNaN_8U_23U_4_nor_3_itm_2;
  assign _0211_ = IsNaN_8U_23U_2_and_9_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15518" *) _2328_ : IsNaN_8U_23U_2_IsNaN_8U_23U_2_nor_2_itm;
  assign _0209_ = IsNaN_8U_23U_2_and_9_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15518" *) _2329_ : IsNaN_8U_23U_2_IsNaN_8U_23U_2_nor_1_itm;
  assign _0215_ = IsNaN_8U_23U_2_and_9_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15518" *) _2330_ : IsNaN_8U_23U_2_IsNaN_8U_23U_2_nor_itm;
  assign _0213_ = _0879_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15506" *) _2327_ : IsNaN_8U_23U_2_IsNaN_8U_23U_2_nor_3_itm;
  assign _0217_ = _0878_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15495" *) _2356_ : IsNaN_8U_23U_4_nor_2_itm_2;
  assign _0219_ = _0877_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15484" *) _2355_ : IsNaN_8U_23U_4_nor_3_itm_3;
  assign _0157_ = _0875_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15475" *) FpCmp_8U_23U_false_is_abs_a_greater_2_lpi_1_dfm_1_mx0w0 : FpCmp_8U_23U_false_is_abs_a_greater_2_lpi_1_dfm_2;
  assign _0212_ = IsNaN_8U_23U_2_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15458" *) _2353_ : IsNaN_8U_23U_2_IsNaN_8U_23U_2_nor_2_itm_1;
  assign _0210_ = IsNaN_8U_23U_2_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15458" *) _2354_ : IsNaN_8U_23U_2_IsNaN_8U_23U_2_nor_1_itm_1;
  assign _0214_ = IsNaN_8U_23U_2_and_6_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15442" *) _2351_ : IsNaN_8U_23U_2_IsNaN_8U_23U_2_nor_3_itm_2;
  assign _0216_ = IsNaN_8U_23U_2_and_6_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15442" *) _2352_ : IsNaN_8U_23U_2_IsNaN_8U_23U_2_nor_itm_2;
  assign _0266_ = _0873_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15432" *) cfg_alu_src_rsci_d : alu_loop_op_2_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_1_svs_2;
  assign _0146_ = FpAlu_8U_23U_and_102_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15411" *) _2374_ : FpAlu_8U_23U_mux1h_152_itm_2;
  assign _0147_ = FpAlu_8U_23U_and_102_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15411" *) _2373_ : FpAlu_8U_23U_mux1h_33_itm_2;
  assign _0293_ = IntSaturation_33U_32U_if_and_9_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15397" *) alu_loop_op_4_IntSaturation_33U_32U_if_acc_1_nl[2] : alu_loop_op_4_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_1_svs_2;
  assign _0254_ = IntSaturation_33U_32U_if_and_9_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15397" *) alu_loop_op_1_IntSaturation_33U_32U_if_acc_nl[2] : alu_loop_op_1_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_svs_2;
  assign _0280_ = IntSaturation_33U_32U_if_and_9_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15397" *) alu_loop_op_3_IntSaturation_33U_32U_if_acc_nl[2] : alu_loop_op_3_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_svs_2;
  assign _0385_ = _0872_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15384" *) alu_loop_op_else_o_mux1h_7_itm[30:0] : reg_alu_loop_op_else_o_32_1_lpi_1_dfm_4_1_itm;
  assign _0386_ = _0864_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15372" *) alu_loop_op_else_o_mux1h_7_itm[31] : reg_alu_loop_op_else_o_32_1_lpi_1_dfm_4_itm;
  assign _0383_ = _0856_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15362" *) alu_loop_op_else_o_mux1h_5_itm[30:0] : reg_alu_loop_op_else_o_32_1_3_lpi_1_dfm_3_1_itm;
  assign _0384_ = _0847_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15351" *) alu_loop_op_else_o_mux1h_5_itm[31] : reg_alu_loop_op_else_o_32_1_3_lpi_1_dfm_3_itm;
  assign _0430_ = and_293_rgt ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) alu_loop_op_2_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_1_svs_2 : alu_loop_op_2_IntSaturation_33U_32U_if_acc_1_nl[2];
  assign _0267_ = _0838_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15338" *) _0430_ : alu_loop_op_2_IntSaturation_33U_32U_if_slc_IntSaturation_33U_32U_if_acc_2_1_svs_3;
  assign _0381_ = _0835_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15328" *) alu_loop_op_else_o_mux1h_3_itm[30:0] : reg_alu_loop_op_else_o_32_1_2_lpi_1_dfm_4_1_itm;
  assign _0382_ = _0828_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15318" *) alu_loop_op_else_o_mux1h_3_itm[31] : reg_alu_loop_op_else_o_32_1_2_lpi_1_dfm_4_itm;
  assign _0379_ = _0819_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15307" *) alu_loop_op_else_o_mux1h_1_itm[30:0] : reg_alu_loop_op_else_o_32_1_1_lpi_1_dfm_3_1_itm;
  assign _0380_ = _0812_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15297" *) alu_loop_op_else_o_mux1h_1_itm[31] : reg_alu_loop_op_else_o_32_1_1_lpi_1_dfm_3_itm;
  assign _0143_ = _0802_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15286" *) FpAlu_8U_23U_equal_tmp_2_mx0w0 : FpAlu_8U_23U_equal_tmp_33;
  assign _0140_ = _0801_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15278" *) FpAlu_8U_23U_equal_tmp_2_mx0w0 : FpAlu_8U_23U_equal_tmp_30;
  assign _0166_ = FpCmp_8U_23U_true_o_and_9_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15268" *) FpCmp_8U_23U_true_o_1_lpi_1_dfm_1_mx0[30:0] : FpCmp_8U_23U_true_o_1_lpi_1_dfm_5_30_0_1;
  assign _0169_ = FpCmp_8U_23U_true_o_and_9_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15268" *) FpCmp_8U_23U_true_o_2_lpi_1_dfm_1_mx0[30:0] : FpCmp_8U_23U_true_o_2_lpi_1_dfm_5_30_0_1;
  assign _0172_ = FpCmp_8U_23U_true_o_and_9_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15268" *) FpCmp_8U_23U_true_o_3_lpi_1_dfm_1_mx0[30:0] : FpCmp_8U_23U_true_o_3_lpi_1_dfm_5_30_0_1;
  assign _0175_ = _0800_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15258" *) FpCmp_8U_23U_true_o_lpi_1_dfm_1_mx0[30:0] : FpCmp_8U_23U_true_o_lpi_1_dfm_5_30_0_1;
  assign _0065_ = AluOut_data_and_17_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15245" *) _2326_ : AluOut_data_0_0_sva_9;
  assign _0066_ = AluOut_data_and_17_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15245" *) _2325_ : AluOut_data_1_0_sva_10;
  assign _0072_ = _0799_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15236" *) AluOut_data_2_0_sva_3_mx0w0 : AluOut_data_2_0_sva_9;
  assign _0152_ = _0798_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15228" *) FpAlu_8U_23U_o_0_sva_2_mx0w0 : FpAlu_8U_23U_o_0_sva_7;
  assign _0223_ = IsNaN_8U_23U_aelse_and_16_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15217" *) IsNaN_8U_23U_land_1_lpi_1_dfm_8 : IsNaN_8U_23U_land_1_lpi_1_dfm_9;
  assign _0229_ = IsNaN_8U_23U_aelse_and_16_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15217" *) IsNaN_8U_23U_land_2_lpi_1_dfm_8 : IsNaN_8U_23U_land_2_lpi_1_dfm_9;
  assign _0235_ = IsNaN_8U_23U_aelse_and_16_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15217" *) IsNaN_8U_23U_land_3_lpi_1_dfm_8 : IsNaN_8U_23U_land_3_lpi_1_dfm_9;
  assign _0241_ = IsNaN_8U_23U_aelse_and_16_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15217" *) IsNaN_8U_23U_land_lpi_1_dfm_8 : IsNaN_8U_23U_land_lpi_1_dfm_9;
  assign _0283_ = IsZero_8U_23U_and_6_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15204" *) alu_loop_op_4_FpAdd_8U_23U_IsZero_8U_23U_or_itm_mx0w0 : alu_loop_op_4_FpAdd_8U_23U_IsZero_8U_23U_or_itm_3;
  assign _0270_ = IsZero_8U_23U_and_6_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15204" *) alu_loop_op_3_FpAdd_8U_23U_IsZero_8U_23U_or_itm_mx0w0 : alu_loop_op_3_FpAdd_8U_23U_IsZero_8U_23U_or_itm_3;
  assign _0257_ = IsZero_8U_23U_and_6_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15204" *) alu_loop_op_2_FpAdd_8U_23U_IsZero_8U_23U_or_itm_mx0w0 : alu_loop_op_2_FpAdd_8U_23U_IsZero_8U_23U_or_itm_3;
  assign _0459_ = FpAdd_8U_23U_qr_lpi_1_dfm_mx0c1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16600|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16599" *) else_AluOp_data_3_lpi_1_dfm_mx1_tmp_30_23 : AluIn_data_sva_127[126:119];
  assign _0126_ = _0797_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15193" *) _0459_ : FpAdd_8U_23U_qr_lpi_1_dfm;
  assign _0458_ = FpAdd_8U_23U_qr_4_lpi_1_dfm_mx0c1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16600|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16599" *) else_AluOp_data_2_lpi_1_dfm_mx1_tmp_30_23 : AluIn_data_sva_127[94:87];
  assign _0123_ = _0794_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15183" *) _0458_ : FpAdd_8U_23U_qr_4_lpi_1_dfm;
  assign _0457_ = FpAdd_8U_23U_qr_3_lpi_1_dfm_mx0c1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16600|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16599" *) else_AluOp_data_1_lpi_1_dfm_mx1_tmp_30_23 : AluIn_data_sva_127[62:55];
  assign _0120_ = _0791_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15173" *) _0457_ : FpAdd_8U_23U_qr_3_lpi_1_dfm;
  assign _0456_ = FpAdd_8U_23U_qr_2_lpi_1_dfm_mx0c1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16600|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16599" *) else_AluOp_data_0_lpi_1_dfm_mx1_tmp_30_23 : AluIn_data_sva_127[30:23];
  assign _0117_ = _0788_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15163" *) _0456_ : FpAdd_8U_23U_qr_2_lpi_1_dfm;
  assign _0129_ = FpAlu_8U_23U_and_94_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15149" *) _0784_ : FpAlu_8U_23U_and_3_itm_2;
  assign _0130_ = FpAlu_8U_23U_and_94_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15149" *) _0785_ : FpAlu_8U_23U_and_6_itm_2;
  assign _0137_ = FpAlu_8U_23U_and_94_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15149" *) FpAlu_8U_23U_equal_tmp_2_mx0w0 : FpAlu_8U_23U_equal_tmp_27;
  assign _0148_ = FpAlu_8U_23U_and_94_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15149" *) FpAlu_8U_23U_nor_dfs_mx0w0 : FpAlu_8U_23U_nor_dfs_4;
  assign _0134_ = FpAlu_8U_23U_and_94_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15149" *) FpAlu_8U_23U_equal_tmp_mx0w0 : FpAlu_8U_23U_equal_tmp_24;
  assign _0131_ = FpAlu_8U_23U_and_94_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15149" *) FpAlu_8U_23U_equal_tmp_1_mx0w0 : FpAlu_8U_23U_equal_tmp_21;
  assign _0343_ = FpAdd_8U_23U_int_mant_p1_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15133" *) else_AluOp_data_2_lpi_1_dfm_2_30_0_1[30:23] : else_AluOp_data_slc_else_AluOp_data_2_30_23_21_itm;
  assign _0339_ = FpAdd_8U_23U_int_mant_p1_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15133" *) else_AluOp_data_1_lpi_1_dfm_2_30_0_1[30:23] : else_AluOp_data_slc_else_AluOp_data_1_30_23_21_itm;
  assign _0335_ = FpAdd_8U_23U_int_mant_p1_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15133" *) else_AluOp_data_0_lpi_1_dfm_2_30_0_1[30:23] : else_AluOp_data_slc_else_AluOp_data_0_30_23_7_itm;
  assign _0347_ = FpAdd_8U_23U_int_mant_p1_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15133" *) else_AluOp_data_3_lpi_1_dfm_2_30_0_1[30:23] : else_AluOp_data_slc_else_AluOp_data_3_30_23_35_itm;
  assign _0345_ = _0783_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15122" *) else_AluOp_data_3_lpi_1_dfm_2_30_0_1[22:0] : else_AluOp_data_slc_else_AluOp_data_3_22_0_12_itm;
  assign _0341_ = _0782_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15113" *) else_AluOp_data_2_lpi_1_dfm_2_30_0_1[22:0] : else_AluOp_data_slc_else_AluOp_data_2_22_0_7_itm;
  assign _0337_ = _0781_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15104" *) else_AluOp_data_1_lpi_1_dfm_2_30_0_1[22:0] : else_AluOp_data_slc_else_AluOp_data_1_22_0_7_itm;
  assign _0333_ = _0780_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15095" *) else_AluOp_data_0_lpi_1_dfm_2_30_0_1[22:0] : else_AluOp_data_slc_else_AluOp_data_0_22_0_2_itm;
  assign _0436_ = and_dcpl_99 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16481|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16480" *) else_AluOp_data_slc_else_AluOp_data_3_22_0_12_itm : else_AluOp_data_3_lpi_1_dfm_2_30_0_1[22:0];
  assign _0346_ = _0779_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15085" *) _0436_ : else_AluOp_data_slc_else_AluOp_data_3_22_0_12_itm_2;
  assign _0435_ = and_dcpl_99 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16481|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16480" *) else_AluOp_data_slc_else_AluOp_data_2_22_0_7_itm : else_AluOp_data_2_lpi_1_dfm_2_30_0_1[22:0];
  assign _0342_ = _0778_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15075" *) _0435_ : else_AluOp_data_slc_else_AluOp_data_2_22_0_7_itm_2;
  assign _0434_ = and_dcpl_99 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16481|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16480" *) else_AluOp_data_slc_else_AluOp_data_1_22_0_7_itm : else_AluOp_data_1_lpi_1_dfm_2_30_0_1[22:0];
  assign _0338_ = _0777_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15065" *) _0434_ : else_AluOp_data_slc_else_AluOp_data_1_22_0_7_itm_2;
  assign _0433_ = and_dcpl_99 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16481|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16480" *) else_AluOp_data_slc_else_AluOp_data_0_22_0_2_itm : else_AluOp_data_0_lpi_1_dfm_2_30_0_1[22:0];
  assign _0334_ = _0776_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15055" *) _0433_ : else_AluOp_data_slc_else_AluOp_data_0_22_0_2_itm_2;
  assign _0361_ = AluOut_data_and_15_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15035" *) _2324_ : mux_177_itm_3;
  assign _0363_ = AluOut_data_and_15_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15035" *) _2323_ : mux_181_itm_3;
  assign _0365_ = AluOut_data_and_15_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15035" *) _2322_ : mux_189_itm_3;
  assign _0075_ = AluOut_data_and_15_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15035" *) _2321_ : AluOut_data_2_31_lpi_1_dfm_6;
  assign _0187_ = _0775_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15022" *) _2415_ : IntSaturation_33U_32U_slc_IntSaturation_33U_32U_o_31_1_1_29_22_itm_2;
  assign _0193_ = _0774_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15011" *) _2414_ : IntSaturation_33U_32U_slc_IntSaturation_33U_32U_o_31_1_2_29_22_itm_3;
  assign _0190_ = _0773_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:15000" *) _2413_ : IntSaturation_33U_32U_slc_IntSaturation_33U_32U_o_31_1_29_22_itm_3;
  assign _0186_ = IntSaturation_33U_32U_and_11_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14988" *) IntSaturation_33U_32U_o_31_1_1_lpi_1_dfm_1[21:0] : IntSaturation_33U_32U_slc_IntSaturation_33U_32U_o_31_1_1_21_0_itm_2;
  assign _0191_ = IntSaturation_33U_32U_and_11_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14988" *) IntSaturation_33U_32U_o_31_1_2_lpi_1_dfm_1[21:0] : IntSaturation_33U_32U_slc_IntSaturation_33U_32U_o_31_1_2_21_0_itm_3;
  assign _0188_ = IntSaturation_33U_32U_and_11_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14988" *) IntSaturation_33U_32U_o_31_1_lpi_1_dfm_1[21:0] : IntSaturation_33U_32U_slc_IntSaturation_33U_32U_o_31_1_21_0_itm_3;
  assign _0194_ = IntSaturation_33U_32U_and_11_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14988" *) IntSaturation_33U_32U_o_31_1_3_lpi_1_dfm_1[21:0] : IntSaturation_33U_32U_slc_IntSaturation_33U_32U_o_31_1_3_21_0_itm_3;
  assign _0196_ = _0772_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14975" *) _2412_ : IntSaturation_33U_32U_slc_IntSaturation_33U_32U_o_31_1_3_29_22_itm_3;
  assign _0144_ = _0770_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14966" *) FpAlu_8U_23U_equal_tmp_33 : FpAlu_8U_23U_equal_tmp_34;
  assign _0158_ = FpCmp_8U_23U_false_o_and_6_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14957" *) reg_alu_loop_op_else_o_32_1_1_lpi_1_dfm_3_1_itm : FpCmp_8U_23U_false_o_1_lpi_1_dfm_6_30_0_1;
  assign _0160_ = FpCmp_8U_23U_false_o_and_6_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14957" *) reg_alu_loop_op_else_o_32_1_2_lpi_1_dfm_4_1_itm : FpCmp_8U_23U_false_o_2_lpi_1_dfm_7_30_0_1;
  assign _0162_ = _0769_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14948" *) reg_alu_loop_op_else_o_32_1_3_lpi_1_dfm_3_1_itm : FpCmp_8U_23U_false_o_3_lpi_1_dfm_7_30_0_1;
  assign _0164_ = _0768_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14940" *) reg_alu_loop_op_else_o_32_1_lpi_1_dfm_4_1_itm : FpCmp_8U_23U_false_o_lpi_1_dfm_8_30_0_1;
  assign _0167_ = FpCmp_8U_23U_true_o_and_5_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14930" *) FpCmp_8U_23U_true_o_1_lpi_1_dfm_5_30_0_1 : FpCmp_8U_23U_true_o_1_lpi_1_dfm_6_30_0_1;
  assign _0170_ = FpCmp_8U_23U_true_o_and_5_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14930" *) FpCmp_8U_23U_true_o_2_lpi_1_dfm_5_30_0_1 : FpCmp_8U_23U_true_o_2_lpi_1_dfm_6_30_0_1;
  assign _0173_ = FpCmp_8U_23U_true_o_and_5_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14930" *) FpCmp_8U_23U_true_o_3_lpi_1_dfm_5_30_0_1 : FpCmp_8U_23U_true_o_3_lpi_1_dfm_6_30_0_1;
  assign _0176_ = _0767_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14920" *) FpCmp_8U_23U_true_o_lpi_1_dfm_5_30_0_1 : FpCmp_8U_23U_true_o_lpi_1_dfm_6_30_0_1;
  assign _0141_ = FpAlu_8U_23U_and_88_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14908" *) FpAlu_8U_23U_equal_tmp_30 : FpAlu_8U_23U_equal_tmp_31;
  assign _0138_ = FpAlu_8U_23U_and_88_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14908" *) FpAlu_8U_23U_equal_tmp_27 : FpAlu_8U_23U_equal_tmp_28;
  assign _0149_ = FpAlu_8U_23U_and_88_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14908" *) FpAlu_8U_23U_nor_dfs_4 : FpAlu_8U_23U_nor_dfs_5;
  assign _0135_ = FpAlu_8U_23U_and_88_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14908" *) FpAlu_8U_23U_equal_tmp_24 : FpAlu_8U_23U_equal_tmp_25;
  assign _0132_ = FpAlu_8U_23U_and_88_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14908" *) FpAlu_8U_23U_equal_tmp_21 : FpAlu_8U_23U_equal_tmp_22;
  assign _0429_ = and_dcpl_165 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) IntSaturation_33U_32U_IntSaturation_33U_32U_or_1_nl : AluOut_data_0_0_sva_9;
  assign _0428_ = and_dcpl_165 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) IntSaturation_33U_32U_IntSaturation_33U_32U_or_2_nl : AluOut_data_1_0_sva_10;
  assign _0427_ = and_dcpl_165 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) IntSaturation_33U_32U_IntSaturation_33U_32U_or_3_nl : AluOut_data_2_0_sva_9;
  assign _0063_ = AluOut_data_and_12_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14891" *) _0429_ : AluOut_data_0_0_sva_10;
  assign _0067_ = AluOut_data_and_12_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14891" *) _0428_ : AluOut_data_1_0_sva_11;
  assign _0070_ = AluOut_data_and_12_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14891" *) _0427_ : AluOut_data_2_0_sva_10;
  assign _0426_ = and_dcpl_165 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) IntSaturation_33U_32U_IntSaturation_33U_32U_or_nl : FpAlu_8U_23U_o_0_sva_7;
  assign _0153_ = _0766_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14880" *) _0426_ : FpAlu_8U_23U_o_0_sva_8;
  assign _0220_ = IsNaN_8U_23U_aelse_and_12_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14868" *) IsNaN_8U_23U_land_1_lpi_1_dfm_9 : IsNaN_8U_23U_land_1_lpi_1_dfm_10;
  assign _0226_ = IsNaN_8U_23U_aelse_and_12_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14868" *) IsNaN_8U_23U_land_2_lpi_1_dfm_9 : IsNaN_8U_23U_land_2_lpi_1_dfm_10;
  assign _0232_ = IsNaN_8U_23U_aelse_and_12_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14868" *) IsNaN_8U_23U_land_3_lpi_1_dfm_9 : IsNaN_8U_23U_land_3_lpi_1_dfm_10;
  assign _0238_ = IsNaN_8U_23U_aelse_and_12_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14868" *) IsNaN_8U_23U_land_lpi_1_dfm_9 : IsNaN_8U_23U_land_lpi_1_dfm_10;
  assign _0127_ = _0765_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14854" *) _2411_ : FpAdd_8U_23U_qr_lpi_1_dfm_6;
  assign _0124_ = _0763_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14843" *) _2410_ : FpAdd_8U_23U_qr_4_lpi_1_dfm_6;
  assign _0121_ = _0761_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14832" *) _2409_ : FpAdd_8U_23U_qr_3_lpi_1_dfm_6;
  assign _0118_ = _0759_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14821" *) _2408_ : FpAdd_8U_23U_qr_2_lpi_1_dfm_6;
  assign _0297_ = _0757_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14813" *) cfg_alu_algo_rsci_d : cfg_alu_algo_1_sva_2;
  assign _0306_ = _0756_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14805" *) cfg_alu_src_rsci_d : cfg_alu_src_1_sva_st;
  assign _0298_ = _0755_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14796" *) cfg_alu_algo_rsci_d : cfg_alu_algo_1_sva_st;
  assign _0299_ = _0754_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14788" *) cfg_alu_algo_rsci_d : cfg_alu_algo_1_sva_st_20;
  assign _0288_ = FpAdd_8U_23U_is_addition_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14773" *) alu_loop_op_4_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_3_svs_mx0w0 : alu_loop_op_4_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_3_svs_st;
  assign _0275_ = FpAdd_8U_23U_is_addition_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14773" *) alu_loop_op_3_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_1_svs_mx0w0 : alu_loop_op_3_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_1_svs_st;
  assign _0261_ = FpAdd_8U_23U_is_addition_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14773" *) alu_loop_op_2_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_2_svs_mx0w0 : alu_loop_op_2_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_2_svs_st;
  assign _0249_ = FpAdd_8U_23U_is_addition_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14773" *) alu_loop_op_1_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_mx0w0 : alu_loop_op_1_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_st;
  assign _0281_ = IsZero_8U_23U_1_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14747" *) alu_loop_op_4_FpAdd_8U_23U_IsZero_8U_23U_1_or_itm_mx0w0 : alu_loop_op_4_FpAdd_8U_23U_IsZero_8U_23U_1_or_itm;
  assign _0268_ = IsZero_8U_23U_1_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14747" *) alu_loop_op_3_FpAdd_8U_23U_IsZero_8U_23U_1_or_itm_mx0w0 : alu_loop_op_3_FpAdd_8U_23U_IsZero_8U_23U_1_or_itm;
  assign _0255_ = IsZero_8U_23U_1_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14747" *) alu_loop_op_2_FpAdd_8U_23U_IsZero_8U_23U_1_or_itm_mx0w0 : alu_loop_op_2_FpAdd_8U_23U_IsZero_8U_23U_1_or_itm;
  assign _0244_ = IsZero_8U_23U_1_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14747" *) alu_loop_op_1_FpAdd_8U_23U_IsZero_8U_23U_1_or_itm_mx0w0 : alu_loop_op_1_FpAdd_8U_23U_IsZero_8U_23U_1_or_itm;
  assign _0081_ = IsZero_8U_23U_1_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14747" *) FpAdd_8U_23U_a_right_shift_qr_3_lpi_1_dfm_mx0w0 : FpAdd_8U_23U_a_right_shift_qr_3_lpi_1_dfm;
  assign _0093_ = IsZero_8U_23U_1_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14747" *) FpAdd_8U_23U_b_right_shift_qr_3_lpi_1_dfm_mx0w0 : FpAdd_8U_23U_b_right_shift_qr_3_lpi_1_dfm;
  assign _0079_ = IsZero_8U_23U_1_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14747" *) FpAdd_8U_23U_a_right_shift_qr_2_lpi_1_dfm_mx0w0 : FpAdd_8U_23U_a_right_shift_qr_2_lpi_1_dfm;
  assign _0091_ = IsZero_8U_23U_1_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14747" *) FpAdd_8U_23U_b_right_shift_qr_2_lpi_1_dfm_mx0w0 : FpAdd_8U_23U_b_right_shift_qr_2_lpi_1_dfm;
  assign _0077_ = IsZero_8U_23U_1_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14747" *) FpAdd_8U_23U_a_right_shift_qr_1_lpi_1_dfm_mx0w0 : FpAdd_8U_23U_a_right_shift_qr_1_lpi_1_dfm;
  assign _0089_ = IsZero_8U_23U_1_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14747" *) FpAdd_8U_23U_b_right_shift_qr_1_lpi_1_dfm_mx0w0 : FpAdd_8U_23U_b_right_shift_qr_1_lpi_1_dfm;
  assign _0083_ = IsZero_8U_23U_1_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14747" *) FpAdd_8U_23U_a_right_shift_qr_lpi_1_dfm_mx0w0 : FpAdd_8U_23U_a_right_shift_qr_lpi_1_dfm;
  assign _0095_ = IsZero_8U_23U_1_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14747" *) FpAdd_8U_23U_b_right_shift_qr_lpi_1_dfm_mx0w0 : FpAdd_8U_23U_b_right_shift_qr_lpi_1_dfm;
  assign _0425_ = and_dcpl_81 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) alu_loop_op_3_FpAdd_8U_23U_IsZero_8U_23U_or_itm_3 : alu_loop_op_3_FpAdd_8U_23U_IsZero_8U_23U_or_itm_mx0w0;
  assign _0424_ = and_dcpl_81 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) alu_loop_op_4_FpAdd_8U_23U_IsZero_8U_23U_or_itm_3 : alu_loop_op_4_FpAdd_8U_23U_IsZero_8U_23U_or_itm_mx0w0;
  assign _0284_ = IsZero_8U_23U_and_4_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14725" *) _0424_ : alu_loop_op_4_FpAdd_8U_23U_IsZero_8U_23U_or_itm_4;
  assign _0271_ = IsZero_8U_23U_and_4_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14725" *) _0425_ : alu_loop_op_3_FpAdd_8U_23U_IsZero_8U_23U_or_itm_4;
  assign _0289_ = FpAdd_8U_23U_if_3_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14713" *) acc_15_nl[50] : alu_loop_op_4_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_3_itm;
  assign _0276_ = FpAdd_8U_23U_if_3_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14713" *) acc_14_nl[50] : alu_loop_op_3_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_1_itm;
  assign _0262_ = FpAdd_8U_23U_if_3_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14713" *) acc_13_nl[50] : alu_loop_op_2_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_2_itm;
  assign _0250_ = FpAdd_8U_23U_if_3_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14713" *) acc_12_nl[50] : alu_loop_op_1_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_itm;
  assign _0182_ = _0753_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14702" *) FpNormalize_8U_49U_if_or_3_itm_mx0w0 : FpNormalize_8U_49U_if_or_3_itm;
  assign _0180_ = _0752_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14694" *) FpNormalize_8U_49U_if_or_2_itm_mx0w0 : FpNormalize_8U_49U_if_or_2_itm;
  assign _0178_ = _0751_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14686" *) FpNormalize_8U_49U_if_or_1_itm_mx0w0 : FpNormalize_8U_49U_if_or_1_itm;
  assign _0103_ = FpAdd_8U_23U_int_mant_p1_and_12_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14675" *) acc_15_nl[50:1] : FpAdd_8U_23U_int_mant_p1_lpi_1_dfm;
  assign _0101_ = FpAdd_8U_23U_int_mant_p1_and_12_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14675" *) acc_14_nl[50:1] : FpAdd_8U_23U_int_mant_p1_3_lpi_1_dfm;
  assign _0099_ = FpAdd_8U_23U_int_mant_p1_and_12_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14675" *) acc_13_nl[50:1] : FpAdd_8U_23U_int_mant_p1_2_lpi_1_dfm;
  assign _0097_ = FpAdd_8U_23U_int_mant_p1_and_12_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14675" *) acc_12_nl[50:1] : FpAdd_8U_23U_int_mant_p1_1_lpi_1_dfm;
  assign _0184_ = _0750_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14664" *) FpNormalize_8U_49U_if_or_itm_mx0w0 : FpNormalize_8U_49U_if_or_itm;
  assign _0207_ = _0748_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14656" *) IsNaN_8U_23U_1_land_lpi_1_dfm_7 : IsNaN_8U_23U_1_land_lpi_1_dfm_8;
  assign _0204_ = _0747_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14648" *) IsNaN_8U_23U_1_land_3_lpi_1_dfm_7 : IsNaN_8U_23U_1_land_3_lpi_1_dfm_8;
  assign _0201_ = _0746_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14640" *) IsNaN_8U_23U_1_land_2_lpi_1_dfm_7 : IsNaN_8U_23U_1_land_2_lpi_1_dfm_8;
  assign _0198_ = _0745_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14632" *) IsNaN_8U_23U_1_land_1_lpi_1_dfm_7 : IsNaN_8U_23U_1_land_1_lpi_1_dfm_8;
  assign _0291_ = FpMantRNE_49U_24U_else_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14621" *) alu_loop_op_4_FpMantRNE_49U_24U_else_and_3_tmp : alu_loop_op_4_FpMantRNE_49U_24U_else_and_3_svs_st;
  assign _0278_ = FpMantRNE_49U_24U_else_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14621" *) alu_loop_op_3_FpMantRNE_49U_24U_else_and_1_tmp : alu_loop_op_3_FpMantRNE_49U_24U_else_and_1_svs_st;
  assign _0264_ = FpMantRNE_49U_24U_else_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14621" *) alu_loop_op_2_FpMantRNE_49U_24U_else_and_2_tmp : alu_loop_op_2_FpMantRNE_49U_24U_else_and_2_svs_st;
  assign _0252_ = FpMantRNE_49U_24U_else_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14621" *) alu_loop_op_1_FpMantRNE_49U_24U_else_and_tmp : alu_loop_op_1_FpMantRNE_49U_24U_else_and_svs_st;
  assign _0286_ = _0744_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14609" *) alu_loop_op_4_FpAdd_8U_23U_if_4_if_acc_6_nl[7] : alu_loop_op_4_FpAdd_8U_23U_if_4_if_slc_FpAdd_8U_23U_if_4_if_acc_1_7_3_svs_st_2;
  assign _0273_ = _0743_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14599" *) alu_loop_op_3_FpAdd_8U_23U_if_4_if_acc_2_nl[7] : alu_loop_op_3_FpAdd_8U_23U_if_4_if_slc_FpAdd_8U_23U_if_4_if_acc_1_7_1_svs_st_2;
  assign _0259_ = _0742_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14589" *) alu_loop_op_2_FpAdd_8U_23U_if_4_if_acc_4_nl[7] : alu_loop_op_2_FpAdd_8U_23U_if_4_if_slc_FpAdd_8U_23U_if_4_if_acc_1_7_2_svs_st_2;
  assign _0247_ = _0741_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14579" *) alu_loop_op_1_FpAdd_8U_23U_if_4_if_acc_1_nl[7] : alu_loop_op_1_FpAdd_8U_23U_if_4_if_slc_FpAdd_8U_23U_if_4_if_acc_1_7_svs_st_2;
  assign _0423_ = and_dcpl_108 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) FpAlu_8U_23U_o_0_sva_8 : AluOut_data_2_0_sva_10;
  assign _0071_ = _0740_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14569" *) _0423_ : AluOut_data_2_0_sva_11;
  assign _0069_ = _0739_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14558" *) _2320_ : AluOut_data_2_0_lpi_1_dfm_3;
  assign _0192_ = IntSaturation_33U_32U_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14548" *) IntSaturation_33U_32U_slc_IntSaturation_33U_32U_o_31_1_2_21_0_itm_3 : IntSaturation_33U_32U_slc_IntSaturation_33U_32U_o_31_1_2_21_0_itm_4;
  assign _0189_ = IntSaturation_33U_32U_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14548" *) IntSaturation_33U_32U_slc_IntSaturation_33U_32U_o_31_1_21_0_itm_3 : IntSaturation_33U_32U_slc_IntSaturation_33U_32U_o_31_1_21_0_itm_4;
  assign _0195_ = IntSaturation_33U_32U_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14548" *) IntSaturation_33U_32U_slc_IntSaturation_33U_32U_o_31_1_3_21_0_itm_3 : IntSaturation_33U_32U_slc_IntSaturation_33U_32U_o_31_1_3_21_0_itm_4;
  assign _0064_ = AluOut_data_and_8_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14537" *) AluOut_data_0_0_sva_10 : AluOut_data_0_0_sva_11;
  assign _0068_ = AluOut_data_and_8_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14537" *) AluOut_data_1_0_sva_11 : AluOut_data_1_0_sva_12;
  assign _0356_ = and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14522" *) io_read_cfg_alu_bypass_rsc_svs_st_6 : io_read_cfg_alu_bypass_rsc_svs_st_7;
  assign _0362_ = and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14522" *) mux_177_itm_3 : mux_177_itm_4;
  assign _0364_ = and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14522" *) mux_181_itm_3 : mux_181_itm_4;
  assign _0366_ = and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14522" *) mux_189_itm_3 : mux_189_itm_4;
  assign _0076_ = and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14522" *) AluOut_data_2_31_lpi_1_dfm_6 : AluOut_data_2_31_lpi_1_dfm_7;
  assign _0352_ = and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14522" *) io_read_cfg_alu_bypass_rsc_svs_7 : io_read_cfg_alu_bypass_rsc_svs_8;
  assign _0296_ = and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14522" *) alu_loop_op_unequal_tmp_7 : alu_loop_op_unequal_tmp_8;
  assign _0303_ = _0738_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14508" *) cfg_alu_algo_1_sva_st_24 : cfg_alu_algo_1_sva_st_25;
  assign _0145_ = _0737_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14500" *) FpAlu_8U_23U_equal_tmp_34 : FpAlu_8U_23U_equal_tmp_35;
  assign _0348_ = _0736_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14492" *) IntSaturation_33U_32U_slc_IntSaturation_33U_32U_o_31_1_29_22_itm_3 : else_AluOp_data_slc_else_AluOp_data_3_30_23_35_itm_3;
  assign _0422_ = and_217_rgt ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) nor_45_cse : FpAdd_8U_23U_is_inf_lpi_1_dfm_2_mx0w0;
  assign _0112_ = _0735_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14483" *) _0422_ : FpAdd_8U_23U_is_inf_lpi_1_dfm_8;
  assign _0155_ = and_524_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14473" *) FpAlu_8U_23U_o_22_1_lpi_1_dfm_2 : FpAlu_8U_23U_o_22_1_lpi_1_dfm_4;
  assign _0156_ = and_524_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14473" *) FpAlu_8U_23U_o_30_23_lpi_1_dfm_2 : FpAlu_8U_23U_o_30_23_lpi_1_dfm_4;
  assign _0165_ = _0732_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14464" *) FpCmp_8U_23U_false_o_lpi_1_dfm_8_30_0_1 : FpCmp_8U_23U_false_o_lpi_1_dfm_9_30_0_1;
  assign _0151_ = _0731_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14456" *) FpAlu_8U_23U_o_0_lpi_1_dfm_2 : FpAlu_8U_23U_o_0_lpi_1_dfm_4;
  assign _0154_ = _0727_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14446" *) FpAlu_8U_23U_o_0_sva_8 : FpAlu_8U_23U_o_0_sva_9;
  assign _0177_ = _0726_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14438" *) FpCmp_8U_23U_true_o_lpi_1_dfm_6_30_0_1 : FpCmp_8U_23U_true_o_lpi_1_dfm_7_30_0_1;
  assign _0336_ = _0725_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14430" *) IntSaturation_33U_32U_slc_IntSaturation_33U_32U_o_31_1_1_29_22_itm_2 : else_AluOp_data_slc_else_AluOp_data_0_30_23_7_itm_3;
  assign _0421_ = and_215_rgt ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) nor_33_cse : FpAdd_8U_23U_is_inf_1_lpi_1_dfm_2_mx0w0;
  assign _0109_ = _0724_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14421" *) _0421_ : FpAdd_8U_23U_is_inf_1_lpi_1_dfm_8;
  assign _0340_ = _0721_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14412" *) IntSaturation_33U_32U_slc_IntSaturation_33U_32U_o_31_1_2_29_22_itm_3 : else_AluOp_data_slc_else_AluOp_data_1_30_23_21_itm_3;
  assign _0420_ = and_213_rgt ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) nor_37_cse : FpAdd_8U_23U_is_inf_2_lpi_1_dfm_2_mx0w0;
  assign _0110_ = _0720_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14403" *) _0420_ : FpAdd_8U_23U_is_inf_2_lpi_1_dfm_8;
  assign _0159_ = FpCmp_8U_23U_false_o_and_1_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14393" *) FpCmp_8U_23U_false_o_1_lpi_1_dfm_6_30_0_1 : FpCmp_8U_23U_false_o_1_lpi_1_dfm_7_30_0_1;
  assign _0161_ = FpCmp_8U_23U_false_o_and_1_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14393" *) FpCmp_8U_23U_false_o_2_lpi_1_dfm_7_30_0_1 : FpCmp_8U_23U_false_o_2_lpi_1_dfm_8_30_0_1;
  assign _0455_ = and_dcpl_127 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16600|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16599" *) IntSaturation_33U_32U_slc_IntSaturation_33U_32U_o_31_1_1_29_22_itm_2 : AluOut_data_2_30_23_lpi_1_dfm_3_mx1w0;
  assign _0074_ = _0717_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14383" *) _0455_ : AluOut_data_2_30_23_lpi_1_dfm_3;
  assign _0344_ = _0714_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14373" *) IntSaturation_33U_32U_slc_IntSaturation_33U_32U_o_31_1_3_29_22_itm_3 : else_AluOp_data_slc_else_AluOp_data_2_30_23_21_itm_3;
  assign _0419_ = and_211_rgt ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) nor_41_cse : FpAdd_8U_23U_is_inf_3_lpi_1_dfm_2_mx0w0;
  assign _0111_ = _0713_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14364" *) _0419_ : FpAdd_8U_23U_is_inf_3_lpi_1_dfm_8;
  assign _0163_ = _0710_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14355" *) FpCmp_8U_23U_false_o_3_lpi_1_dfm_7_30_0_1 : FpCmp_8U_23U_false_o_3_lpi_1_dfm_8_30_0_1;
  assign _0432_ = and_dcpl_127 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16464|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16463" *) IntSaturation_33U_32U_slc_IntSaturation_33U_32U_o_31_1_1_21_0_itm_2 : AluOut_data_2_22_1_lpi_1_dfm_3_mx1w0;
  assign _0073_ = _0709_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14346" *) _0432_ : AluOut_data_2_22_1_lpi_1_dfm_3;
  assign _0168_ = FpCmp_8U_23U_true_o_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14335" *) FpCmp_8U_23U_true_o_1_lpi_1_dfm_6_30_0_1 : FpCmp_8U_23U_true_o_1_lpi_1_dfm_7_30_0_1;
  assign _0171_ = FpCmp_8U_23U_true_o_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14335" *) FpCmp_8U_23U_true_o_2_lpi_1_dfm_6_30_0_1 : FpCmp_8U_23U_true_o_2_lpi_1_dfm_7_30_0_1;
  assign _0174_ = FpCmp_8U_23U_true_o_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14335" *) FpCmp_8U_23U_true_o_3_lpi_1_dfm_6_30_0_1 : FpCmp_8U_23U_true_o_3_lpi_1_dfm_7_30_0_1;
  assign _0142_ = FpAlu_8U_23U_and_82_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14321" *) FpAlu_8U_23U_equal_tmp_31 : FpAlu_8U_23U_equal_tmp_32;
  assign _0139_ = FpAlu_8U_23U_and_82_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14321" *) FpAlu_8U_23U_equal_tmp_28 : FpAlu_8U_23U_equal_tmp_29;
  assign _0150_ = FpAlu_8U_23U_and_82_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14321" *) FpAlu_8U_23U_nor_dfs_5 : FpAlu_8U_23U_nor_dfs_6;
  assign _0136_ = FpAlu_8U_23U_and_82_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14321" *) FpAlu_8U_23U_equal_tmp_25 : FpAlu_8U_23U_equal_tmp_26;
  assign _0133_ = FpAlu_8U_23U_and_82_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14321" *) FpAlu_8U_23U_equal_tmp_22 : FpAlu_8U_23U_equal_tmp_23;
  assign _0369_ = _0706_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14309" *) AluIn_data_mux1h_13_itm[22:0] : reg_AluIn_data_sva_4_30_0_1_itm;
  assign _0370_ = _0700_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14299" *) AluIn_data_mux1h_13_itm[30:23] : reg_AluIn_data_sva_4_30_0_itm;
  assign _0371_ = _0697_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14290" *) AluIn_data_mux1h_11_itm[22:0] : reg_AluIn_data_sva_4_62_32_1_itm;
  assign _0372_ = _0691_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14280" *) AluIn_data_mux1h_11_itm[30:23] : reg_AluIn_data_sva_4_62_32_itm;
  assign _0373_ = _0688_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14271" *) AluIn_data_mux1h_9_itm[22:0] : reg_AluIn_data_sva_4_94_64_1_itm;
  assign _0374_ = _0682_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14261" *) AluIn_data_mux1h_9_itm[30:23] : reg_AluIn_data_sva_4_94_64_itm;
  assign _0418_ = and_dcpl_99 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) alu_loop_op_1_FpMantRNE_49U_24U_else_and_svs_st : alu_loop_op_1_FpMantRNE_49U_24U_else_and_tmp;
  assign _0417_ = and_dcpl_99 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) alu_loop_op_2_FpMantRNE_49U_24U_else_and_2_svs_st : alu_loop_op_2_FpMantRNE_49U_24U_else_and_2_tmp;
  assign _0416_ = and_dcpl_99 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) alu_loop_op_3_FpMantRNE_49U_24U_else_and_1_svs_st : alu_loop_op_3_FpMantRNE_49U_24U_else_and_1_tmp;
  assign _0415_ = and_dcpl_99 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) alu_loop_op_4_FpMantRNE_49U_24U_else_and_3_svs_st : alu_loop_op_4_FpMantRNE_49U_24U_else_and_3_tmp;
  assign _0292_ = FpMantRNE_49U_24U_else_and_4_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14245" *) _0415_ : alu_loop_op_4_FpMantRNE_49U_24U_else_and_3_svs_st_2;
  assign _0279_ = FpMantRNE_49U_24U_else_and_4_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14245" *) _0416_ : alu_loop_op_3_FpMantRNE_49U_24U_else_and_1_svs_st_2;
  assign _0265_ = FpMantRNE_49U_24U_else_and_4_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14245" *) _0417_ : alu_loop_op_2_FpMantRNE_49U_24U_else_and_2_svs_st_2;
  assign _0253_ = FpMantRNE_49U_24U_else_and_4_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14245" *) _0418_ : alu_loop_op_1_FpMantRNE_49U_24U_else_and_svs_st_2;
  assign _0087_ = IsNaN_8U_23U_1_aelse_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14223" *) _0679_ : FpAdd_8U_23U_and_3_tmp_3;
  assign _0088_ = IsNaN_8U_23U_1_aelse_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14223" *) _0678_ : FpAdd_8U_23U_and_tmp_2;
  assign _0085_ = IsNaN_8U_23U_1_aelse_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14223" *) _0677_ : FpAdd_8U_23U_and_1_tmp_3;
  assign _0086_ = IsNaN_8U_23U_1_aelse_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14223" *) _0676_ : FpAdd_8U_23U_and_2_tmp_3;
  assign _0208_ = IsNaN_8U_23U_1_aelse_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14223" *) IsNaN_8U_23U_1_land_lpi_1_dfm_8 : IsNaN_8U_23U_1_land_lpi_1_dfm_9;
  assign _0205_ = IsNaN_8U_23U_1_aelse_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14223" *) IsNaN_8U_23U_1_land_3_lpi_1_dfm_8 : IsNaN_8U_23U_1_land_3_lpi_1_dfm_9;
  assign _0202_ = IsNaN_8U_23U_1_aelse_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14223" *) IsNaN_8U_23U_1_land_2_lpi_1_dfm_8 : IsNaN_8U_23U_1_land_2_lpi_1_dfm_9;
  assign _0199_ = IsNaN_8U_23U_1_aelse_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14223" *) IsNaN_8U_23U_1_land_1_lpi_1_dfm_8 : IsNaN_8U_23U_1_land_1_lpi_1_dfm_9;
  assign _0239_ = IsNaN_8U_23U_aelse_and_8_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14205" *) IsNaN_8U_23U_land_lpi_1_dfm_10 : IsNaN_8U_23U_land_lpi_1_dfm_11;
  assign _0233_ = IsNaN_8U_23U_aelse_and_8_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14205" *) IsNaN_8U_23U_land_3_lpi_1_dfm_10 : IsNaN_8U_23U_land_3_lpi_1_dfm_11;
  assign _0227_ = IsNaN_8U_23U_aelse_and_8_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14205" *) IsNaN_8U_23U_land_2_lpi_1_dfm_10 : IsNaN_8U_23U_land_2_lpi_1_dfm_11;
  assign _0221_ = IsNaN_8U_23U_aelse_and_8_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14205" *) IsNaN_8U_23U_land_1_lpi_1_dfm_10 : IsNaN_8U_23U_land_1_lpi_1_dfm_11;
  assign _0367_ = _0675_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14194" *) AluIn_data_mux1h_7_itm[22:0] : reg_AluIn_data_sva_4_126_96_1_itm;
  assign _0368_ = _0669_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14184" *) AluIn_data_mux1h_7_itm[30:23] : reg_AluIn_data_sva_4_126_96_itm;
  assign _0414_ = and_dcpl_99 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) alu_loop_op_4_FpAdd_8U_23U_if_4_if_slc_FpAdd_8U_23U_if_4_if_acc_1_7_3_svs_st_2 : alu_loop_op_4_FpAdd_8U_23U_if_4_if_acc_6_nl[7];
  assign _0287_ = _0664_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14173" *) _0414_ : alu_loop_op_4_FpAdd_8U_23U_if_4_if_slc_FpAdd_8U_23U_if_4_if_acc_1_7_3_svs_st_3;
  assign _0413_ = and_dcpl_99 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) alu_loop_op_3_FpAdd_8U_23U_if_4_if_slc_FpAdd_8U_23U_if_4_if_acc_1_7_1_svs_st_2 : alu_loop_op_3_FpAdd_8U_23U_if_4_if_acc_2_nl[7];
  assign _0274_ = _0663_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14161" *) _0413_ : alu_loop_op_3_FpAdd_8U_23U_if_4_if_slc_FpAdd_8U_23U_if_4_if_acc_1_7_1_svs_st_3;
  assign _0412_ = and_dcpl_99 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) alu_loop_op_2_FpAdd_8U_23U_if_4_if_slc_FpAdd_8U_23U_if_4_if_acc_1_7_2_svs_st_2 : alu_loop_op_2_FpAdd_8U_23U_if_4_if_acc_4_nl[7];
  assign _0260_ = _0662_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14149" *) _0412_ : alu_loop_op_2_FpAdd_8U_23U_if_4_if_slc_FpAdd_8U_23U_if_4_if_acc_1_7_2_svs_st_3;
  assign _0411_ = and_dcpl_99 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) alu_loop_op_1_FpAdd_8U_23U_if_4_if_slc_FpAdd_8U_23U_if_4_if_acc_1_7_svs_st_2 : alu_loop_op_1_FpAdd_8U_23U_if_4_if_acc_1_nl[7];
  assign _0248_ = _0661_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14137" *) _0411_ : alu_loop_op_1_FpAdd_8U_23U_if_4_if_slc_FpAdd_8U_23U_if_4_if_acc_1_7_svs_st_3;
  assign _0116_ = _0660_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14127" *) FpAdd_8U_23U_o_expo_lpi_1_dfm_2_mx0w0 : FpAdd_8U_23U_o_expo_lpi_1_dfm_13;
  assign _0454_ = and_dcpl_108 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16600|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16599" *) IntSaturation_33U_32U_slc_IntSaturation_33U_32U_o_31_1_29_22_itm_3 : FpAdd_8U_23U_o_expo_3_lpi_1_dfm_2_mx0w0;
  assign _0115_ = _0659_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14118" *) _0454_ : FpAdd_8U_23U_o_expo_3_lpi_1_dfm_13;
  assign _0453_ = and_dcpl_108 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16600|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16599" *) IntSaturation_33U_32U_slc_IntSaturation_33U_32U_o_31_1_3_29_22_itm_3 : FpAdd_8U_23U_o_expo_2_lpi_1_dfm_2_mx0w0;
  assign _0114_ = _0658_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14108" *) _0453_ : FpAdd_8U_23U_o_expo_2_lpi_1_dfm_13;
  assign _0452_ = and_dcpl_108 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16600|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16599" *) IntSaturation_33U_32U_slc_IntSaturation_33U_32U_o_31_1_2_29_22_itm_3 : FpAdd_8U_23U_o_expo_1_lpi_1_dfm_2_mx0w0;
  assign _0113_ = _0657_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14098" *) _0452_ : FpAdd_8U_23U_o_expo_1_lpi_1_dfm_13;
  assign _0360_ = _0655_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14089" *) _1363_ : main_stage_v_4;
  assign _0060_ = and_550_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14074" *) AluIn_data_sva_128[30:0] : AluIn_data_sva_3_30_0_1;
  assign _0061_ = and_550_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14074" *) AluIn_data_sva_128[62:32] : AluIn_data_sva_3_62_32_1;
  assign _0062_ = and_550_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14074" *) AluIn_data_sva_128[94:64] : AluIn_data_sva_3_94_64_1;
  assign _0059_ = and_550_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14074" *) AluIn_data_sva_128[126:96] : AluIn_data_sva_3_126_96_1;
  assign _0295_ = and_550_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14074" *) alu_loop_op_unequal_tmp_6 : alu_loop_op_unequal_tmp_7;
  assign _0355_ = and_550_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14074" *) io_read_cfg_alu_bypass_rsc_svs_st_5 : io_read_cfg_alu_bypass_rsc_svs_st_6;
  assign _0351_ = and_550_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14074" *) io_read_cfg_alu_bypass_rsc_svs_6 : io_read_cfg_alu_bypass_rsc_svs_7;
  assign _0302_ = _0653_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14060" *) cfg_alu_algo_1_sva_st_23 : cfg_alu_algo_1_sva_st_24;
  assign _0410_ = and_dcpl_99 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) FpNormalize_8U_49U_if_or_3_itm : FpNormalize_8U_49U_if_or_3_itm_mx0w0;
  assign _0183_ = _0652_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14051" *) _0410_ : FpNormalize_8U_49U_if_or_3_itm_2;
  assign _0409_ = and_dcpl_99 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) FpNormalize_8U_49U_if_or_2_itm : FpNormalize_8U_49U_if_or_2_itm_mx0w0;
  assign _0181_ = _0651_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14041" *) _0409_ : FpNormalize_8U_49U_if_or_2_itm_2;
  assign _0408_ = and_dcpl_99 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) FpNormalize_8U_49U_if_or_1_itm : FpNormalize_8U_49U_if_or_1_itm_mx0w0;
  assign _0179_ = _0650_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14031" *) _0408_ : FpNormalize_8U_49U_if_or_1_itm_2;
  assign _0407_ = and_dcpl_99 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) FpNormalize_8U_49U_if_or_itm : FpNormalize_8U_49U_if_or_itm_mx0w0;
  assign _0185_ = _0649_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:14021" *) _0407_ : FpNormalize_8U_49U_if_or_itm_2;
  assign _0406_ = and_dcpl_99 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) alu_loop_op_1_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_itm : acc_12_nl[50];
  assign _0405_ = and_dcpl_99 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) alu_loop_op_2_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_2_itm : acc_13_nl[50];
  assign _0404_ = and_dcpl_99 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) alu_loop_op_3_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_1_itm : acc_14_nl[50];
  assign _0403_ = and_dcpl_99 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) alu_loop_op_4_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_3_itm : acc_15_nl[50];
  assign _0443_ = FpAdd_8U_23U_int_mant_p1_or_3_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16566|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16565" *) FpAdd_8U_23U_int_mant_p1_lpi_1_dfm : acc_15_nl[50:1];
  assign _0442_ = FpAdd_8U_23U_int_mant_p1_or_3_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16566|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16565" *) FpAdd_8U_23U_int_mant_p1_3_lpi_1_dfm : acc_14_nl[50:1];
  assign _0441_ = FpAdd_8U_23U_int_mant_p1_or_3_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16566|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16565" *) FpAdd_8U_23U_int_mant_p1_2_lpi_1_dfm : acc_13_nl[50:1];
  assign _0440_ = FpAdd_8U_23U_int_mant_p1_or_3_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16566|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16565" *) FpAdd_8U_23U_int_mant_p1_1_lpi_1_dfm : acc_12_nl[50:1];
  assign _0290_ = FpAdd_8U_23U_int_mant_p1_and_4_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13997" *) _0403_ : alu_loop_op_4_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_3_itm_2;
  assign _0277_ = FpAdd_8U_23U_int_mant_p1_and_4_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13997" *) _0404_ : alu_loop_op_3_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_1_itm_2;
  assign _0263_ = FpAdd_8U_23U_int_mant_p1_and_4_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13997" *) _0405_ : alu_loop_op_2_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_2_itm_2;
  assign _0251_ = FpAdd_8U_23U_int_mant_p1_and_4_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13997" *) _0406_ : alu_loop_op_1_FpAdd_8U_23U_slc_FpAdd_8U_23U_int_mant_p1_49_itm_2;
  assign _0104_ = FpAdd_8U_23U_int_mant_p1_and_4_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13997" *) _0443_ : FpAdd_8U_23U_int_mant_p1_lpi_1_dfm_5;
  assign _0102_ = FpAdd_8U_23U_int_mant_p1_and_4_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13997" *) _0442_ : FpAdd_8U_23U_int_mant_p1_3_lpi_1_dfm_5;
  assign _0100_ = FpAdd_8U_23U_int_mant_p1_and_4_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13997" *) _0441_ : FpAdd_8U_23U_int_mant_p1_2_lpi_1_dfm_5;
  assign _0098_ = FpAdd_8U_23U_int_mant_p1_and_4_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13997" *) _0440_ : FpAdd_8U_23U_int_mant_p1_1_lpi_1_dfm_5;
  assign _0128_ = FpAdd_8U_23U_and_39_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13975" *) FpAdd_8U_23U_qr_lpi_1_dfm_6 : FpAdd_8U_23U_qr_lpi_1_dfm_7;
  assign _0125_ = FpAdd_8U_23U_and_39_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13975" *) FpAdd_8U_23U_qr_4_lpi_1_dfm_6 : FpAdd_8U_23U_qr_4_lpi_1_dfm_7;
  assign _0122_ = FpAdd_8U_23U_and_39_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13975" *) FpAdd_8U_23U_qr_3_lpi_1_dfm_6 : FpAdd_8U_23U_qr_3_lpi_1_dfm_7;
  assign _0119_ = FpAdd_8U_23U_and_39_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13975" *) FpAdd_8U_23U_qr_2_lpi_1_dfm_6 : FpAdd_8U_23U_qr_2_lpi_1_dfm_7;
  assign _0243_ = FpAdd_8U_23U_and_39_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13975" *) IsNaN_8U_23U_land_lpi_1_dfm_st_4 : IsNaN_8U_23U_land_lpi_1_dfm_st_5;
  assign _0237_ = FpAdd_8U_23U_and_39_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13975" *) IsNaN_8U_23U_land_3_lpi_1_dfm_st_4 : IsNaN_8U_23U_land_3_lpi_1_dfm_st_5;
  assign _0231_ = FpAdd_8U_23U_and_39_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13975" *) IsNaN_8U_23U_land_2_lpi_1_dfm_st_4 : IsNaN_8U_23U_land_2_lpi_1_dfm_st_5;
  assign _0225_ = FpAdd_8U_23U_and_39_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13975" *) IsNaN_8U_23U_land_1_lpi_1_dfm_st_4 : IsNaN_8U_23U_land_1_lpi_1_dfm_st_5;
  assign _0359_ = _0648_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13960" *) _1362_ : main_stage_v_3;
  assign _0350_ = AluIn_data_and_1_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13945" *) io_read_cfg_alu_bypass_rsc_svs_5 : io_read_cfg_alu_bypass_rsc_svs_6;
  assign _0058_ = AluIn_data_and_1_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13945" *) AluIn_data_sva_127 : AluIn_data_sva_128;
  assign _0294_ = AluIn_data_and_1_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13945" *) _1361_ : alu_loop_op_unequal_tmp_6;
  assign _0354_ = AluIn_data_and_1_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13945" *) io_read_cfg_alu_bypass_rsc_svs_st_1 : io_read_cfg_alu_bypass_rsc_svs_st_5;
  assign _0197_ = AluIn_data_and_1_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13945" *) IsNaN_8U_23U_1_land_1_lpi_1_dfm_mx0w0 : IsNaN_8U_23U_1_land_1_lpi_1_dfm_7;
  assign _0200_ = AluIn_data_and_1_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13945" *) IsNaN_8U_23U_1_land_2_lpi_1_dfm_mx0w0 : IsNaN_8U_23U_1_land_2_lpi_1_dfm_7;
  assign _0203_ = AluIn_data_and_1_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13945" *) IsNaN_8U_23U_1_land_3_lpi_1_dfm_mx0w0 : IsNaN_8U_23U_1_land_3_lpi_1_dfm_7;
  assign _0206_ = AluIn_data_and_1_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13945" *) IsNaN_8U_23U_1_land_lpi_1_dfm_mx0w0 : IsNaN_8U_23U_1_land_lpi_1_dfm_7;
  assign _0438_ = _1877_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16515|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16514" *) chn_alu_op_rsci_d_mxwt[126:96] : cfg_alu_op_1_sva_1[30:0];
  assign _0332_ = else_AluOp_data_and_10_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13925" *) _0438_ : else_AluOp_data_3_lpi_1_dfm_2_30_0_1;
  assign _0330_ = else_AluOp_data_and_10_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13925" *) else_AluOp_data_1_lpi_1_dfm_mx0[30:0] : else_AluOp_data_1_lpi_1_dfm_2_30_0_1;
  assign _0331_ = else_AluOp_data_and_10_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13925" *) else_AluOp_data_2_lpi_1_dfm_mx0[30:0] : else_AluOp_data_2_lpi_1_dfm_2_30_0_1;
  assign _0329_ = else_AluOp_data_and_10_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13925" *) else_AluOp_data_0_lpi_1_dfm_mx0[30:0] : else_AluOp_data_0_lpi_1_dfm_2_30_0_1;
  assign _0301_ = else_AluOp_data_and_10_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13925" *) cfg_alu_algo_1_sva_st_22 : cfg_alu_algo_1_sva_st_23;
  assign _0451_ = and_dcpl_99 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16600|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16599" *) FpAdd_8U_23U_a_right_shift_qr_1_lpi_1_dfm : FpAdd_8U_23U_a_right_shift_qr_1_lpi_1_dfm_mx0w0;
  assign _0450_ = and_dcpl_99 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16600|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16599" *) FpAdd_8U_23U_b_right_shift_qr_1_lpi_1_dfm : FpAdd_8U_23U_b_right_shift_qr_1_lpi_1_dfm_mx0w0;
  assign _0402_ = and_dcpl_99 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) alu_loop_op_1_FpAdd_8U_23U_IsZero_8U_23U_1_or_itm : alu_loop_op_1_FpAdd_8U_23U_IsZero_8U_23U_1_or_itm_mx0w0;
  assign _0401_ = and_dcpl_99 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) alu_loop_op_1_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_st : alu_loop_op_1_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_mx0w0;
  assign _0449_ = and_dcpl_99 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16600|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16599" *) FpAdd_8U_23U_a_right_shift_qr_2_lpi_1_dfm : FpAdd_8U_23U_a_right_shift_qr_2_lpi_1_dfm_mx0w0;
  assign _0448_ = and_dcpl_99 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16600|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16599" *) FpAdd_8U_23U_b_right_shift_qr_2_lpi_1_dfm : FpAdd_8U_23U_b_right_shift_qr_2_lpi_1_dfm_mx0w0;
  assign _0400_ = and_dcpl_99 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) alu_loop_op_2_FpAdd_8U_23U_IsZero_8U_23U_1_or_itm : alu_loop_op_2_FpAdd_8U_23U_IsZero_8U_23U_1_or_itm_mx0w0;
  assign _0399_ = and_dcpl_99 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) alu_loop_op_2_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_2_svs_st : alu_loop_op_2_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_2_svs_mx0w0;
  assign _0447_ = and_dcpl_99 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16600|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16599" *) FpAdd_8U_23U_a_right_shift_qr_3_lpi_1_dfm : FpAdd_8U_23U_a_right_shift_qr_3_lpi_1_dfm_mx0w0;
  assign _0446_ = and_dcpl_99 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16600|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16599" *) FpAdd_8U_23U_b_right_shift_qr_3_lpi_1_dfm : FpAdd_8U_23U_b_right_shift_qr_3_lpi_1_dfm_mx0w0;
  assign _0398_ = and_dcpl_99 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) alu_loop_op_3_FpAdd_8U_23U_IsZero_8U_23U_1_or_itm : alu_loop_op_3_FpAdd_8U_23U_IsZero_8U_23U_1_or_itm_mx0w0;
  assign _0397_ = and_dcpl_99 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) alu_loop_op_3_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_1_svs_st : alu_loop_op_3_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_1_svs_mx0w0;
  assign _0445_ = and_dcpl_99 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16600|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16599" *) FpAdd_8U_23U_a_right_shift_qr_lpi_1_dfm : FpAdd_8U_23U_a_right_shift_qr_lpi_1_dfm_mx0w0;
  assign _0444_ = and_dcpl_99 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16600|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16599" *) FpAdd_8U_23U_b_right_shift_qr_lpi_1_dfm : FpAdd_8U_23U_b_right_shift_qr_lpi_1_dfm_mx0w0;
  assign _0396_ = and_dcpl_99 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) alu_loop_op_4_FpAdd_8U_23U_IsZero_8U_23U_1_or_itm : alu_loop_op_4_FpAdd_8U_23U_IsZero_8U_23U_1_or_itm_mx0w0;
  assign _0395_ = and_dcpl_99 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) alu_loop_op_4_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_3_svs_st : alu_loop_op_4_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_3_svs_mx0w0;
  assign _0375_ = FpAdd_8U_23U_is_addition_and_8_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13874" *) _0401_ : reg_alu_loop_op_1_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_1_cse;
  assign _0376_ = FpAdd_8U_23U_is_addition_and_8_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13874" *) _0399_ : reg_alu_loop_op_2_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_2_svs_1_cse;
  assign _0377_ = FpAdd_8U_23U_is_addition_and_8_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13874" *) _0397_ : reg_alu_loop_op_3_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_1_svs_1_cse;
  assign _0378_ = FpAdd_8U_23U_is_addition_and_8_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13874" *) _0395_ : reg_alu_loop_op_4_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_3_svs_1_cse;
  assign _0282_ = FpAdd_8U_23U_is_addition_and_8_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13874" *) _0396_ : alu_loop_op_4_FpAdd_8U_23U_IsZero_8U_23U_1_or_itm_2;
  assign _0269_ = FpAdd_8U_23U_is_addition_and_8_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13874" *) _0398_ : alu_loop_op_3_FpAdd_8U_23U_IsZero_8U_23U_1_or_itm_2;
  assign _0256_ = FpAdd_8U_23U_is_addition_and_8_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13874" *) _0400_ : alu_loop_op_2_FpAdd_8U_23U_IsZero_8U_23U_1_or_itm_2;
  assign _0245_ = FpAdd_8U_23U_is_addition_and_8_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13874" *) _0402_ : alu_loop_op_1_FpAdd_8U_23U_IsZero_8U_23U_1_or_itm_2;
  assign _0096_ = FpAdd_8U_23U_is_addition_and_8_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13874" *) _0444_ : FpAdd_8U_23U_b_right_shift_qr_lpi_1_dfm_5;
  assign _0084_ = FpAdd_8U_23U_is_addition_and_8_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13874" *) _0445_ : FpAdd_8U_23U_a_right_shift_qr_lpi_1_dfm_5;
  assign _0094_ = FpAdd_8U_23U_is_addition_and_8_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13874" *) _0446_ : FpAdd_8U_23U_b_right_shift_qr_3_lpi_1_dfm_5;
  assign _0082_ = FpAdd_8U_23U_is_addition_and_8_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13874" *) _0447_ : FpAdd_8U_23U_a_right_shift_qr_3_lpi_1_dfm_5;
  assign _0092_ = FpAdd_8U_23U_is_addition_and_8_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13874" *) _0448_ : FpAdd_8U_23U_b_right_shift_qr_2_lpi_1_dfm_5;
  assign _0080_ = FpAdd_8U_23U_is_addition_and_8_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13874" *) _0449_ : FpAdd_8U_23U_a_right_shift_qr_2_lpi_1_dfm_5;
  assign _0090_ = FpAdd_8U_23U_is_addition_and_8_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13874" *) _0450_ : FpAdd_8U_23U_b_right_shift_qr_1_lpi_1_dfm_5;
  assign _0078_ = FpAdd_8U_23U_is_addition_and_8_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13874" *) _0451_ : FpAdd_8U_23U_a_right_shift_qr_1_lpi_1_dfm_5;
  assign _0246_ = IsNaN_8U_23U_aelse_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13836" *) IsNaN_8U_23U_4_nor_2_itm_2 : alu_loop_op_1_FpAdd_8U_23U_IsZero_8U_23U_or_itm_3;
  assign _0108_ = IsNaN_8U_23U_aelse_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13836" *) FpAdd_8U_23U_is_a_greater_lor_lpi_1_dfm_1_mx0w0 : FpAdd_8U_23U_is_a_greater_lor_lpi_1_dfm_6;
  assign _0107_ = IsNaN_8U_23U_aelse_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13836" *) FpAdd_8U_23U_is_a_greater_lor_3_lpi_1_dfm_1_mx0w0 : FpAdd_8U_23U_is_a_greater_lor_3_lpi_1_dfm_6;
  assign _0105_ = IsNaN_8U_23U_aelse_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13836" *) FpAdd_8U_23U_is_a_greater_lor_1_lpi_1_dfm_1_mx0w0 : FpAdd_8U_23U_is_a_greater_lor_1_lpi_1_dfm_6;
  assign _0106_ = IsNaN_8U_23U_aelse_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13836" *) FpAdd_8U_23U_is_a_greater_lor_2_lpi_1_dfm_1_mx0w0 : FpAdd_8U_23U_is_a_greater_lor_2_lpi_1_dfm_6;
  assign _0236_ = IsNaN_8U_23U_aelse_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13836" *) IsNaN_8U_23U_2_IsNaN_8U_23U_2_nor_3_itm_2 : IsNaN_8U_23U_land_3_lpi_1_dfm_st_4;
  assign _0230_ = IsNaN_8U_23U_aelse_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13836" *) IsNaN_8U_23U_2_IsNaN_8U_23U_2_nor_2_itm_1 : IsNaN_8U_23U_land_2_lpi_1_dfm_st_4;
  assign _0224_ = IsNaN_8U_23U_aelse_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13836" *) IsNaN_8U_23U_2_IsNaN_8U_23U_2_nor_1_itm_1 : IsNaN_8U_23U_land_1_lpi_1_dfm_st_4;
  assign _0285_ = IsNaN_8U_23U_aelse_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13836" *) alu_loop_op_4_FpAdd_8U_23U_IsZero_8U_23U_or_itm_4 : alu_loop_op_4_FpAdd_8U_23U_IsZero_8U_23U_or_itm_5;
  assign _0272_ = IsNaN_8U_23U_aelse_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13836" *) alu_loop_op_3_FpAdd_8U_23U_IsZero_8U_23U_or_itm_4 : alu_loop_op_3_FpAdd_8U_23U_IsZero_8U_23U_or_itm_5;
  assign _0258_ = IsNaN_8U_23U_aelse_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13836" *) IsNaN_8U_23U_4_nor_3_itm_3 : alu_loop_op_2_FpAdd_8U_23U_IsZero_8U_23U_or_itm_4;
  assign _0242_ = IsNaN_8U_23U_aelse_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13836" *) IsNaN_8U_23U_2_IsNaN_8U_23U_2_nor_itm_2 : IsNaN_8U_23U_land_lpi_1_dfm_st_4;
  assign _0358_ = _0647_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13817" *) _1360_ : main_stage_v_2;
  assign _0353_ = _0646_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13809" *) cfg_alu_bypass_rsci_d : io_read_cfg_alu_bypass_rsc_svs_st_1;
  assign _0394_ = cfg_alu_src_1_sva_st_1_mx0c1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) cfg_alu_src_1_sva_st : cfg_alu_src_rsci_d;
  assign _0307_ = _0645_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13799" *) _0394_ : cfg_alu_src_1_sva_st_1;
  assign _0439_ = and_167_rgt ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16532|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16531" *) chn_alu_op_rsci_d_mxwt[127:96] : cfg_alu_op_rsci_d;
  assign _0305_ = _0643_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13788" *) _0439_ : cfg_alu_op_1_sva_1;
  assign _0437_ = and_dcpl_81 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16498|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16497" *) cfg_alu_algo_1_sva_st : cfg_alu_algo_rsci_d;
  assign _0300_ = _0641_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13779" *) _0437_ : cfg_alu_algo_1_sva_st_22;
  assign _0387_ = _0640_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13771" *) cfg_alu_algo_cfg_alu_algo_mux_3_itm : reg_cfg_alu_algo_1_sva_st_13_cse;
  assign _0304_ = _0639_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13763" *) cfg_alu_algo_cfg_alu_algo_mux_3_itm : cfg_alu_algo_1_sva_st_28;
  assign _0349_ = AluIn_data_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13750" *) cfg_alu_bypass_rsci_d : io_read_cfg_alu_bypass_rsc_svs_5;
  assign _0057_ = AluIn_data_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13750" *) chn_alu_in_rsci_d_mxwt : AluIn_data_sva_127;
  assign _0222_ = AluIn_data_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13750" *) IsNaN_8U_23U_2_IsNaN_8U_23U_2_nor_itm_mx0w0 : IsNaN_8U_23U_land_1_lpi_1_dfm_8;
  assign _0228_ = AluIn_data_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13750" *) IsNaN_8U_23U_2_IsNaN_8U_23U_2_nor_1_itm_mx0w0 : IsNaN_8U_23U_land_2_lpi_1_dfm_8;
  assign _0234_ = AluIn_data_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13750" *) IsNaN_8U_23U_2_IsNaN_8U_23U_2_nor_2_itm_mx0w0 : IsNaN_8U_23U_land_3_lpi_1_dfm_8;
  assign _0240_ = AluIn_data_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13750" *) IsNaN_8U_23U_2_IsNaN_8U_23U_2_nor_3_itm_mx0w0 : IsNaN_8U_23U_land_lpi_1_dfm_8;
  assign _0357_ = _0638_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13737" *) _1355_ : main_stage_v_1;
  assign _0311_ = _0637_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13729" *) _1354_ : chn_alu_op_rsci_ld_core_psct;
  assign _0389_ = _0633_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13720" *) _1353_ : reg_chn_alu_out_rsci_ld_core_psct_cse;
  assign _0324_ = chn_alu_out_and_18_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13711" *) AluOut_data_2_22_1_lpi_1_dfm_3_mx1w0 : chn_alu_out_rsci_d_86_65;
  assign _0325_ = chn_alu_out_and_18_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13711" *) AluOut_data_2_30_23_lpi_1_dfm_3_mx1w0 : chn_alu_out_rsci_d_94_87;
  assign _0393_ = and_dcpl_40 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) alu_loop_op_mux_204_mx1w1 : reg_AluIn_data_sva_4_94_64_1_itm[0];
  assign _0323_ = _0632_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13701" *) _0393_ : chn_alu_out_rsci_d_64;
  assign _0317_ = chn_alu_out_and_1_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13680" *) _2405_ : chn_alu_out_rsci_d_30_23;
  assign _0318_ = chn_alu_out_and_1_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13680" *) mux_177_itm_4 : chn_alu_out_rsci_d_31;
  assign _0321_ = chn_alu_out_and_1_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13680" *) _2406_ : chn_alu_out_rsci_d_62_55;
  assign _0322_ = chn_alu_out_and_1_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13680" *) mux_181_itm_4 : chn_alu_out_rsci_d_63;
  assign _0326_ = chn_alu_out_and_1_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13680" *) AluOut_data_2_31_lpi_1_dfm_7 : chn_alu_out_rsci_d_95;
  assign _0313_ = chn_alu_out_and_1_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13680" *) _2382_ : chn_alu_out_rsci_d_118_97;
  assign _0314_ = chn_alu_out_and_1_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13680" *) _2407_ : chn_alu_out_rsci_d_126_119;
  assign _0315_ = chn_alu_out_and_1_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13680" *) mux_189_itm_4 : chn_alu_out_rsci_d_127;
  assign _0320_ = and_734_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13662" *) _2381_ : chn_alu_out_rsci_d_54_33;
  assign _0316_ = and_734_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13662" *) _2380_ : chn_alu_out_rsci_d_22_1;
  assign _0392_ = and_dcpl_40 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) alu_loop_op_mux_212_nl : reg_AluIn_data_sva_4_126_96_1_itm[0];
  assign _0391_ = and_dcpl_40 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) alu_loop_op_mux_210_nl : reg_AluIn_data_sva_4_62_32_1_itm[0];
  assign _0390_ = and_dcpl_40 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16447|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:16446" *) alu_loop_op_mux_209_nl : reg_AluIn_data_sva_4_30_0_1_itm[0];
  assign _0319_ = chn_alu_out_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13648" *) _0391_ : chn_alu_out_rsci_d_32;
  assign _0327_ = chn_alu_out_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13648" *) _0392_ : chn_alu_out_rsci_d_96;
  assign _0312_ = chn_alu_out_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13648" *) _0390_ : chn_alu_out_rsci_d_0;
  assign _0309_ = _0631_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13638" *) chn_alu_in_rsci_ld_core_psct_mx0c0 : chn_alu_in_rsci_ld_core_psct;
  assign _0388_ = core_wen ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13627" *) or_tmp_695 : reg_cfg_alu_algo_rsc_triosy_obj_ld_core_psct_cse;
  assign _0308_ = core_wen ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13627" *) _1352_ : chn_alu_in_rsci_iswt0;
  assign _0310_ = core_wen ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13627" *) and_357_cse : chn_alu_op_rsci_iswt0;
  assign _0328_ = core_wen ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:13627" *) and_dcpl_43 : chn_alu_out_rsci_iswt0;
  assign _2435_ = AluIn_data_sva_127[127] ^ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12657" *) else_AluOp_data_3_lpi_1_dfm_mx0[31];
  assign _2436_ = AluIn_data_sva_127[95] ^ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12667" *) else_AluOp_data_2_lpi_1_dfm_mx0[31];
  assign _2437_ = AluIn_data_sva_127[63] ^ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12678" *) else_AluOp_data_1_lpi_1_dfm_mx0[31];
  assign _2438_ = AluIn_data_sva_127[31] ^ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12689" *) else_AluOp_data_0_lpi_1_dfm_mx0[31];
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12227" *)
  SDP_Y_CORE_Y_alu_core_cfg_alu_algo_rsc_triosy_obj Y_alu_core_cfg_alu_algo_rsc_triosy_obj_inst (
    .cfg_alu_algo_rsc_triosy_lz(cfg_alu_algo_rsc_triosy_lz),
    .cfg_alu_algo_rsc_triosy_obj_bawt(cfg_alu_algo_rsc_triosy_obj_bawt),
    .cfg_alu_algo_rsc_triosy_obj_iswt0(reg_cfg_alu_algo_rsc_triosy_obj_ld_core_psct_cse),
    .cfg_alu_algo_rsc_triosy_obj_oswt(cfg_alu_algo_rsc_triosy_obj_oswt),
    .core_wen(core_wen),
    .core_wten(core_wten),
    .nvdla_core_clk(nvdla_core_clk),
    .nvdla_core_rstn(nvdla_core_rstn)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12194" *)
  SDP_Y_CORE_Y_alu_core_cfg_alu_bypass_rsc_triosy_obj Y_alu_core_cfg_alu_bypass_rsc_triosy_obj_inst (
    .cfg_alu_bypass_rsc_triosy_lz(cfg_alu_bypass_rsc_triosy_lz),
    .cfg_alu_bypass_rsc_triosy_obj_bawt(cfg_alu_bypass_rsc_triosy_obj_bawt),
    .cfg_alu_bypass_rsc_triosy_obj_iswt0(reg_cfg_alu_algo_rsc_triosy_obj_ld_core_psct_cse),
    .cfg_alu_bypass_rsc_triosy_obj_oswt(cfg_alu_bypass_rsc_triosy_obj_oswt),
    .core_wen(core_wen),
    .core_wten(core_wten),
    .nvdla_core_clk(nvdla_core_clk),
    .nvdla_core_rstn(nvdla_core_rstn)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12216" *)
  SDP_Y_CORE_Y_alu_core_cfg_alu_op_rsc_triosy_obj Y_alu_core_cfg_alu_op_rsc_triosy_obj_inst (
    .cfg_alu_op_rsc_triosy_lz(cfg_alu_op_rsc_triosy_lz),
    .cfg_alu_op_rsc_triosy_obj_bawt(cfg_alu_op_rsc_triosy_obj_bawt),
    .cfg_alu_op_rsc_triosy_obj_iswt0(reg_cfg_alu_algo_rsc_triosy_obj_ld_core_psct_cse),
    .cfg_alu_op_rsc_triosy_obj_oswt(cfg_alu_op_rsc_triosy_obj_oswt),
    .core_wen(core_wen),
    .core_wten(core_wten),
    .nvdla_core_clk(nvdla_core_clk),
    .nvdla_core_rstn(nvdla_core_rstn)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12205" *)
  SDP_Y_CORE_Y_alu_core_cfg_alu_src_rsc_triosy_obj Y_alu_core_cfg_alu_src_rsc_triosy_obj_inst (
    .cfg_alu_src_rsc_triosy_lz(cfg_alu_src_rsc_triosy_lz),
    .cfg_alu_src_rsc_triosy_obj_bawt(cfg_alu_src_rsc_triosy_obj_bawt),
    .cfg_alu_src_rsc_triosy_obj_iswt0(reg_cfg_alu_algo_rsc_triosy_obj_ld_core_psct_cse),
    .cfg_alu_src_rsc_triosy_obj_oswt(cfg_alu_src_rsc_triosy_obj_oswt),
    .core_wen(core_wen),
    .core_wten(core_wten),
    .nvdla_core_clk(nvdla_core_clk),
    .nvdla_core_rstn(nvdla_core_rstn)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12149" *)
  SDP_Y_CORE_Y_alu_core_chn_alu_in_rsci Y_alu_core_chn_alu_in_rsci_inst (
    .chn_alu_in_rsc_lz(chn_alu_in_rsc_lz),
    .chn_alu_in_rsc_vz(chn_alu_in_rsc_vz),
    .chn_alu_in_rsc_z(chn_alu_in_rsc_z),
    .chn_alu_in_rsci_bawt(chn_alu_in_rsci_bawt),
    .chn_alu_in_rsci_d_mxwt(chn_alu_in_rsci_d_mxwt),
    .chn_alu_in_rsci_iswt0(chn_alu_in_rsci_iswt0),
    .chn_alu_in_rsci_ld_core_psct(chn_alu_in_rsci_ld_core_psct),
    .chn_alu_in_rsci_oswt(chn_alu_in_rsci_oswt),
    .chn_alu_in_rsci_wen_comp(chn_alu_in_rsci_wen_comp),
    .core_wen(core_wen),
    .core_wten(core_wten),
    .nvdla_core_clk(nvdla_core_clk),
    .nvdla_core_rstn(nvdla_core_rstn)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12164" *)
  SDP_Y_CORE_Y_alu_core_chn_alu_op_rsci Y_alu_core_chn_alu_op_rsci_inst (
    .chn_alu_op_rsc_lz(chn_alu_op_rsc_lz),
    .chn_alu_op_rsc_vz(chn_alu_op_rsc_vz),
    .chn_alu_op_rsc_z(chn_alu_op_rsc_z),
    .chn_alu_op_rsci_bawt(chn_alu_op_rsci_bawt),
    .chn_alu_op_rsci_d_mxwt(chn_alu_op_rsci_d_mxwt),
    .chn_alu_op_rsci_iswt0(chn_alu_op_rsci_iswt0),
    .chn_alu_op_rsci_ld_core_psct(chn_alu_op_rsci_ld_core_psct),
    .chn_alu_op_rsci_oswt(chn_alu_op_rsci_oswt),
    .chn_alu_op_rsci_wen_comp(chn_alu_op_rsci_wen_comp),
    .core_wen(core_wen),
    .core_wten(core_wten),
    .nvdla_core_clk(nvdla_core_clk),
    .nvdla_core_rstn(nvdla_core_rstn)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12179" *)
  SDP_Y_CORE_Y_alu_core_chn_alu_out_rsci Y_alu_core_chn_alu_out_rsci_inst (
    .chn_alu_out_rsc_lz(chn_alu_out_rsc_lz),
    .chn_alu_out_rsc_vz(chn_alu_out_rsc_vz),
    .chn_alu_out_rsc_z(chn_alu_out_rsc_z),
    .chn_alu_out_rsci_bawt(chn_alu_out_rsci_bawt),
    .chn_alu_out_rsci_d({ chn_alu_out_rsci_d_127, chn_alu_out_rsci_d_126_119, chn_alu_out_rsci_d_118_97, chn_alu_out_rsci_d_96, chn_alu_out_rsci_d_95, chn_alu_out_rsci_d_94_87, chn_alu_out_rsci_d_86_65, chn_alu_out_rsci_d_64, chn_alu_out_rsci_d_63, chn_alu_out_rsci_d_62_55, chn_alu_out_rsci_d_54_33, chn_alu_out_rsci_d_32, chn_alu_out_rsci_d_31, chn_alu_out_rsci_d_30_23, chn_alu_out_rsci_d_22_1, chn_alu_out_rsci_d_0 }),
    .chn_alu_out_rsci_iswt0(chn_alu_out_rsci_iswt0),
    .chn_alu_out_rsci_ld_core_psct(reg_chn_alu_out_rsci_ld_core_psct_cse),
    .chn_alu_out_rsci_oswt(chn_alu_out_rsci_oswt),
    .chn_alu_out_rsci_wen_comp(chn_alu_out_rsci_wen_comp),
    .core_wen(core_wen),
    .core_wten(core_wten),
    .nvdla_core_clk(nvdla_core_clk),
    .nvdla_core_rstn(nvdla_core_rstn)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12247" *)
  SDP_Y_CORE_Y_alu_core_core_fsm Y_alu_core_core_fsm_inst (
    .core_wen(core_wen),
    .fsm_output(fsm_output),
    .nvdla_core_clk(nvdla_core_clk),
    .nvdla_core_rstn(nvdla_core_rstn)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12238" *)
  SDP_Y_CORE_Y_alu_core_staller Y_alu_core_staller_inst (
    .chn_alu_in_rsci_wen_comp(chn_alu_in_rsci_wen_comp),
    .chn_alu_op_rsci_wen_comp(chn_alu_op_rsci_wen_comp),
    .chn_alu_out_rsci_wen_comp(chn_alu_out_rsci_wen_comp),
    .core_wen(core_wen),
    .core_wten(core_wten),
    .nvdla_core_clk(nvdla_core_clk),
    .nvdla_core_rstn(nvdla_core_rstn)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12093" *)
  \$paramod\SDP_Y_CORE_mgc_shift_bl_v4\width_a=24\signd_a=0\width_s=9\width_z=49  alu_loop_op_1_FpAdd_8U_23U_a_int_mant_p1_lshift_rg (
    .a({ alu_loop_op_1_FpAdd_8U_23U_IsZero_8U_23U_or_itm_3, AluIn_data_sva_128[22:0] }),
    .s({ alu_loop_op_1_FpAdd_8U_23U_a_left_shift_acc_nl, nl_alu_loop_op_1_FpAdd_8U_23U_a_int_mant_p1_lshift_rg_s[0] }),
    .z(FpAdd_8U_23U_a_int_mant_p1_1_sva)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12037" *)
  \$paramod\SDP_Y_CORE_mgc_shift_bl_v4\width_a=24\signd_a=0\width_s=9\width_z=49  alu_loop_op_1_FpAdd_8U_23U_b_int_mant_p1_lshift_rg (
    .a({ alu_loop_op_1_FpAdd_8U_23U_IsZero_8U_23U_1_or_itm_2, else_AluOp_data_0_lpi_1_dfm_2_30_0_1[22:0] }),
    .s({ alu_loop_op_1_FpAdd_8U_23U_b_left_shift_acc_nl, nl_alu_loop_op_1_FpAdd_8U_23U_b_int_mant_p1_lshift_rg_s[0] }),
    .z(FpAdd_8U_23U_addend_larger_asn_19_mx0w1)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12141" *)
  \$paramod\SDP_Y_CORE_mgc_shift_l_v4\width_a=49\signd_a=0\width_s=6\width_z=49  alu_loop_op_1_FpNormalize_8U_49U_else_lshift_rg (
    .a(FpAdd_8U_23U_int_mant_p1_1_lpi_1_dfm_5[48:0]),
    .s(libraries_leading_sign_49_0_78e877fc94067377fcee479dbb0ed8e083a3_4),
    .z(alu_loop_op_1_FpNormalize_8U_49U_else_lshift_itm)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12101" *)
  SDP_Y_CORE_leading_sign_49_0 alu_loop_op_1_leading_sign_49_0_rg (
    .mantissa(FpAdd_8U_23U_int_mant_p1_1_lpi_1_dfm_5[48:0]),
    .rtn(libraries_leading_sign_49_0_78e877fc94067377fcee479dbb0ed8e083a3_4)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12085" *)
  \$paramod\SDP_Y_CORE_mgc_shift_bl_v4\width_a=24\signd_a=0\width_s=9\width_z=49  alu_loop_op_2_FpAdd_8U_23U_a_int_mant_p1_lshift_2_rg (
    .a({ alu_loop_op_2_FpAdd_8U_23U_IsZero_8U_23U_or_itm_4, AluIn_data_sva_128[54:32] }),
    .s({ alu_loop_op_2_FpAdd_8U_23U_a_left_shift_acc_2_nl, nl_alu_loop_op_2_FpAdd_8U_23U_a_int_mant_p1_lshift_2_rg_s[0] }),
    .z(FpAdd_8U_23U_a_int_mant_p1_2_sva)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12045" *)
  \$paramod\SDP_Y_CORE_mgc_shift_bl_v4\width_a=24\signd_a=0\width_s=9\width_z=49  alu_loop_op_2_FpAdd_8U_23U_b_int_mant_p1_lshift_2_rg (
    .a({ alu_loop_op_2_FpAdd_8U_23U_IsZero_8U_23U_1_or_itm_2, else_AluOp_data_1_lpi_1_dfm_2_30_0_1[22:0] }),
    .s({ alu_loop_op_2_FpAdd_8U_23U_b_left_shift_acc_2_nl, nl_alu_loop_op_2_FpAdd_8U_23U_b_int_mant_p1_lshift_2_rg_s[0] }),
    .z(FpAdd_8U_23U_addend_larger_asn_13_mx0w1)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12133" *)
  \$paramod\SDP_Y_CORE_mgc_shift_l_v4\width_a=49\signd_a=0\width_s=6\width_z=49  alu_loop_op_2_FpNormalize_8U_49U_else_lshift_2_rg (
    .a(FpAdd_8U_23U_int_mant_p1_2_lpi_1_dfm_5[48:0]),
    .s(libraries_leading_sign_49_0_78e877fc94067377fcee479dbb0ed8e083a3_5),
    .z(alu_loop_op_2_FpNormalize_8U_49U_else_lshift_2_itm)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12105" *)
  SDP_Y_CORE_leading_sign_49_0 alu_loop_op_2_leading_sign_49_0_2_rg (
    .mantissa(FpAdd_8U_23U_int_mant_p1_2_lpi_1_dfm_5[48:0]),
    .rtn(libraries_leading_sign_49_0_78e877fc94067377fcee479dbb0ed8e083a3_5)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12077" *)
  \$paramod\SDP_Y_CORE_mgc_shift_bl_v4\width_a=24\signd_a=0\width_s=9\width_z=49  alu_loop_op_3_FpAdd_8U_23U_a_int_mant_p1_lshift_1_rg (
    .a({ alu_loop_op_3_FpAdd_8U_23U_IsZero_8U_23U_or_itm_5, AluIn_data_sva_128[86:64] }),
    .s({ alu_loop_op_3_FpAdd_8U_23U_a_left_shift_acc_1_nl, nl_alu_loop_op_3_FpAdd_8U_23U_a_int_mant_p1_lshift_1_rg_s[0] }),
    .z(FpAdd_8U_23U_a_int_mant_p1_3_sva)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12053" *)
  \$paramod\SDP_Y_CORE_mgc_shift_bl_v4\width_a=24\signd_a=0\width_s=9\width_z=49  alu_loop_op_3_FpAdd_8U_23U_b_int_mant_p1_lshift_1_rg (
    .a({ alu_loop_op_3_FpAdd_8U_23U_IsZero_8U_23U_1_or_itm_2, else_AluOp_data_2_lpi_1_dfm_2_30_0_1[22:0] }),
    .s({ alu_loop_op_3_FpAdd_8U_23U_b_left_shift_acc_1_nl, nl_alu_loop_op_3_FpAdd_8U_23U_b_int_mant_p1_lshift_1_rg_s[0] }),
    .z(FpAdd_8U_23U_addend_larger_asn_7_mx0w1)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12125" *)
  \$paramod\SDP_Y_CORE_mgc_shift_l_v4\width_a=49\signd_a=0\width_s=6\width_z=49  alu_loop_op_3_FpNormalize_8U_49U_else_lshift_1_rg (
    .a(FpAdd_8U_23U_int_mant_p1_3_lpi_1_dfm_5[48:0]),
    .s(libraries_leading_sign_49_0_78e877fc94067377fcee479dbb0ed8e083a3_6),
    .z(alu_loop_op_3_FpNormalize_8U_49U_else_lshift_1_itm)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12109" *)
  SDP_Y_CORE_leading_sign_49_0 alu_loop_op_3_leading_sign_49_0_1_rg (
    .mantissa(FpAdd_8U_23U_int_mant_p1_3_lpi_1_dfm_5[48:0]),
    .rtn(libraries_leading_sign_49_0_78e877fc94067377fcee479dbb0ed8e083a3_6)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12069" *)
  \$paramod\SDP_Y_CORE_mgc_shift_bl_v4\width_a=24\signd_a=0\width_s=9\width_z=49  alu_loop_op_4_FpAdd_8U_23U_a_int_mant_p1_lshift_3_rg (
    .a({ alu_loop_op_4_FpAdd_8U_23U_IsZero_8U_23U_or_itm_5, AluIn_data_sva_128[118:96] }),
    .s({ alu_loop_op_4_FpAdd_8U_23U_a_left_shift_acc_3_nl, nl_alu_loop_op_4_FpAdd_8U_23U_a_int_mant_p1_lshift_3_rg_s[0] }),
    .z(FpAdd_8U_23U_a_int_mant_p1_sva)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12061" *)
  \$paramod\SDP_Y_CORE_mgc_shift_bl_v4\width_a=24\signd_a=0\width_s=9\width_z=49  alu_loop_op_4_FpAdd_8U_23U_b_int_mant_p1_lshift_3_rg (
    .a({ alu_loop_op_4_FpAdd_8U_23U_IsZero_8U_23U_1_or_itm_2, else_AluOp_data_3_lpi_1_dfm_2_30_0_1[22:0] }),
    .s({ alu_loop_op_4_FpAdd_8U_23U_b_left_shift_acc_3_nl, nl_alu_loop_op_4_FpAdd_8U_23U_b_int_mant_p1_lshift_3_rg_s[0] }),
    .z(FpAdd_8U_23U_addend_larger_asn_1_mx0w1)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12117" *)
  \$paramod\SDP_Y_CORE_mgc_shift_l_v4\width_a=49\signd_a=0\width_s=6\width_z=49  alu_loop_op_4_FpNormalize_8U_49U_else_lshift_3_rg (
    .a(FpAdd_8U_23U_int_mant_p1_lpi_1_dfm_5[48:0]),
    .s(libraries_leading_sign_49_0_78e877fc94067377fcee479dbb0ed8e083a3_7),
    .z(alu_loop_op_4_FpNormalize_8U_49U_else_lshift_3_itm)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:12113" *)
  SDP_Y_CORE_leading_sign_49_0 alu_loop_op_4_leading_sign_49_0_3_rg (
    .mantissa(FpAdd_8U_23U_int_mant_p1_lpi_1_dfm_5[48:0]),
    .rtn(libraries_leading_sign_49_0_78e877fc94067377fcee479dbb0ed8e083a3_7)
  );
  assign _0041_[1] = _0041_[2];
  assign _0042_[1] = _0042_[2];
  assign _0043_[1] = _0043_[2];
  assign _0044_[1] = _0044_[2];
  assign _0045_[7:0] = { _0045_[8], FpNormalize_8U_49U_else_mux_4_nl, 1'b1 };
  assign _0046_[7:0] = { _0046_[8], FpNormalize_8U_49U_else_mux_5_nl, 1'b1 };
  assign _0047_[7:0] = { _0047_[8], FpNormalize_8U_49U_else_mux_6_nl, 1'b1 };
  assign _0048_[7:0] = { _0048_[8], FpNormalize_8U_49U_else_mux_7_nl, 1'b1 };
  assign _1135_[6:0] = _1059_;
  assign FpAdd_8U_23U_is_a_greater_oif_aelse_acc_1_itm_23_1 = FpAdd_8U_23U_is_a_greater_oif_aelse_acc_1_nl[23];
  assign FpAdd_8U_23U_is_a_greater_oif_aelse_acc_2_itm_23_1 = FpAdd_8U_23U_is_a_greater_oif_aelse_acc_2_nl[23];
  assign FpAdd_8U_23U_is_a_greater_oif_aelse_acc_3_itm_23_1 = FpAdd_8U_23U_is_a_greater_oif_aelse_acc_3_nl[23];
  assign FpAdd_8U_23U_is_a_greater_oif_aelse_acc_itm_23_1 = FpAdd_8U_23U_is_a_greater_oif_aelse_acc_nl[23];
  assign FpCmp_8U_23U_false_else_if_acc_6_itm_8 = FpCmp_8U_23U_false_else_if_acc_6_nl[8];
  assign FpCmp_8U_23U_true_else_else_if_acc_4_itm_23 = FpCmp_8U_23U_true_else_else_if_acc_4_nl[23];
  assign FpCmp_8U_23U_true_if_acc_10_itm_8 = FpCmp_8U_23U_true_if_acc_10_nl[8];
  assign FpCmp_8U_23U_true_if_acc_4_itm_8 = FpCmp_8U_23U_true_if_acc_4_nl[8];
  assign FpCmp_8U_23U_true_if_acc_6_itm_8 = FpCmp_8U_23U_true_if_acc_6_nl[8];
  assign FpCmp_8U_23U_true_if_acc_8_itm_8 = FpCmp_8U_23U_true_if_acc_8_nl[8];
  assign alu_loop_op_1_FpAdd_8U_23U_if_3_if_acc_1_itm_7_1 = alu_loop_op_1_FpAdd_8U_23U_if_3_if_acc_1_nl[7];
  assign alu_loop_op_1_FpAdd_8U_23U_if_4_if_acc_1_itm_7_1 = alu_loop_op_1_FpAdd_8U_23U_if_4_if_acc_1_nl[7];
  assign alu_loop_op_1_IntSaturation_33U_32U_else_if_acc_itm_2_1 = alu_loop_op_1_IntSaturation_33U_32U_else_if_acc_nl[2];
  assign alu_loop_op_1_IntSaturation_33U_32U_if_acc_itm_2 = alu_loop_op_1_IntSaturation_33U_32U_if_acc_nl[2];
  assign alu_loop_op_2_FpAdd_8U_23U_if_3_if_acc_4_itm_7_1 = alu_loop_op_2_FpAdd_8U_23U_if_3_if_acc_4_nl[7];
  assign alu_loop_op_2_FpAdd_8U_23U_if_4_if_acc_4_itm_7_1 = alu_loop_op_2_FpAdd_8U_23U_if_4_if_acc_4_nl[7];
  assign alu_loop_op_2_IntSaturation_33U_32U_else_if_acc_1_itm_2_1 = alu_loop_op_2_IntSaturation_33U_32U_else_if_acc_1_nl[2];
  assign alu_loop_op_2_IntSaturation_33U_32U_if_acc_1_itm_2 = alu_loop_op_2_IntSaturation_33U_32U_if_acc_1_nl[2];
  assign alu_loop_op_3_FpAdd_8U_23U_if_3_if_acc_2_itm_7_1 = alu_loop_op_3_FpAdd_8U_23U_if_3_if_acc_2_nl[7];
  assign alu_loop_op_3_FpAdd_8U_23U_if_4_if_acc_2_itm_7_1 = alu_loop_op_3_FpAdd_8U_23U_if_4_if_acc_2_nl[7];
  assign alu_loop_op_3_IntSaturation_33U_32U_else_if_acc_itm_2_1 = alu_loop_op_3_IntSaturation_33U_32U_else_if_acc_nl[2];
  assign alu_loop_op_3_IntSaturation_33U_32U_if_acc_itm_2 = alu_loop_op_3_IntSaturation_33U_32U_if_acc_nl[2];
  assign alu_loop_op_4_FpAdd_8U_23U_if_3_if_acc_6_itm_7_1 = alu_loop_op_4_FpAdd_8U_23U_if_3_if_acc_6_nl[7];
  assign alu_loop_op_4_FpAdd_8U_23U_if_4_if_acc_6_itm_7_1 = alu_loop_op_4_FpAdd_8U_23U_if_4_if_acc_6_nl[7];
  assign alu_loop_op_4_IntSaturation_33U_32U_else_if_acc_1_itm_2_1 = alu_loop_op_4_IntSaturation_33U_32U_else_if_acc_1_nl[2];
  assign alu_loop_op_4_IntSaturation_33U_32U_if_acc_1_itm_2 = alu_loop_op_4_IntSaturation_33U_32U_if_acc_1_nl[2];
  assign and_729_nl = and_218_nl;
  assign cfg_alu_bypass_rsc_triosy_obj_oswt_unreg_pff = and_dcpl_64;
  assign chn_alu_in_rsci_oswt_unreg = or_tmp_695;
  assign nl_FpAdd_8U_23U_is_a_greater_oif_aelse_acc_1_nl[23:0] = FpAdd_8U_23U_is_a_greater_oif_aelse_acc_1_nl;
  assign nl_FpAdd_8U_23U_is_a_greater_oif_aelse_acc_2_nl[23:0] = FpAdd_8U_23U_is_a_greater_oif_aelse_acc_2_nl;
  assign nl_FpAdd_8U_23U_is_a_greater_oif_aelse_acc_3_nl[23:0] = FpAdd_8U_23U_is_a_greater_oif_aelse_acc_3_nl;
  assign nl_FpAdd_8U_23U_is_a_greater_oif_aelse_acc_nl[23:0] = FpAdd_8U_23U_is_a_greater_oif_aelse_acc_nl;
  assign nl_FpCmp_8U_23U_false_else_if_acc_10_nl[8:0] = FpCmp_8U_23U_false_else_if_acc_10_nl;
  assign nl_FpCmp_8U_23U_false_else_if_acc_4_nl[8:0] = FpCmp_8U_23U_false_else_if_acc_4_nl;
  assign nl_FpCmp_8U_23U_false_else_if_acc_6_nl[8:0] = FpCmp_8U_23U_false_else_if_acc_6_nl;
  assign nl_FpCmp_8U_23U_false_else_if_acc_8_nl[8:0] = FpCmp_8U_23U_false_else_if_acc_8_nl;
  assign nl_FpCmp_8U_23U_true_else_else_if_acc_4_nl[23:0] = FpCmp_8U_23U_true_else_else_if_acc_4_nl;
  assign nl_FpCmp_8U_23U_true_else_else_if_acc_6_nl[23:0] = FpCmp_8U_23U_true_else_else_if_acc_6_nl;
  assign nl_FpCmp_8U_23U_true_else_else_if_acc_7_nl[23:0] = FpCmp_8U_23U_true_else_else_if_acc_7_nl;
  assign nl_FpCmp_8U_23U_true_else_else_if_acc_8_nl[23:0] = FpCmp_8U_23U_true_else_else_if_acc_8_nl;
  assign nl_FpCmp_8U_23U_true_if_acc_10_nl[8:0] = FpCmp_8U_23U_true_if_acc_10_nl;
  assign nl_FpCmp_8U_23U_true_if_acc_4_nl[8:0] = FpCmp_8U_23U_true_if_acc_4_nl;
  assign nl_FpCmp_8U_23U_true_if_acc_6_nl[8:0] = FpCmp_8U_23U_true_if_acc_6_nl;
  assign nl_FpCmp_8U_23U_true_if_acc_8_nl[8:0] = FpCmp_8U_23U_true_if_acc_8_nl;
  assign nl_Y_alu_core_chn_alu_out_rsci_inst_chn_alu_out_rsci_d = { chn_alu_out_rsci_d_127, chn_alu_out_rsci_d_126_119, chn_alu_out_rsci_d_118_97, chn_alu_out_rsci_d_96, chn_alu_out_rsci_d_95, chn_alu_out_rsci_d_94_87, chn_alu_out_rsci_d_86_65, chn_alu_out_rsci_d_64, chn_alu_out_rsci_d_63, chn_alu_out_rsci_d_62_55, chn_alu_out_rsci_d_54_33, chn_alu_out_rsci_d_32, chn_alu_out_rsci_d_31, chn_alu_out_rsci_d_30_23, chn_alu_out_rsci_d_22_1, chn_alu_out_rsci_d_0 };
  assign nl_acc_10_nl[33:0] = acc_10_nl;
  assign nl_acc_11_nl[33:0] = acc_11_nl;
  assign nl_acc_12_nl[50:0] = acc_12_nl;
  assign nl_acc_13_nl[50:0] = acc_13_nl;
  assign nl_acc_14_nl[50:0] = acc_14_nl;
  assign nl_acc_15_nl[50:0] = acc_15_nl;
  assign nl_acc_1_nl[8:0] = acc_1_nl;
  assign nl_acc_2_nl[8:0] = acc_2_nl;
  assign nl_acc_3_nl[8:0] = acc_3_nl;
  assign nl_acc_4_nl[8:0] = acc_4_nl;
  assign nl_acc_5_nl[8:0] = acc_5_nl;
  assign nl_acc_6_nl[8:0] = acc_6_nl;
  assign nl_acc_7_nl[8:0] = acc_7_nl;
  assign nl_acc_8_nl[33:0] = acc_8_nl;
  assign nl_acc_9_nl[33:0] = acc_9_nl;
  assign nl_acc_nl[8:0] = acc_nl;
  assign nl_alu_loop_op_1_FpAdd_8U_23U_a_int_mant_p1_lshift_rg_a = { alu_loop_op_1_FpAdd_8U_23U_IsZero_8U_23U_or_itm_3, AluIn_data_sva_128[22:0] };
  assign nl_alu_loop_op_1_FpAdd_8U_23U_a_int_mant_p1_lshift_rg_s[8:1] = alu_loop_op_1_FpAdd_8U_23U_a_left_shift_acc_nl;
  assign nl_alu_loop_op_1_FpAdd_8U_23U_a_left_shift_acc_nl[7:0] = alu_loop_op_1_FpAdd_8U_23U_a_left_shift_acc_nl;
  assign nl_alu_loop_op_1_FpAdd_8U_23U_b_int_mant_p1_lshift_rg_a = { alu_loop_op_1_FpAdd_8U_23U_IsZero_8U_23U_1_or_itm_2, else_AluOp_data_0_lpi_1_dfm_2_30_0_1[22:0] };
  assign nl_alu_loop_op_1_FpAdd_8U_23U_b_int_mant_p1_lshift_rg_s[8:1] = alu_loop_op_1_FpAdd_8U_23U_b_left_shift_acc_nl;
  assign nl_alu_loop_op_1_FpAdd_8U_23U_b_left_shift_acc_nl[7:0] = alu_loop_op_1_FpAdd_8U_23U_b_left_shift_acc_nl;
  assign nl_alu_loop_op_1_FpAdd_8U_23U_if_3_if_acc_1_nl[7:0] = alu_loop_op_1_FpAdd_8U_23U_if_3_if_acc_1_nl;
  assign nl_alu_loop_op_1_FpAdd_8U_23U_if_4_if_acc_1_nl[7:0] = alu_loop_op_1_FpAdd_8U_23U_if_4_if_acc_1_nl;
  assign nl_alu_loop_op_1_FpAdd_8U_23U_if_4_if_acc_nl[7:0] = alu_loop_op_1_FpAdd_8U_23U_if_4_if_acc_nl;
  assign nl_alu_loop_op_1_FpMantRNE_49U_24U_else_acc_nl[22:0] = alu_loop_op_1_FpMantRNE_49U_24U_else_acc_nl;
  assign nl_alu_loop_op_1_FpNormalize_8U_49U_acc_nl[8:0] = alu_loop_op_1_FpNormalize_8U_49U_acc_nl;
  assign nl_alu_loop_op_1_FpNormalize_8U_49U_else_lshift_rg_a = FpAdd_8U_23U_int_mant_p1_1_lpi_1_dfm_5[48:0];
  assign nl_alu_loop_op_1_IntSaturation_33U_32U_else_if_acc_nl[2:0] = alu_loop_op_1_IntSaturation_33U_32U_else_if_acc_nl;
  assign nl_alu_loop_op_1_IntSaturation_33U_32U_if_acc_nl[2:0] = alu_loop_op_1_IntSaturation_33U_32U_if_acc_nl;
  assign nl_alu_loop_op_1_leading_sign_49_0_rg_mantissa = FpAdd_8U_23U_int_mant_p1_1_lpi_1_dfm_5[48:0];
  assign nl_alu_loop_op_2_FpAdd_8U_23U_a_int_mant_p1_lshift_2_rg_a = { alu_loop_op_2_FpAdd_8U_23U_IsZero_8U_23U_or_itm_4, AluIn_data_sva_128[54:32] };
  assign nl_alu_loop_op_2_FpAdd_8U_23U_a_int_mant_p1_lshift_2_rg_s[8:1] = alu_loop_op_2_FpAdd_8U_23U_a_left_shift_acc_2_nl;
  assign nl_alu_loop_op_2_FpAdd_8U_23U_a_left_shift_acc_2_nl[7:0] = alu_loop_op_2_FpAdd_8U_23U_a_left_shift_acc_2_nl;
  assign nl_alu_loop_op_2_FpAdd_8U_23U_b_int_mant_p1_lshift_2_rg_a = { alu_loop_op_2_FpAdd_8U_23U_IsZero_8U_23U_1_or_itm_2, else_AluOp_data_1_lpi_1_dfm_2_30_0_1[22:0] };
  assign nl_alu_loop_op_2_FpAdd_8U_23U_b_int_mant_p1_lshift_2_rg_s[8:1] = alu_loop_op_2_FpAdd_8U_23U_b_left_shift_acc_2_nl;
  assign nl_alu_loop_op_2_FpAdd_8U_23U_b_left_shift_acc_2_nl[7:0] = alu_loop_op_2_FpAdd_8U_23U_b_left_shift_acc_2_nl;
  assign nl_alu_loop_op_2_FpAdd_8U_23U_if_3_if_acc_4_nl[7:0] = alu_loop_op_2_FpAdd_8U_23U_if_3_if_acc_4_nl;
  assign nl_alu_loop_op_2_FpAdd_8U_23U_if_4_if_acc_4_nl[7:0] = alu_loop_op_2_FpAdd_8U_23U_if_4_if_acc_4_nl;
  assign nl_alu_loop_op_2_FpAdd_8U_23U_if_4_if_acc_5_nl[7:0] = alu_loop_op_2_FpAdd_8U_23U_if_4_if_acc_5_nl;
  assign nl_alu_loop_op_2_FpMantRNE_49U_24U_else_acc_2_nl[22:0] = alu_loop_op_2_FpMantRNE_49U_24U_else_acc_2_nl;
  assign nl_alu_loop_op_2_FpNormalize_8U_49U_acc_2_nl[8:0] = alu_loop_op_2_FpNormalize_8U_49U_acc_2_nl;
  assign nl_alu_loop_op_2_FpNormalize_8U_49U_else_lshift_2_rg_a = FpAdd_8U_23U_int_mant_p1_2_lpi_1_dfm_5[48:0];
  assign nl_alu_loop_op_2_IntSaturation_33U_32U_else_if_acc_1_nl[2:0] = alu_loop_op_2_IntSaturation_33U_32U_else_if_acc_1_nl;
  assign nl_alu_loop_op_2_IntSaturation_33U_32U_if_acc_1_nl[2:0] = alu_loop_op_2_IntSaturation_33U_32U_if_acc_1_nl;
  assign nl_alu_loop_op_2_leading_sign_49_0_2_rg_mantissa = FpAdd_8U_23U_int_mant_p1_2_lpi_1_dfm_5[48:0];
  assign nl_alu_loop_op_3_FpAdd_8U_23U_a_int_mant_p1_lshift_1_rg_a = { alu_loop_op_3_FpAdd_8U_23U_IsZero_8U_23U_or_itm_5, AluIn_data_sva_128[86:64] };
  assign nl_alu_loop_op_3_FpAdd_8U_23U_a_int_mant_p1_lshift_1_rg_s[8:1] = alu_loop_op_3_FpAdd_8U_23U_a_left_shift_acc_1_nl;
  assign nl_alu_loop_op_3_FpAdd_8U_23U_a_left_shift_acc_1_nl[7:0] = alu_loop_op_3_FpAdd_8U_23U_a_left_shift_acc_1_nl;
  assign nl_alu_loop_op_3_FpAdd_8U_23U_b_int_mant_p1_lshift_1_rg_a = { alu_loop_op_3_FpAdd_8U_23U_IsZero_8U_23U_1_or_itm_2, else_AluOp_data_2_lpi_1_dfm_2_30_0_1[22:0] };
  assign nl_alu_loop_op_3_FpAdd_8U_23U_b_int_mant_p1_lshift_1_rg_s[8:1] = alu_loop_op_3_FpAdd_8U_23U_b_left_shift_acc_1_nl;
  assign nl_alu_loop_op_3_FpAdd_8U_23U_b_left_shift_acc_1_nl[7:0] = alu_loop_op_3_FpAdd_8U_23U_b_left_shift_acc_1_nl;
  assign nl_alu_loop_op_3_FpAdd_8U_23U_if_3_if_acc_2_nl[7:0] = alu_loop_op_3_FpAdd_8U_23U_if_3_if_acc_2_nl;
  assign nl_alu_loop_op_3_FpAdd_8U_23U_if_4_if_acc_2_nl[7:0] = alu_loop_op_3_FpAdd_8U_23U_if_4_if_acc_2_nl;
  assign nl_alu_loop_op_3_FpAdd_8U_23U_if_4_if_acc_3_nl[7:0] = alu_loop_op_3_FpAdd_8U_23U_if_4_if_acc_3_nl;
  assign nl_alu_loop_op_3_FpMantRNE_49U_24U_else_acc_1_nl[22:0] = alu_loop_op_3_FpMantRNE_49U_24U_else_acc_1_nl;
  assign nl_alu_loop_op_3_FpNormalize_8U_49U_acc_1_nl[8:0] = alu_loop_op_3_FpNormalize_8U_49U_acc_1_nl;
  assign nl_alu_loop_op_3_FpNormalize_8U_49U_else_lshift_1_rg_a = FpAdd_8U_23U_int_mant_p1_3_lpi_1_dfm_5[48:0];
  assign nl_alu_loop_op_3_IntSaturation_33U_32U_else_if_acc_nl[2:0] = alu_loop_op_3_IntSaturation_33U_32U_else_if_acc_nl;
  assign nl_alu_loop_op_3_IntSaturation_33U_32U_if_acc_nl[2:0] = alu_loop_op_3_IntSaturation_33U_32U_if_acc_nl;
  assign nl_alu_loop_op_3_leading_sign_49_0_1_rg_mantissa = FpAdd_8U_23U_int_mant_p1_3_lpi_1_dfm_5[48:0];
  assign nl_alu_loop_op_4_FpAdd_8U_23U_a_int_mant_p1_lshift_3_rg_a = { alu_loop_op_4_FpAdd_8U_23U_IsZero_8U_23U_or_itm_5, AluIn_data_sva_128[118:96] };
  assign nl_alu_loop_op_4_FpAdd_8U_23U_a_int_mant_p1_lshift_3_rg_s[8:1] = alu_loop_op_4_FpAdd_8U_23U_a_left_shift_acc_3_nl;
  assign nl_alu_loop_op_4_FpAdd_8U_23U_a_left_shift_acc_3_nl[7:0] = alu_loop_op_4_FpAdd_8U_23U_a_left_shift_acc_3_nl;
  assign nl_alu_loop_op_4_FpAdd_8U_23U_b_int_mant_p1_lshift_3_rg_a = { alu_loop_op_4_FpAdd_8U_23U_IsZero_8U_23U_1_or_itm_2, else_AluOp_data_3_lpi_1_dfm_2_30_0_1[22:0] };
  assign nl_alu_loop_op_4_FpAdd_8U_23U_b_int_mant_p1_lshift_3_rg_s[8:1] = alu_loop_op_4_FpAdd_8U_23U_b_left_shift_acc_3_nl;
  assign nl_alu_loop_op_4_FpAdd_8U_23U_b_left_shift_acc_3_nl[7:0] = alu_loop_op_4_FpAdd_8U_23U_b_left_shift_acc_3_nl;
  assign nl_alu_loop_op_4_FpAdd_8U_23U_if_3_if_acc_6_nl[7:0] = alu_loop_op_4_FpAdd_8U_23U_if_3_if_acc_6_nl;
  assign nl_alu_loop_op_4_FpAdd_8U_23U_if_4_if_acc_6_nl[7:0] = alu_loop_op_4_FpAdd_8U_23U_if_4_if_acc_6_nl;
  assign nl_alu_loop_op_4_FpAdd_8U_23U_if_4_if_acc_7_nl[7:0] = alu_loop_op_4_FpAdd_8U_23U_if_4_if_acc_7_nl;
  assign nl_alu_loop_op_4_FpMantRNE_49U_24U_else_acc_3_nl[22:0] = alu_loop_op_4_FpMantRNE_49U_24U_else_acc_3_nl;
  assign nl_alu_loop_op_4_FpNormalize_8U_49U_acc_3_nl[8:0] = alu_loop_op_4_FpNormalize_8U_49U_acc_3_nl;
  assign nl_alu_loop_op_4_FpNormalize_8U_49U_else_lshift_3_rg_a = FpAdd_8U_23U_int_mant_p1_lpi_1_dfm_5[48:0];
  assign nl_alu_loop_op_4_IntSaturation_33U_32U_else_if_acc_1_nl[2:0] = alu_loop_op_4_IntSaturation_33U_32U_else_if_acc_1_nl;
  assign nl_alu_loop_op_4_IntSaturation_33U_32U_if_acc_1_nl[2:0] = alu_loop_op_4_IntSaturation_33U_32U_if_acc_1_nl;
  assign nl_alu_loop_op_4_leading_sign_49_0_3_rg_mantissa = FpAdd_8U_23U_int_mant_p1_lpi_1_dfm_5[48:0];
  assign nl_alu_loop_op_else_else_else_else_ac_int_cctor_1_sva[32:0] = alu_loop_op_else_else_else_else_ac_int_cctor_1_sva;
  assign nl_alu_loop_op_else_else_else_else_ac_int_cctor_2_sva[32:0] = alu_loop_op_else_else_else_else_ac_int_cctor_2_sva;
  assign nl_alu_loop_op_else_else_else_else_ac_int_cctor_3_sva[32:0] = alu_loop_op_else_else_else_else_ac_int_cctor_3_sva;
  assign nl_alu_loop_op_else_else_else_else_ac_int_cctor_sva[32:0] = alu_loop_op_else_else_else_else_ac_int_cctor_sva;
  assign or_937_cse = or_16_cse;
  assign z_out_12 = acc_12_nl[50:1];
  assign z_out_13 = acc_13_nl[50:1];
  assign z_out_14 = acc_14_nl[50:1];
  assign z_out_15 = acc_15_nl[50:1];
  assign z_out_4 = acc_4_nl[8:1];
  assign z_out_5 = acc_5_nl[8:1];
  assign z_out_6 = acc_6_nl[8:1];
  assign z_out_7 = acc_7_nl[8:1];
endmodule
