module aes_top_fifo(clk, rst, wr, addr, data_in, data_out, ack, stb, xram_data_in, aes_state, aes_addr, aes_len, aes_ctr, aes_key0, aes_step, addr_fifo_out, data_fifo_out, wr_fifo_out);
  logic [15:0] _0000_;
  logic [15:0] _0001_;
  logic [15:0] _0002_;
  logic [15:0] _0003_;
  logic [15:0] _0004_;
  logic [15:0] _0005_;
  logic [15:0] _0006_;
  logic [15:0] _0007_;
  logic [15:0] _0008_;
  logic [15:0] _0009_;
  logic [15:0] _0010_;
  logic [15:0] _0011_;
  logic [15:0] _0012_;
  logic [15:0] _0013_;
  logic [15:0] _0014_;
  logic [15:0] _0015_;
  logic [15:0] _0016_;
  logic [15:0] _0017_;
  logic [15:0] _0018_;
  logic [15:0] _0019_;
  logic [15:0] _0020_;
  logic [15:0] _0021_;
  logic [15:0] _0022_;
  logic [15:0] _0023_;
  logic [15:0] _0024_;
  logic [15:0] _0025_;
  logic [15:0] _0026_;
  logic [15:0] _0027_;
  logic [15:0] _0028_;
  logic [15:0] _0029_;
  logic [15:0] _0030_;
  logic [15:0] _0031_;
  logic [15:0] _0032_;
  logic [15:0] _0033_;
  logic [15:0] _0034_;
  logic [15:0] _0035_;
  logic [15:0] _0036_;
  logic [15:0] _0037_;
  logic [15:0] _0038_;
  logic [15:0] _0039_;
  logic [15:0] _0040_;
  logic [15:0] _0041_;
  logic [15:0] _0042_;
  logic [15:0] _0043_;
  logic [15:0] _0044_;
  logic [15:0] _0045_;
  logic [15:0] _0046_;
  logic [15:0] _0047_;
  logic [15:0] _0048_;
  logic [15:0] _0049_;
  logic [15:0] _0050_;
  logic [15:0] _0051_;
  logic [15:0] _0052_;
  logic [15:0] _0053_;
  logic [15:0] _0054_;
  logic [15:0] _0055_;
  logic [15:0] _0056_;
  logic [15:0] _0057_;
  logic [15:0] _0058_;
  logic [15:0] _0059_;
  logic [15:0] _0060_;
  logic [15:0] _0061_;
  logic [15:0] _0062_;
  logic [15:0] _0063_;
  logic [15:0] _0064_;
  logic [15:0] _0065_;
  logic [15:0] _0066_;
  logic [15:0] _0067_;
  logic [15:0] _0068_;
  logic [15:0] _0069_;
  logic [15:0] _0070_;
  logic [15:0] _0071_;
  logic [15:0] _0072_;
  logic [15:0] _0073_;
  logic [15:0] _0074_;
  logic [15:0] _0075_;
  logic [15:0] _0076_;
  logic [15:0] _0077_;
  logic [15:0] _0078_;
  logic [15:0] _0079_;
  logic [1:0] _0080_;
  logic [4:0] _0081_;
  logic [15:0] _0082_;
  logic [3:0] _0083_;
  logic [127:0] _0084_;
  logic [127:0] _0085_;
  logic [15:0] _0086_;
  logic [127:0] _0087_;
  logic [15:0] _0088_;
  logic [15:0] _0089_;
  logic [3:0] _0090_;
  logic [15:0] _0091_;
  logic [127:0] _0092_;
  logic [4:0] _0093_;
  logic [31:0] _0094_;
  logic [31:0] _0095_;
  logic [31:0] _0096_;
  logic _0097_;
  logic _0098_;
  logic _0099_;
  logic _0100_;
  logic _0101_;
  logic _0102_;
  logic _0103_;
  logic _0104_;
  logic _0105_;
  logic _0106_;
  logic _0107_;
  logic _0108_;
  logic _0109_;
  logic _0110_;
  logic _0111_;
  logic _0112_;
  logic _0113_;
  logic _0114_;
  logic _0115_;
  logic _0116_;
  logic _0117_;
  logic _0118_;
  logic _0119_;
  logic _0120_;
  logic _0121_;
  logic _0122_;
  logic _0123_;
  logic _0124_;
  logic _0125_;
  logic _0126_;
  logic _0127_;
  logic _0128_;
  logic _0129_;
  logic _0130_;
  logic _0131_;
  logic _0132_;
  logic _0133_;
  logic _0134_;
  logic _0135_;
  logic [7:0] _0136_;
  logic [7:0] _0137_;
  logic [7:0] _0138_;
  logic [7:0] _0139_;
  logic [1:0] _0140_;
  logic [1:0] _0141_;
  logic [1:0] _0142_;
  logic [1:0] _0143_;
  logic [127:0] _0144_;
  logic [4:0] _0145_;
  logic [7:0] _0146_;
  logic [7:0] _0147_;
  logic [7:0] _0148_;
  logic [7:0] _0149_;
  logic [7:0] _0150_;
  logic [7:0] _0151_;
  logic [7:0] _0152_;
  logic [7:0] _0153_;
  logic [7:0] _0154_;
  logic [7:0] _0155_;
  logic [7:0] _0156_;
  logic [7:0] _0157_;
  logic [7:0] _0158_;
  logic [7:0] _0159_;
  logic [127:0] _0160_;
  logic _0161_;
  logic _0162_;
  logic _0163_;
  logic _0164_;
  logic _0165_;
  logic _0166_;
  logic _0167_;
  logic _0168_;
  logic _0169_;
  logic _0170_;
  logic _0171_;
  logic _0172_;
  logic _0173_;
  logic _0174_;
  logic _0175_;
  logic _0176_;
  logic _0177_;
  logic [7:0] _0178_;
  logic [7:0] _0179_;
  logic [7:0] _0180_;
  logic [7:0] _0181_;
  logic [7:0] _0182_;
  logic [7:0] _0183_;
  logic [7:0] _0184_;
  logic [7:0] _0185_;
  logic [7:0] _0186_;
  logic [7:0] _0187_;
  logic [7:0] _0188_;
  logic [7:0] _0189_;
  logic [7:0] _0190_;
  logic [7:0] _0191_;
  logic [127:0] _0192_;
  logic _0193_;
  logic [7:0] _0194_;
  logic [7:0] _0195_;
  logic [7:0] _0196_;
  logic [7:0] _0197_;
  logic [7:0] _0198_;
  logic [7:0] _0199_;
  logic [7:0] _0200_;
  logic [7:0] _0201_;
  logic [7:0] _0202_;
  logic [7:0] _0203_;
  logic [7:0] _0204_;
  logic [7:0] _0205_;
  logic [7:0] _0206_;
  logic [7:0] _0207_;
  logic [15:0] _0208_;
  logic _0209_;
  logic _0210_;
  logic [15:0] _0211_;
  logic _0212_;
  logic [7:0] _0213_;
  logic [7:0] _0214_;
  logic [7:0] _0215_;
  logic [7:0] _0216_;
  logic [7:0] _0217_;
  logic [7:0] _0218_;
  logic [7:0] _0219_;
  logic [7:0] _0220_;
  logic [7:0] _0221_;
  logic [7:0] _0222_;
  logic [7:0] _0223_;
  logic [7:0] _0224_;
  logic [7:0] _0225_;
  logic [7:0] _0226_;
  logic [7:0] _0227_;
  logic [7:0] _0228_;
  logic [7:0] _0229_;
  logic [7:0] _0230_;
  logic [7:0] _0231_;
  logic [7:0] _0232_;
  logic [7:0] _0233_;
  logic [7:0] _0234_;
  logic [7:0] _0235_;
  logic [7:0] _0236_;
  logic [7:0] _0237_;
  logic [7:0] _0238_;
  logic [7:0] _0239_;
  logic [7:0] _0240_;
  logic [7:0] _0241_;
  logic [7:0] _0242_;
  logic [7:0] _0243_;
  logic [7:0] _0244_;
  logic [7:0] _0245_;
  logic [7:0] _0246_;
  logic [7:0] _0247_;
  logic [7:0] _0248_;
  logic [7:0] _0249_;
  logic [7:0] _0250_;
  logic [7:0] _0251_;
  logic [7:0] _0252_;
  logic [7:0] _0253_;
  logic [7:0] _0254_;
  logic [7:0] _0255_;
  logic [7:0] _0256_;
  logic [7:0] _0257_;
  logic [7:0] _0258_;
  logic [7:0] _0259_;
  logic [7:0] _0260_;
  logic [7:0] _0261_;
  logic [7:0] _0262_;
  logic [7:0] _0263_;
  logic [7:0] _0264_;
  logic [7:0] _0265_;
  logic [7:0] _0266_;
  logic [7:0] _0267_;
  logic [7:0] _0268_;
  logic [7:0] _0269_;
  logic [7:0] _0270_;
  logic [7:0] _0271_;
  logic [7:0] _0272_;
  logic [7:0] _0273_;
  logic [7:0] _0274_;
  logic [7:0] _0275_;
  logic [7:0] _0276_;
  logic [7:0] _0277_;
  logic [7:0] _0278_;
  logic [7:0] _0279_;
  logic [7:0] _0280_;
  logic [7:0] _0281_;
  logic [7:0] _0282_;
  logic [7:0] _0283_;
  logic [7:0] _0284_;
  logic [7:0] _0285_;
  logic [7:0] _0286_;
  logic [7:0] _0287_;
  logic [7:0] _0288_;
  logic [7:0] _0289_;
  logic [7:0] _0290_;
  logic [7:0] _0291_;
  logic [7:0] _0292_;
  logic _0293_;
  logic _0294_;
  logic _0295_;
  logic _0296_;
  logic _0297_;
  logic _0298_;
  logic _0299_;
  logic _0300_;
  logic _0301_;
  logic _0302_;
  logic _0303_;
  logic _0304_;
  logic _0305_;
  logic _0306_;
  logic _0307_;
  logic _0308_;
  logic _0309_;
  logic _0310_;
  logic _0311_;
  logic _0312_;
  logic _0313_;
  logic _0314_;
  logic _0315_;
  logic _0316_;
  logic _0317_;
  logic _0318_;
  logic _0319_;
  logic _0320_;
  logic _0321_;
  logic _0322_;
  logic _0323_;
  logic _0324_;
  logic _0325_;
  logic _0326_;
  logic _0327_;
  logic _0328_;
  logic _0329_;
  logic _0330_;
  logic _0331_;
  logic _0332_;
  logic _0333_;
  logic _0334_;
  logic _0335_;
  logic _0336_;
  logic _0337_;
  logic _0338_;
  logic _0339_;
  logic _0340_;
  logic _0341_;
  logic _0342_;
  logic _0343_;
  logic _0344_;
  logic _0345_;
  logic _0346_;
  logic _0347_;
  logic _0348_;
  logic _0349_;
  logic _0350_;
  logic _0351_;
  logic _0352_;
  logic _0353_;
  logic _0354_;
  logic _0355_;
  logic _0356_;
  logic _0357_;
  logic _0358_;
  logic _0359_;
  logic _0360_;
  logic _0361_;
  logic _0362_;
  logic _0363_;
  logic _0364_;
  logic _0365_;
  logic _0366_;
  logic _0367_;
  logic _0368_;
  logic _0369_;
  logic _0370_;
  logic _0371_;
  logic _0372_;
  output ack;
  input [15:0] addr;
  logic \addr_fifo.ack ;
  logic \addr_fifo.clk ;
  logic [15:0] \addr_fifo.in ;
  logic [15:0] \addr_fifo.out ;
  logic [15:0] \addr_fifo.r0 ;
  logic [15:0] \addr_fifo.r1 ;
  logic [15:0] \addr_fifo.r10 ;
  logic [15:0] \addr_fifo.r11 ;
  logic [15:0] \addr_fifo.r12 ;
  logic [15:0] \addr_fifo.r13 ;
  logic [15:0] \addr_fifo.r14 ;
  logic [15:0] \addr_fifo.r15 ;
  logic [15:0] \addr_fifo.r16 ;
  logic [15:0] \addr_fifo.r17 ;
  logic [15:0] \addr_fifo.r18 ;
  logic [15:0] \addr_fifo.r19 ;
  logic [15:0] \addr_fifo.r2 ;
  logic [15:0] \addr_fifo.r20 ;
  logic [15:0] \addr_fifo.r21 ;
  logic [15:0] \addr_fifo.r22 ;
  logic [15:0] \addr_fifo.r23 ;
  logic [15:0] \addr_fifo.r24 ;
  logic [15:0] \addr_fifo.r25 ;
  logic [15:0] \addr_fifo.r26 ;
  logic [15:0] \addr_fifo.r27 ;
  logic [15:0] \addr_fifo.r28 ;
  logic [15:0] \addr_fifo.r29 ;
  logic [15:0] \addr_fifo.r3 ;
  logic [15:0] \addr_fifo.r30 ;
  logic [15:0] \addr_fifo.r31 ;
  logic [15:0] \addr_fifo.r32 ;
  logic [15:0] \addr_fifo.r33 ;
  logic [15:0] \addr_fifo.r34 ;
  logic [15:0] \addr_fifo.r35 ;
  logic [15:0] \addr_fifo.r36 ;
  logic [15:0] \addr_fifo.r37 ;
  logic [15:0] \addr_fifo.r38 ;
  logic [15:0] \addr_fifo.r39 ;
  logic [15:0] \addr_fifo.r4 ;
  logic [15:0] \addr_fifo.r5 ;
  logic [15:0] \addr_fifo.r6 ;
  logic [15:0] \addr_fifo.r7 ;
  logic [15:0] \addr_fifo.r8 ;
  logic [15:0] \addr_fifo.r9 ;
  logic \addr_fifo.rst ;
  logic \addr_fifo.stb ;
  logic \addr_fifo.wr ;
  output [15:0] addr_fifo_out;
  output [15:0] aes_addr;
  output [127:0] aes_ctr;
  output [127:0] aes_key0;
  output [15:0] aes_len;
  output [1:0] aes_state;
  output aes_step;
  logic \aes_top_0.ack ;
  logic [15:0] \aes_top_0.addr ;
  logic [15:0] \aes_top_0.aes_addr ;
  logic [7:0] \aes_top_0.aes_addr_dataout ;
  logic [127:0] \aes_top_0.aes_ctr ;
  logic [7:0] \aes_top_0.aes_ctr_dataout ;
  logic [127:0] \aes_top_0.aes_curr_key ;
  logic [127:0] \aes_top_0.aes_key0 ;
  logic [7:0] \aes_top_0.aes_key0_dataout ;
  logic [15:0] \aes_top_0.aes_len ;
  logic [7:0] \aes_top_0.aes_len_dataout ;
  logic [127:0] \aes_top_0.aes_out ;
  logic [127:0] \aes_top_0.aes_reg_ctr ;
  logic [3:0] \aes_top_0.aes_reg_ctr_i.addr ;
  logic \aes_top_0.aes_reg_ctr_i.clk ;
  logic [7:0] \aes_top_0.aes_reg_ctr_i.data_in ;
  logic [7:0] \aes_top_0.aes_reg_ctr_i.data_out ;
  logic [7:0] \aes_top_0.aes_reg_ctr_i.data_out_mux ;
  logic \aes_top_0.aes_reg_ctr_i.en ;
  logic [7:0] \aes_top_0.aes_reg_ctr_i.reg0_next ;
  logic [7:0] \aes_top_0.aes_reg_ctr_i.reg10_next ;
  logic [7:0] \aes_top_0.aes_reg_ctr_i.reg11_next ;
  logic [7:0] \aes_top_0.aes_reg_ctr_i.reg12_next ;
  logic [7:0] \aes_top_0.aes_reg_ctr_i.reg13_next ;
  logic [7:0] \aes_top_0.aes_reg_ctr_i.reg14_next ;
  logic [7:0] \aes_top_0.aes_reg_ctr_i.reg15_next ;
  logic [7:0] \aes_top_0.aes_reg_ctr_i.reg1_next ;
  logic [7:0] \aes_top_0.aes_reg_ctr_i.reg2_next ;
  logic [7:0] \aes_top_0.aes_reg_ctr_i.reg3_next ;
  logic [7:0] \aes_top_0.aes_reg_ctr_i.reg4_next ;
  logic [7:0] \aes_top_0.aes_reg_ctr_i.reg5_next ;
  logic [7:0] \aes_top_0.aes_reg_ctr_i.reg6_next ;
  logic [7:0] \aes_top_0.aes_reg_ctr_i.reg7_next ;
  logic [7:0] \aes_top_0.aes_reg_ctr_i.reg8_next ;
  logic [7:0] \aes_top_0.aes_reg_ctr_i.reg9_next ;
  logic [127:0] \aes_top_0.aes_reg_ctr_i.reg_out ;
  logic \aes_top_0.aes_reg_ctr_i.rst ;
  logic \aes_top_0.aes_reg_ctr_i.wr ;
  logic \aes_top_0.aes_reg_ctr_i.wr0 ;
  logic \aes_top_0.aes_reg_ctr_i.wr1 ;
  logic \aes_top_0.aes_reg_ctr_i.wr10 ;
  logic \aes_top_0.aes_reg_ctr_i.wr11 ;
  logic \aes_top_0.aes_reg_ctr_i.wr12 ;
  logic \aes_top_0.aes_reg_ctr_i.wr13 ;
  logic \aes_top_0.aes_reg_ctr_i.wr14 ;
  logic \aes_top_0.aes_reg_ctr_i.wr15 ;
  logic \aes_top_0.aes_reg_ctr_i.wr2 ;
  logic \aes_top_0.aes_reg_ctr_i.wr3 ;
  logic \aes_top_0.aes_reg_ctr_i.wr4 ;
  logic \aes_top_0.aes_reg_ctr_i.wr5 ;
  logic \aes_top_0.aes_reg_ctr_i.wr6 ;
  logic \aes_top_0.aes_reg_ctr_i.wr7 ;
  logic \aes_top_0.aes_reg_ctr_i.wr8 ;
  logic \aes_top_0.aes_reg_ctr_i.wr9 ;
  logic [127:0] \aes_top_0.aes_reg_key0 ;
  logic [3:0] \aes_top_0.aes_reg_key0_i.addr ;
  logic \aes_top_0.aes_reg_key0_i.clk ;
  logic [7:0] \aes_top_0.aes_reg_key0_i.data_in ;
  logic [7:0] \aes_top_0.aes_reg_key0_i.data_out ;
  logic [7:0] \aes_top_0.aes_reg_key0_i.data_out_mux ;
  logic \aes_top_0.aes_reg_key0_i.en ;
  logic [7:0] \aes_top_0.aes_reg_key0_i.reg0_next ;
  logic [7:0] \aes_top_0.aes_reg_key0_i.reg10_next ;
  logic [7:0] \aes_top_0.aes_reg_key0_i.reg11_next ;
  logic [7:0] \aes_top_0.aes_reg_key0_i.reg12_next ;
  logic [7:0] \aes_top_0.aes_reg_key0_i.reg13_next ;
  logic [7:0] \aes_top_0.aes_reg_key0_i.reg14_next ;
  logic [7:0] \aes_top_0.aes_reg_key0_i.reg15_next ;
  logic [7:0] \aes_top_0.aes_reg_key0_i.reg1_next ;
  logic [7:0] \aes_top_0.aes_reg_key0_i.reg2_next ;
  logic [7:0] \aes_top_0.aes_reg_key0_i.reg3_next ;
  logic [7:0] \aes_top_0.aes_reg_key0_i.reg4_next ;
  logic [7:0] \aes_top_0.aes_reg_key0_i.reg5_next ;
  logic [7:0] \aes_top_0.aes_reg_key0_i.reg6_next ;
  logic [7:0] \aes_top_0.aes_reg_key0_i.reg7_next ;
  logic [7:0] \aes_top_0.aes_reg_key0_i.reg8_next ;
  logic [7:0] \aes_top_0.aes_reg_key0_i.reg9_next ;
  logic [127:0] \aes_top_0.aes_reg_key0_i.reg_out ;
  logic \aes_top_0.aes_reg_key0_i.rst ;
  logic \aes_top_0.aes_reg_key0_i.wr ;
  logic \aes_top_0.aes_reg_key0_i.wr0 ;
  logic \aes_top_0.aes_reg_key0_i.wr1 ;
  logic \aes_top_0.aes_reg_key0_i.wr10 ;
  logic \aes_top_0.aes_reg_key0_i.wr11 ;
  logic \aes_top_0.aes_reg_key0_i.wr12 ;
  logic \aes_top_0.aes_reg_key0_i.wr13 ;
  logic \aes_top_0.aes_reg_key0_i.wr14 ;
  logic \aes_top_0.aes_reg_key0_i.wr15 ;
  logic \aes_top_0.aes_reg_key0_i.wr2 ;
  logic \aes_top_0.aes_reg_key0_i.wr3 ;
  logic \aes_top_0.aes_reg_key0_i.wr4 ;
  logic \aes_top_0.aes_reg_key0_i.wr5 ;
  logic \aes_top_0.aes_reg_key0_i.wr6 ;
  logic \aes_top_0.aes_reg_key0_i.wr7 ;
  logic \aes_top_0.aes_reg_key0_i.wr8 ;
  logic \aes_top_0.aes_reg_key0_i.wr9 ;
  logic [15:0] \aes_top_0.aes_reg_opaddr ;
  logic \aes_top_0.aes_reg_opaddr_i.addr ;
  logic \aes_top_0.aes_reg_opaddr_i.clk ;
  logic [7:0] \aes_top_0.aes_reg_opaddr_i.data_in ;
  logic [7:0] \aes_top_0.aes_reg_opaddr_i.data_out ;
  logic [7:0] \aes_top_0.aes_reg_opaddr_i.data_out_mux ;
  logic \aes_top_0.aes_reg_opaddr_i.en ;
  logic [7:0] \aes_top_0.aes_reg_opaddr_i.reg0_next ;
  logic [7:0] \aes_top_0.aes_reg_opaddr_i.reg1_next ;
  logic [15:0] \aes_top_0.aes_reg_opaddr_i.reg_out ;
  logic \aes_top_0.aes_reg_opaddr_i.rst ;
  logic \aes_top_0.aes_reg_opaddr_i.wr ;
  logic \aes_top_0.aes_reg_opaddr_i.wr0 ;
  logic \aes_top_0.aes_reg_opaddr_i.wr1 ;
  logic [15:0] \aes_top_0.aes_reg_oplen ;
  logic \aes_top_0.aes_reg_oplen_i.addr ;
  logic \aes_top_0.aes_reg_oplen_i.clk ;
  logic [7:0] \aes_top_0.aes_reg_oplen_i.data_in ;
  logic [7:0] \aes_top_0.aes_reg_oplen_i.data_out ;
  logic [7:0] \aes_top_0.aes_reg_oplen_i.data_out_mux ;
  logic \aes_top_0.aes_reg_oplen_i.en ;
  logic [7:0] \aes_top_0.aes_reg_oplen_i.reg0_next ;
  logic [7:0] \aes_top_0.aes_reg_oplen_i.reg1_next ;
  logic [15:0] \aes_top_0.aes_reg_oplen_i.reg_out ;
  logic \aes_top_0.aes_reg_oplen_i.rst ;
  logic \aes_top_0.aes_reg_oplen_i.wr ;
  logic \aes_top_0.aes_reg_oplen_i.wr0 ;
  logic \aes_top_0.aes_reg_oplen_i.wr1 ;
  logic [1:0] \aes_top_0.aes_reg_state ;
  logic [1:0] \aes_top_0.aes_reg_state_next ;
  logic \aes_top_0.aes_reg_state_next_idle ;
  logic \aes_top_0.aes_reg_state_next_operate ;
  logic [1:0] \aes_top_0.aes_reg_state_next_read_data ;
  logic [1:0] \aes_top_0.aes_reg_state_next_write_data ;
  logic [1:0] \aes_top_0.aes_state ;
  logic \aes_top_0.aes_state_idle ;
  logic \aes_top_0.aes_state_operate ;
  logic \aes_top_0.aes_state_read_data ;
  logic \aes_top_0.aes_state_write_data ;
  logic \aes_top_0.aes_step ;
  logic [4:0] \aes_top_0.aes_time_counter ;
  logic [4:0] \aes_top_0.aes_time_counter_next ;
  logic \aes_top_0.aes_time_enough ;
  logic [15:0] \aes_top_0.block_counter ;
  logic [15:0] \aes_top_0.block_counter_next ;
  logic [3:0] \aes_top_0.byte_counter ;
  logic [3:0] \aes_top_0.byte_counter_next ;
  logic \aes_top_0.clk ;
  logic [7:0] \aes_top_0.data_in ;
  logic [7:0] \aes_top_0.data_out ;
  logic [127:0] \aes_top_0.encrypted_data ;
  logic [127:0] \aes_top_0.encrypted_data_buf ;
  logic [127:0] \aes_top_0.encrypted_data_buf_next ;
  logic \aes_top_0.in_addr_range ;
  logic \aes_top_0.incr_byte_counter ;
  logic \aes_top_0.last_byte_acked ;
  logic [127:0] \aes_top_0.mem_data_buf ;
  logic [127:0] \aes_top_0.mem_data_buf_next ;
  logic \aes_top_0.more_blocks ;
  logic [15:0] \aes_top_0.operated_bytes_count ;
  logic [15:0] \aes_top_0.operated_bytes_count_next ;
  logic \aes_top_0.reset_byte_counter ;
  logic \aes_top_0.rst ;
  logic \aes_top_0.sel_reg_addr ;
  logic \aes_top_0.sel_reg_ctr ;
  logic \aes_top_0.sel_reg_key0 ;
  logic \aes_top_0.sel_reg_len ;
  logic \aes_top_0.sel_reg_start ;
  logic \aes_top_0.sel_reg_state ;
  logic \aes_top_0.start_op ;
  logic \aes_top_0.stb ;
  logic [127:0] \aes_top_0.uaes_ctr ;
  logic [127:0] \aes_top_0.uaes_ctr_nxt ;
  logic \aes_top_0.wr ;
  logic \aes_top_0.wren ;
  logic \aes_top_0.xram_ack ;
  logic [15:0] \aes_top_0.xram_addr ;
  logic [7:0] \aes_top_0.xram_data_in ;
  logic [7:0] \aes_top_0.xram_data_out ;
  logic \aes_top_0.xram_stb ;
  logic \aes_top_0.xram_wr ;
  input clk;
  logic \data_fifo.ack ;
  logic \data_fifo.clk ;
  logic [7:0] \data_fifo.in ;
  logic [7:0] \data_fifo.out ;
  logic [7:0] \data_fifo.r0 ;
  logic [7:0] \data_fifo.r1 ;
  logic [7:0] \data_fifo.r10 ;
  logic [7:0] \data_fifo.r11 ;
  logic [7:0] \data_fifo.r12 ;
  logic [7:0] \data_fifo.r13 ;
  logic [7:0] \data_fifo.r14 ;
  logic [7:0] \data_fifo.r15 ;
  logic [7:0] \data_fifo.r16 ;
  logic [7:0] \data_fifo.r17 ;
  logic [7:0] \data_fifo.r18 ;
  logic [7:0] \data_fifo.r19 ;
  logic [7:0] \data_fifo.r2 ;
  logic [7:0] \data_fifo.r20 ;
  logic [7:0] \data_fifo.r21 ;
  logic [7:0] \data_fifo.r22 ;
  logic [7:0] \data_fifo.r23 ;
  logic [7:0] \data_fifo.r24 ;
  logic [7:0] \data_fifo.r25 ;
  logic [7:0] \data_fifo.r26 ;
  logic [7:0] \data_fifo.r27 ;
  logic [7:0] \data_fifo.r28 ;
  logic [7:0] \data_fifo.r29 ;
  logic [7:0] \data_fifo.r3 ;
  logic [7:0] \data_fifo.r30 ;
  logic [7:0] \data_fifo.r31 ;
  logic [7:0] \data_fifo.r32 ;
  logic [7:0] \data_fifo.r33 ;
  logic [7:0] \data_fifo.r34 ;
  logic [7:0] \data_fifo.r35 ;
  logic [7:0] \data_fifo.r36 ;
  logic [7:0] \data_fifo.r37 ;
  logic [7:0] \data_fifo.r38 ;
  logic [7:0] \data_fifo.r39 ;
  logic [7:0] \data_fifo.r4 ;
  logic [7:0] \data_fifo.r5 ;
  logic [7:0] \data_fifo.r6 ;
  logic [7:0] \data_fifo.r7 ;
  logic [7:0] \data_fifo.r8 ;
  logic [7:0] \data_fifo.r9 ;
  logic \data_fifo.rst ;
  logic \data_fifo.stb ;
  logic \data_fifo.wr ;
  output [7:0] data_fifo_out;
  input [7:0] data_in;
  output [7:0] data_out;
  input rst;
  input stb;
  input wr;
  logic \wr_fifo.ack ;
  logic \wr_fifo.clk ;
  logic \wr_fifo.in ;
  logic \wr_fifo.out ;
  logic \wr_fifo.r0 ;
  logic \wr_fifo.r1 ;
  logic \wr_fifo.r10 ;
  logic \wr_fifo.r11 ;
  logic \wr_fifo.r12 ;
  logic \wr_fifo.r13 ;
  logic \wr_fifo.r14 ;
  logic \wr_fifo.r15 ;
  logic \wr_fifo.r16 ;
  logic \wr_fifo.r17 ;
  logic \wr_fifo.r18 ;
  logic \wr_fifo.r19 ;
  logic \wr_fifo.r2 ;
  logic \wr_fifo.r20 ;
  logic \wr_fifo.r21 ;
  logic \wr_fifo.r22 ;
  logic \wr_fifo.r23 ;
  logic \wr_fifo.r24 ;
  logic \wr_fifo.r25 ;
  logic \wr_fifo.r26 ;
  logic \wr_fifo.r27 ;
  logic \wr_fifo.r28 ;
  logic \wr_fifo.r29 ;
  logic \wr_fifo.r3 ;
  logic \wr_fifo.r30 ;
  logic \wr_fifo.r31 ;
  logic \wr_fifo.r32 ;
  logic \wr_fifo.r33 ;
  logic \wr_fifo.r34 ;
  logic \wr_fifo.r35 ;
  logic \wr_fifo.r36 ;
  logic \wr_fifo.r37 ;
  logic \wr_fifo.r38 ;
  logic \wr_fifo.r39 ;
  logic \wr_fifo.r4 ;
  logic \wr_fifo.r5 ;
  logic \wr_fifo.r6 ;
  logic \wr_fifo.r7 ;
  logic \wr_fifo.r8 ;
  logic \wr_fifo.r9 ;
  logic \wr_fifo.rst ;
  logic \wr_fifo.stb ;
  logic \wr_fifo.wr ;
  output wr_fifo_out;
  logic xram_ack;
  logic [15:0] xram_addr;
  input [7:0] xram_data_in;
  logic [7:0] xram_data_out;
  logic xram_stb;
  logic xram_wr;
  always @(posedge clk)
      \addr_fifo.r1 <= _0011_;
  always @(posedge clk)
      \addr_fifo.r2 <= _0022_;
  always @(posedge clk)
      \addr_fifo.r3 <= _0033_;
  always @(posedge clk)
      \addr_fifo.r4 <= _0034_;
  always @(posedge clk)
      \addr_fifo.r5 <= _0035_;
  always @(posedge clk)
      \addr_fifo.r6 <= _0036_;
  always @(posedge clk)
      \addr_fifo.r7 <= _0037_;
  always @(posedge clk)
      \addr_fifo.r8 <= _0038_;
  always @(posedge clk)
      \addr_fifo.r9 <= _0039_;
  always @(posedge clk)
      \addr_fifo.r0 <= _0000_;
  always @(posedge clk)
      \addr_fifo.r10 <= _0001_;
  always @(posedge clk)
      \addr_fifo.r11 <= _0002_;
  always @(posedge clk)
      \addr_fifo.r12 <= _0003_;
  always @(posedge clk)
      \addr_fifo.r13 <= _0004_;
  always @(posedge clk)
      \addr_fifo.r14 <= _0005_;
  always @(posedge clk)
      \addr_fifo.r15 <= _0006_;
  always @(posedge clk)
      \addr_fifo.r16 <= _0007_;
  always @(posedge clk)
      \addr_fifo.r17 <= _0008_;
  always @(posedge clk)
      \addr_fifo.r18 <= _0009_;
  always @(posedge clk)
      \addr_fifo.r19 <= _0010_;
  always @(posedge clk)
      \addr_fifo.r20 <= _0012_;
  always @(posedge clk)
      \addr_fifo.r21 <= _0013_;
  always @(posedge clk)
      \addr_fifo.r22 <= _0014_;
  always @(posedge clk)
      \addr_fifo.r23 <= _0015_;
  always @(posedge clk)
      \addr_fifo.r24 <= _0016_;
  always @(posedge clk)
      \addr_fifo.r25 <= _0017_;
  always @(posedge clk)
      \addr_fifo.r26 <= _0018_;
  always @(posedge clk)
      \addr_fifo.r27 <= _0019_;
  always @(posedge clk)
      \addr_fifo.r28 <= _0020_;
  always @(posedge clk)
      \addr_fifo.r29 <= _0021_;
  always @(posedge clk)
      \addr_fifo.r30 <= _0023_;
  always @(posedge clk)
      \addr_fifo.r31 <= _0024_;
  always @(posedge clk)
      \addr_fifo.r32 <= _0025_;
  always @(posedge clk)
      \addr_fifo.r33 <= _0026_;
  always @(posedge clk)
      \addr_fifo.r34 <= _0027_;
  always @(posedge clk)
      \addr_fifo.r35 <= _0028_;
  always @(posedge clk)
      \addr_fifo.r36 <= _0029_;
  always @(posedge clk)
      \addr_fifo.r37 <= _0030_;
  always @(posedge clk)
      \addr_fifo.r38 <= _0031_;
  always @(posedge clk)
      \addr_fifo.r39 <= _0032_;
  assign _0040_ = \addr_fifo.wr ? \addr_fifo.r38 : \addr_fifo.r39 ;
  assign _0032_ = rst ? 16'b0000000000000000 : _0040_;
  assign _0041_ = \addr_fifo.wr ? \addr_fifo.r37 : \addr_fifo.r38 ;
  assign _0031_ = rst ? 16'b0000000000000000 : _0041_;
  assign _0042_ = \addr_fifo.wr ? \addr_fifo.r36 : \addr_fifo.r37 ;
  assign _0030_ = rst ? 16'b0000000000000000 : _0042_;
  assign _0043_ = \addr_fifo.wr ? \addr_fifo.r35 : \addr_fifo.r36 ;
  assign _0029_ = rst ? 16'b0000000000000000 : _0043_;
  assign _0044_ = \addr_fifo.wr ? \addr_fifo.r34 : \addr_fifo.r35 ;
  assign _0028_ = rst ? 16'b0000000000000000 : _0044_;
  assign _0045_ = \addr_fifo.wr ? \addr_fifo.r33 : \addr_fifo.r34 ;
  assign _0027_ = rst ? 16'b0000000000000000 : _0045_;
  assign _0046_ = \addr_fifo.wr ? \addr_fifo.r32 : \addr_fifo.r33 ;
  assign _0026_ = rst ? 16'b0000000000000000 : _0046_;
  assign _0047_ = \addr_fifo.wr ? \addr_fifo.r31 : \addr_fifo.r32 ;
  assign _0025_ = rst ? 16'b0000000000000000 : _0047_;
  assign _0048_ = \addr_fifo.wr ? \addr_fifo.r30 : \addr_fifo.r31 ;
  assign _0024_ = rst ? 16'b0000000000000000 : _0048_;
  assign _0049_ = \addr_fifo.wr ? \addr_fifo.r29 : \addr_fifo.r30 ;
  assign _0023_ = rst ? 16'b0000000000000000 : _0049_;
  assign _0050_ = \addr_fifo.wr ? \addr_fifo.r28 : \addr_fifo.r29 ;
  assign _0021_ = rst ? 16'b0000000000000000 : _0050_;
  assign _0051_ = \addr_fifo.wr ? \addr_fifo.r27 : \addr_fifo.r28 ;
  assign _0020_ = rst ? 16'b0000000000000000 : _0051_;
  assign _0052_ = \addr_fifo.wr ? \addr_fifo.r26 : \addr_fifo.r27 ;
  assign _0019_ = rst ? 16'b0000000000000000 : _0052_;
  assign _0053_ = \addr_fifo.wr ? \addr_fifo.r25 : \addr_fifo.r26 ;
  assign _0018_ = rst ? 16'b0000000000000000 : _0053_;
  assign _0054_ = \addr_fifo.wr ? \addr_fifo.r24 : \addr_fifo.r25 ;
  assign _0017_ = rst ? 16'b0000000000000000 : _0054_;
  assign _0055_ = \addr_fifo.wr ? \addr_fifo.r23 : \addr_fifo.r24 ;
  assign _0016_ = rst ? 16'b0000000000000000 : _0055_;
  assign _0056_ = \addr_fifo.wr ? \addr_fifo.r22 : \addr_fifo.r23 ;
  assign _0015_ = rst ? 16'b0000000000000000 : _0056_;
  assign _0057_ = \addr_fifo.wr ? \addr_fifo.r21 : \addr_fifo.r22 ;
  assign _0014_ = rst ? 16'b0000000000000000 : _0057_;
  assign _0058_ = \addr_fifo.wr ? \addr_fifo.r20 : \addr_fifo.r21 ;
  assign _0013_ = rst ? 16'b0000000000000000 : _0058_;
  assign _0059_ = \addr_fifo.wr ? \addr_fifo.r19 : \addr_fifo.r20 ;
  assign _0012_ = rst ? 16'b0000000000000000 : _0059_;
  assign _0060_ = \addr_fifo.wr ? \addr_fifo.r18 : \addr_fifo.r19 ;
  assign _0010_ = rst ? 16'b0000000000000000 : _0060_;
  assign _0061_ = \addr_fifo.wr ? \addr_fifo.r17 : \addr_fifo.r18 ;
  assign _0009_ = rst ? 16'b0000000000000000 : _0061_;
  assign _0062_ = \addr_fifo.wr ? \addr_fifo.r16 : \addr_fifo.r17 ;
  assign _0008_ = rst ? 16'b0000000000000000 : _0062_;
  assign _0063_ = \addr_fifo.wr ? \addr_fifo.r15 : \addr_fifo.r16 ;
  assign _0007_ = rst ? 16'b0000000000000000 : _0063_;
  assign _0064_ = \addr_fifo.wr ? \addr_fifo.r14 : \addr_fifo.r15 ;
  assign _0006_ = rst ? 16'b0000000000000000 : _0064_;
  assign _0065_ = \addr_fifo.wr ? \addr_fifo.r13 : \addr_fifo.r14 ;
  assign _0005_ = rst ? 16'b0000000000000000 : _0065_;
  assign _0066_ = \addr_fifo.wr ? \addr_fifo.r12 : \addr_fifo.r13 ;
  assign _0004_ = rst ? 16'b0000000000000000 : _0066_;
  assign _0067_ = \addr_fifo.wr ? \addr_fifo.r11 : \addr_fifo.r12 ;
  assign _0003_ = rst ? 16'b0000000000000000 : _0067_;
  assign _0068_ = \addr_fifo.wr ? \addr_fifo.r10 : \addr_fifo.r11 ;
  assign _0002_ = rst ? 16'b0000000000000000 : _0068_;
  assign _0069_ = \addr_fifo.wr ? \addr_fifo.r9 : \addr_fifo.r10 ;
  assign _0001_ = rst ? 16'b0000000000000000 : _0069_;
  assign _0070_ = \addr_fifo.wr ? \addr_fifo.in : \addr_fifo.r0 ;
  assign _0000_ = rst ? 16'b0000000000000000 : _0070_;
  assign _0071_ = \addr_fifo.wr ? \addr_fifo.r8 : \addr_fifo.r9 ;
  assign _0039_ = rst ? 16'b0000000000000000 : _0071_;
  assign _0072_ = \addr_fifo.wr ? \addr_fifo.r7 : \addr_fifo.r8 ;
  assign _0038_ = rst ? 16'b0000000000000000 : _0072_;
  assign _0073_ = \addr_fifo.wr ? \addr_fifo.r6 : \addr_fifo.r7 ;
  assign _0037_ = rst ? 16'b0000000000000000 : _0073_;
  assign _0074_ = \addr_fifo.wr ? \addr_fifo.r5 : \addr_fifo.r6 ;
  assign _0036_ = rst ? 16'b0000000000000000 : _0074_;
  assign _0075_ = \addr_fifo.wr ? \addr_fifo.r4 : \addr_fifo.r5 ;
  assign _0035_ = rst ? 16'b0000000000000000 : _0075_;
  assign _0076_ = \addr_fifo.wr ? \addr_fifo.r3 : \addr_fifo.r4 ;
  assign _0034_ = rst ? 16'b0000000000000000 : _0076_;
  assign _0077_ = \addr_fifo.wr ? \addr_fifo.r2 : \addr_fifo.r3 ;
  assign _0033_ = rst ? 16'b0000000000000000 : _0077_;
  assign _0078_ = \addr_fifo.wr ? \addr_fifo.r1 : \addr_fifo.r2 ;
  assign _0022_ = rst ? 16'b0000000000000000 : _0078_;
  assign _0079_ = \addr_fifo.wr ? \addr_fifo.r0 : \addr_fifo.r1 ;
  assign _0011_ = rst ? 16'b0000000000000000 : _0079_;
  assign _0088_ = \aes_top_0.operated_bytes_count + 5'b10000;
  assign _0089_ = \aes_top_0.block_counter + 5'b10000;
  assign _0090_ = \aes_top_0.byte_counter + 1'b1;
  assign _0091_ = \aes_top_0.aes_reg_opaddr_i.reg_out + \aes_top_0.block_counter ;
  assign \addr_fifo.in = _0091_ + \aes_top_0.byte_counter ;
  assign _0092_ = \aes_top_0.uaes_ctr + 5'b10000;
  assign _0093_ = \aes_top_0.aes_time_counter + 1'b1;
  assign \aes_top_0.sel_reg_start = addr == 16'b1111111100000000;
  assign \aes_top_0.sel_reg_state = addr == 16'b1111111100000001;
  assign \aes_top_0.aes_reg_opaddr_i.en = addr[15:1] == 15'b111111110000001;
  assign \aes_top_0.aes_reg_oplen_i.en = addr[15:1] == 15'b111111110000010;
  assign \aes_top_0.aes_reg_ctr_i.en = addr[15:4] == 12'b111111110010;
  assign \aes_top_0.aes_reg_key0_i.en = addr[15:4] == 12'b111111110001;
  assign \aes_top_0.aes_state_idle = ! \aes_top_0.aes_reg_state ;
  assign \aes_top_0.aes_state_read_data = \aes_top_0.aes_reg_state == 1'b1;
  assign \aes_top_0.aes_state_operate = \aes_top_0.aes_reg_state == 2'b10;
  assign \addr_fifo.wr = \aes_top_0.aes_reg_state == 2'b11;
  assign _0097_ = \aes_top_0.byte_counter == 4'b1111;
  assign _0098_ = ! \aes_top_0.byte_counter ;
  assign _0099_ = \aes_top_0.byte_counter == 1'b1;
  assign _0100_ = \aes_top_0.byte_counter == 2'b10;
  assign _0101_ = \aes_top_0.byte_counter == 2'b11;
  assign _0102_ = \aes_top_0.byte_counter == 3'b100;
  assign _0103_ = \aes_top_0.byte_counter == 3'b101;
  assign _0104_ = \aes_top_0.byte_counter == 3'b110;
  assign _0105_ = \aes_top_0.byte_counter == 3'b111;
  assign _0106_ = \aes_top_0.byte_counter == 4'b1000;
  assign _0107_ = \aes_top_0.byte_counter == 4'b1001;
  assign _0108_ = \aes_top_0.byte_counter == 4'b1010;
  assign _0109_ = \aes_top_0.byte_counter == 4'b1011;
  assign _0110_ = \aes_top_0.byte_counter == 4'b1100;
  assign _0111_ = \aes_top_0.byte_counter == 4'b1101;
  assign _0112_ = \aes_top_0.byte_counter == 4'b1110;
  assign _0113_ = addr >= 16'b1111111100000000;
  assign \aes_top_0.aes_time_enough = \aes_top_0.aes_time_counter >= 5'b10101;
  assign \aes_top_0.in_addr_range = _0113_ && _0133_;
  assign \aes_top_0.ack = stb && \aes_top_0.in_addr_range ;
  assign \aes_top_0.wren = wr && \aes_top_0.aes_state_idle ;
  assign _0114_ = \aes_top_0.sel_reg_start && data_in[0];
  assign \aes_top_0.reset_byte_counter = _0114_ && \aes_top_0.wren ;
  assign \aes_top_0.aes_reg_opaddr_i.wr = \aes_top_0.aes_reg_opaddr_i.en && \aes_top_0.wren ;
  assign \aes_top_0.aes_reg_oplen_i.wr = \aes_top_0.aes_reg_oplen_i.en && \aes_top_0.wren ;
  assign \aes_top_0.aes_reg_ctr_i.wr = \aes_top_0.aes_reg_ctr_i.en && \aes_top_0.wren ;
  assign \aes_top_0.aes_reg_key0_i.wr = \aes_top_0.aes_reg_key0_i.en && \aes_top_0.wren ;
  assign _0115_ = \aes_top_0.last_byte_acked && \addr_fifo.wr ;
  assign \aes_top_0.last_byte_acked = _0097_ && \aes_top_0.xram_ack ;
  assign \aes_top_0.more_blocks = _0115_ && _0134_;
  assign _0116_ = \aes_top_0.last_byte_acked && \aes_top_0.more_blocks ;
  assign _0117_ = \aes_top_0.xram_ack && _0098_;
  assign _0118_ = \aes_top_0.xram_ack && _0099_;
  assign _0119_ = \aes_top_0.xram_ack && _0100_;
  assign _0120_ = \aes_top_0.xram_ack && _0101_;
  assign _0121_ = \aes_top_0.xram_ack && _0102_;
  assign _0122_ = \aes_top_0.xram_ack && _0103_;
  assign _0123_ = \aes_top_0.xram_ack && _0104_;
  assign _0124_ = \aes_top_0.xram_ack && _0105_;
  assign _0125_ = \aes_top_0.xram_ack && _0106_;
  assign _0126_ = \aes_top_0.xram_ack && _0107_;
  assign _0127_ = \aes_top_0.xram_ack && _0108_;
  assign _0128_ = \aes_top_0.xram_ack && _0109_;
  assign _0129_ = \aes_top_0.xram_ack && _0110_;
  assign _0130_ = \aes_top_0.xram_ack && _0111_;
  assign _0131_ = \aes_top_0.xram_ack && _0112_;
  assign \aes_top_0.xram_ack = \aes_top_0.aes_state_read_data || \addr_fifo.wr ;
  assign _0132_ = \aes_top_0.more_blocks || \aes_top_0.reset_byte_counter ;
  assign _0133_ = addr < 16'b1111111100110000;
  assign _0134_ = \aes_top_0.operated_bytes_count_next < \aes_top_0.aes_reg_oplen_i.reg_out ;
  assign _0135_ = \aes_top_0.aes_time_counter < 5'b11111;
  assign \aes_top_0.aes_step = \aes_top_0.aes_reg_state != \aes_top_0.aes_reg_state_next ;
  always @(posedge clk)
      \aes_top_0.aes_reg_state <= _0080_;
  always @(posedge clk)
      \aes_top_0.operated_bytes_count <= _0086_;
  always @(posedge clk)
      \aes_top_0.block_counter <= _0082_;
  always @(posedge clk)
      \aes_top_0.byte_counter <= _0083_;
  always @(posedge clk)
      \aes_top_0.mem_data_buf <= _0085_;
  always @(posedge clk)
      \aes_top_0.encrypted_data_buf <= _0084_;
  always @(posedge clk)
      \aes_top_0.aes_time_counter <= _0081_;
  always @(posedge clk)
      \aes_top_0.uaes_ctr <= _0087_;
  assign _0084_ = rst ? \aes_top_0.encrypted_data_buf : \aes_top_0.encrypted_data_buf_next ;
  assign _0085_ = rst ? \aes_top_0.mem_data_buf : \aes_top_0.mem_data_buf_next ;
  assign _0083_ = rst ? 4'b0000 : \aes_top_0.byte_counter_next ;
  assign _0082_ = rst ? 16'b0000000000000000 : \aes_top_0.block_counter_next ;
  assign _0086_ = rst ? 16'b0000000000000000 : \aes_top_0.operated_bytes_count_next ;
  assign _0080_ = rst ? 2'b00 : \aes_top_0.aes_reg_state_next ;
  assign _0081_ = rst ? 5'b00000 : \aes_top_0.aes_time_counter_next ;
  assign _0087_ = rst ? 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 : \aes_top_0.uaes_ctr_nxt ;
  assign _0136_ = \aes_top_0.aes_reg_key0_i.en ? \aes_top_0.aes_key0_dataout : 8'b00000000;
  assign _0137_ = \aes_top_0.aes_reg_ctr_i.en ? \aes_top_0.aes_ctr_dataout : _0136_;
  assign _0138_ = \aes_top_0.aes_reg_oplen_i.en ? \aes_top_0.aes_len_dataout : _0137_;
  assign _0139_ = \aes_top_0.aes_reg_opaddr_i.en ? \aes_top_0.aes_addr_dataout : _0138_;
  logic [7:0] fangyuan0;
  assign fangyuan0 = { 6'b000000, \aes_top_0.aes_reg_state };
  assign \aes_top_0.data_out = \aes_top_0.sel_reg_state ? fangyuan0 : _0139_;
  assign _0094_[15:0] = _0115_ ? _0088_ : \aes_top_0.operated_bytes_count ;
  assign \aes_top_0.operated_bytes_count_next = \aes_top_0.reset_byte_counter ? 16'b0000000000000000 : _0094_[15:0];
  assign _0095_[15:0] = \aes_top_0.more_blocks ? _0089_ : \aes_top_0.block_counter ;
  assign \aes_top_0.block_counter_next = \aes_top_0.reset_byte_counter ? 16'b0000000000000000 : _0095_[15:0];
  assign _0096_[3:0] = \aes_top_0.xram_ack ? _0090_ : \aes_top_0.byte_counter ;
  assign \aes_top_0.byte_counter_next = \aes_top_0.reset_byte_counter ? 4'b0000 : _0096_[3:0];
  assign \aes_top_0.aes_reg_state_next_read_data = \aes_top_0.last_byte_acked ? 2'b10 : 2'b01;
  assign _0140_ = \aes_top_0.last_byte_acked ? 2'b00 : 2'b11;
  assign \aes_top_0.aes_reg_state_next_write_data = _0116_ ? 2'b01 : _0140_;
  assign _0141_ = \addr_fifo.wr ? \aes_top_0.aes_reg_state_next_write_data : 2'b00;
  logic [1:0] fangyuan1;
  assign fangyuan1 = { 1'b1, \aes_top_0.aes_time_enough };
  assign _0142_ = \aes_top_0.aes_state_operate ? fangyuan1 : _0141_;
  assign _0143_ = \aes_top_0.aes_state_read_data ? \aes_top_0.aes_reg_state_next_read_data : _0142_;
  logic [1:0] fangyuan2;
  assign fangyuan2 = { 1'b0, \aes_top_0.reset_byte_counter };
  assign \aes_top_0.aes_reg_state_next = \aes_top_0.aes_state_idle ? fangyuan2 : _0143_;
  assign \aes_top_0.mem_data_buf_next [7:0] = _0117_ ? xram_data_in : \aes_top_0.mem_data_buf [7:0];
  assign \aes_top_0.mem_data_buf_next [15:8] = _0118_ ? xram_data_in : \aes_top_0.mem_data_buf [15:8];
  assign \aes_top_0.mem_data_buf_next [23:16] = _0119_ ? xram_data_in : \aes_top_0.mem_data_buf [23:16];
  assign \aes_top_0.mem_data_buf_next [31:24] = _0120_ ? xram_data_in : \aes_top_0.mem_data_buf [31:24];
  assign \aes_top_0.mem_data_buf_next [39:32] = _0121_ ? xram_data_in : \aes_top_0.mem_data_buf [39:32];
  assign \aes_top_0.mem_data_buf_next [47:40] = _0122_ ? xram_data_in : \aes_top_0.mem_data_buf [47:40];
  assign \aes_top_0.mem_data_buf_next [55:48] = _0123_ ? xram_data_in : \aes_top_0.mem_data_buf [55:48];
  assign \aes_top_0.mem_data_buf_next [63:56] = _0124_ ? xram_data_in : \aes_top_0.mem_data_buf [63:56];
  assign \aes_top_0.mem_data_buf_next [71:64] = _0125_ ? xram_data_in : \aes_top_0.mem_data_buf [71:64];
  assign \aes_top_0.mem_data_buf_next [79:72] = _0126_ ? xram_data_in : \aes_top_0.mem_data_buf [79:72];
  assign \aes_top_0.mem_data_buf_next [87:80] = _0127_ ? xram_data_in : \aes_top_0.mem_data_buf [87:80];
  assign \aes_top_0.mem_data_buf_next [95:88] = _0128_ ? xram_data_in : \aes_top_0.mem_data_buf [95:88];
  assign \aes_top_0.mem_data_buf_next [103:96] = _0129_ ? xram_data_in : \aes_top_0.mem_data_buf [103:96];
  assign \aes_top_0.mem_data_buf_next [111:104] = _0130_ ? xram_data_in : \aes_top_0.mem_data_buf [111:104];
  assign \aes_top_0.mem_data_buf_next [119:112] = _0131_ ? xram_data_in : \aes_top_0.mem_data_buf [119:112];
  assign \aes_top_0.mem_data_buf_next [127:120] = \aes_top_0.last_byte_acked ? xram_data_in : \aes_top_0.mem_data_buf [127:120];
  assign _0144_ = \aes_top_0.more_blocks ? _0092_ : \aes_top_0.uaes_ctr ;
  assign \aes_top_0.uaes_ctr_nxt = \aes_top_0.reset_byte_counter ? \aes_top_0.aes_reg_ctr_i.reg_out : _0144_;
  assign _0145_ = _0135_ ? _0093_ : \aes_top_0.aes_time_counter ;
  assign \aes_top_0.aes_time_counter_next = _0132_ ? 5'b00000 : _0145_;
  assign \aes_top_0.encrypted_data_buf_next = \aes_top_0.aes_state_operate ? \aes_top_0.encrypted_data : \aes_top_0.encrypted_data_buf ;
  assign _0146_ = _0112_ ? \aes_top_0.encrypted_data_buf [119:112] : \aes_top_0.encrypted_data_buf [127:120];
  assign _0147_ = _0111_ ? \aes_top_0.encrypted_data_buf [111:104] : _0146_;
  assign _0148_ = _0110_ ? \aes_top_0.encrypted_data_buf [103:96] : _0147_;
  assign _0149_ = _0109_ ? \aes_top_0.encrypted_data_buf [95:88] : _0148_;
  assign _0150_ = _0108_ ? \aes_top_0.encrypted_data_buf [87:80] : _0149_;
  assign _0151_ = _0107_ ? \aes_top_0.encrypted_data_buf [79:72] : _0150_;
  assign _0152_ = _0106_ ? \aes_top_0.encrypted_data_buf [71:64] : _0151_;
  assign _0153_ = _0105_ ? \aes_top_0.encrypted_data_buf [63:56] : _0152_;
  assign _0154_ = _0104_ ? \aes_top_0.encrypted_data_buf [55:48] : _0153_;
  assign _0155_ = _0103_ ? \aes_top_0.encrypted_data_buf [47:40] : _0154_;
  assign _0156_ = _0102_ ? \aes_top_0.encrypted_data_buf [39:32] : _0155_;
  assign _0157_ = _0101_ ? \aes_top_0.encrypted_data_buf [31:24] : _0156_;
  assign _0158_ = _0100_ ? \aes_top_0.encrypted_data_buf [23:16] : _0157_;
  assign _0159_ = _0099_ ? \aes_top_0.encrypted_data_buf [15:8] : _0158_;
  assign \aes_top_0.xram_data_out = _0098_ ? \aes_top_0.encrypted_data_buf [7:0] : _0159_;
  assign \aes_top_0.encrypted_data = \aes_top_0.aes_out ^ \aes_top_0.mem_data_buf ;
  assign _0161_ = ! addr[3:0];
  assign _0162_ = addr[3:0] == 1'b1;
  assign _0163_ = addr[3:0] == 2'b10;
  assign _0164_ = addr[3:0] == 2'b11;
  assign _0165_ = addr[3:0] == 3'b100;
  assign _0166_ = addr[3:0] == 3'b101;
  assign _0167_ = addr[3:0] == 3'b110;
  assign _0168_ = addr[3:0] == 3'b111;
  assign _0169_ = addr[3:0] == 4'b1000;
  assign _0170_ = addr[3:0] == 4'b1001;
  assign _0171_ = addr[3:0] == 4'b1010;
  assign _0172_ = addr[3:0] == 4'b1011;
  assign _0173_ = addr[3:0] == 4'b1100;
  assign _0174_ = addr[3:0] == 4'b1101;
  assign _0175_ = addr[3:0] == 4'b1110;
  assign _0176_ = addr[3:0] == 4'b1111;
  assign _0177_ = \aes_top_0.aes_reg_ctr_i.en && \aes_top_0.aes_reg_ctr_i.wr ;
  assign \aes_top_0.aes_reg_ctr_i.wr0 = _0177_ && _0161_;
  assign \aes_top_0.aes_reg_ctr_i.wr1 = _0177_ && _0162_;
  assign \aes_top_0.aes_reg_ctr_i.wr2 = _0177_ && _0163_;
  assign \aes_top_0.aes_reg_ctr_i.wr3 = _0177_ && _0164_;
  assign \aes_top_0.aes_reg_ctr_i.wr4 = _0177_ && _0165_;
  assign \aes_top_0.aes_reg_ctr_i.wr5 = _0177_ && _0166_;
  assign \aes_top_0.aes_reg_ctr_i.wr6 = _0177_ && _0167_;
  assign \aes_top_0.aes_reg_ctr_i.wr7 = _0177_ && _0168_;
  assign \aes_top_0.aes_reg_ctr_i.wr8 = _0177_ && _0169_;
  assign \aes_top_0.aes_reg_ctr_i.wr9 = _0177_ && _0170_;
  assign \aes_top_0.aes_reg_ctr_i.wr10 = _0177_ && _0171_;
  assign \aes_top_0.aes_reg_ctr_i.wr11 = _0177_ && _0172_;
  assign \aes_top_0.aes_reg_ctr_i.wr12 = _0177_ && _0173_;
  assign \aes_top_0.aes_reg_ctr_i.wr13 = _0177_ && _0174_;
  assign \aes_top_0.aes_reg_ctr_i.wr14 = _0177_ && _0175_;
  assign \aes_top_0.aes_reg_ctr_i.wr15 = _0177_ && _0176_;
  always @(posedge clk)
      \aes_top_0.aes_reg_ctr_i.reg_out <= _0160_;
  assign _0160_[127:120] = rst ? 8'b00000000 : \aes_top_0.aes_reg_ctr_i.reg15_next ;
  assign _0160_[119:112] = rst ? 8'b00000000 : \aes_top_0.aes_reg_ctr_i.reg14_next ;
  assign _0160_[111:104] = rst ? 8'b00000000 : \aes_top_0.aes_reg_ctr_i.reg13_next ;
  assign _0160_[103:96] = rst ? 8'b00000000 : \aes_top_0.aes_reg_ctr_i.reg12_next ;
  assign _0160_[95:88] = rst ? 8'b00000000 : \aes_top_0.aes_reg_ctr_i.reg11_next ;
  assign _0160_[87:80] = rst ? 8'b00000000 : \aes_top_0.aes_reg_ctr_i.reg10_next ;
  assign _0160_[79:72] = rst ? 8'b00000000 : \aes_top_0.aes_reg_ctr_i.reg9_next ;
  assign _0160_[71:64] = rst ? 8'b00000000 : \aes_top_0.aes_reg_ctr_i.reg8_next ;
  assign _0160_[63:56] = rst ? 8'b00000000 : \aes_top_0.aes_reg_ctr_i.reg7_next ;
  assign _0160_[55:48] = rst ? 8'b00000000 : \aes_top_0.aes_reg_ctr_i.reg6_next ;
  assign _0160_[47:40] = rst ? 8'b00000000 : \aes_top_0.aes_reg_ctr_i.reg5_next ;
  assign _0160_[39:32] = rst ? 8'b00000000 : \aes_top_0.aes_reg_ctr_i.reg4_next ;
  assign _0160_[31:24] = rst ? 8'b00000000 : \aes_top_0.aes_reg_ctr_i.reg3_next ;
  assign _0160_[23:16] = rst ? 8'b00000000 : \aes_top_0.aes_reg_ctr_i.reg2_next ;
  assign _0160_[15:8] = rst ? 8'b00000000 : \aes_top_0.aes_reg_ctr_i.reg1_next ;
  assign _0160_[7:0] = rst ? 8'b00000000 : \aes_top_0.aes_reg_ctr_i.reg0_next ;
  assign \aes_top_0.aes_reg_ctr_i.reg0_next = \aes_top_0.aes_reg_ctr_i.wr0 ? data_in : \aes_top_0.aes_reg_ctr_i.reg_out [7:0];
  assign \aes_top_0.aes_reg_ctr_i.reg1_next = \aes_top_0.aes_reg_ctr_i.wr1 ? data_in : \aes_top_0.aes_reg_ctr_i.reg_out [15:8];
  assign \aes_top_0.aes_reg_ctr_i.reg2_next = \aes_top_0.aes_reg_ctr_i.wr2 ? data_in : \aes_top_0.aes_reg_ctr_i.reg_out [23:16];
  assign \aes_top_0.aes_reg_ctr_i.reg3_next = \aes_top_0.aes_reg_ctr_i.wr3 ? data_in : \aes_top_0.aes_reg_ctr_i.reg_out [31:24];
  assign \aes_top_0.aes_reg_ctr_i.reg4_next = \aes_top_0.aes_reg_ctr_i.wr4 ? data_in : \aes_top_0.aes_reg_ctr_i.reg_out [39:32];
  assign \aes_top_0.aes_reg_ctr_i.reg5_next = \aes_top_0.aes_reg_ctr_i.wr5 ? data_in : \aes_top_0.aes_reg_ctr_i.reg_out [47:40];
  assign \aes_top_0.aes_reg_ctr_i.reg6_next = \aes_top_0.aes_reg_ctr_i.wr6 ? data_in : \aes_top_0.aes_reg_ctr_i.reg_out [55:48];
  assign \aes_top_0.aes_reg_ctr_i.reg7_next = \aes_top_0.aes_reg_ctr_i.wr7 ? data_in : \aes_top_0.aes_reg_ctr_i.reg_out [63:56];
  assign \aes_top_0.aes_reg_ctr_i.reg8_next = \aes_top_0.aes_reg_ctr_i.wr8 ? data_in : \aes_top_0.aes_reg_ctr_i.reg_out [71:64];
  assign \aes_top_0.aes_reg_ctr_i.reg9_next = \aes_top_0.aes_reg_ctr_i.wr9 ? data_in : \aes_top_0.aes_reg_ctr_i.reg_out [79:72];
  assign \aes_top_0.aes_reg_ctr_i.reg10_next = \aes_top_0.aes_reg_ctr_i.wr10 ? data_in : \aes_top_0.aes_reg_ctr_i.reg_out [87:80];
  assign \aes_top_0.aes_reg_ctr_i.reg11_next = \aes_top_0.aes_reg_ctr_i.wr11 ? data_in : \aes_top_0.aes_reg_ctr_i.reg_out [95:88];
  assign \aes_top_0.aes_reg_ctr_i.reg12_next = \aes_top_0.aes_reg_ctr_i.wr12 ? data_in : \aes_top_0.aes_reg_ctr_i.reg_out [103:96];
  assign \aes_top_0.aes_reg_ctr_i.reg13_next = \aes_top_0.aes_reg_ctr_i.wr13 ? data_in : \aes_top_0.aes_reg_ctr_i.reg_out [111:104];
  assign \aes_top_0.aes_reg_ctr_i.reg14_next = \aes_top_0.aes_reg_ctr_i.wr14 ? data_in : \aes_top_0.aes_reg_ctr_i.reg_out [119:112];
  assign \aes_top_0.aes_reg_ctr_i.reg15_next = \aes_top_0.aes_reg_ctr_i.wr15 ? data_in : \aes_top_0.aes_reg_ctr_i.reg_out [127:120];
  assign _0178_ = _0175_ ? \aes_top_0.aes_reg_ctr_i.reg_out [119:112] : \aes_top_0.aes_reg_ctr_i.reg_out [127:120];
  assign _0179_ = _0174_ ? \aes_top_0.aes_reg_ctr_i.reg_out [111:104] : _0178_;
  assign _0180_ = _0173_ ? \aes_top_0.aes_reg_ctr_i.reg_out [103:96] : _0179_;
  assign _0181_ = _0172_ ? \aes_top_0.aes_reg_ctr_i.reg_out [95:88] : _0180_;
  assign _0182_ = _0171_ ? \aes_top_0.aes_reg_ctr_i.reg_out [87:80] : _0181_;
  assign _0183_ = _0170_ ? \aes_top_0.aes_reg_ctr_i.reg_out [79:72] : _0182_;
  assign _0184_ = _0169_ ? \aes_top_0.aes_reg_ctr_i.reg_out [71:64] : _0183_;
  assign _0185_ = _0168_ ? \aes_top_0.aes_reg_ctr_i.reg_out [63:56] : _0184_;
  assign _0186_ = _0167_ ? \aes_top_0.aes_reg_ctr_i.reg_out [55:48] : _0185_;
  assign _0187_ = _0166_ ? \aes_top_0.aes_reg_ctr_i.reg_out [47:40] : _0186_;
  assign _0188_ = _0165_ ? \aes_top_0.aes_reg_ctr_i.reg_out [39:32] : _0187_;
  assign _0189_ = _0164_ ? \aes_top_0.aes_reg_ctr_i.reg_out [31:24] : _0188_;
  assign _0190_ = _0163_ ? \aes_top_0.aes_reg_ctr_i.reg_out [23:16] : _0189_;
  assign _0191_ = _0162_ ? \aes_top_0.aes_reg_ctr_i.reg_out [15:8] : _0190_;
  assign \aes_top_0.aes_ctr_dataout = _0161_ ? \aes_top_0.aes_reg_ctr_i.reg_out [7:0] : _0191_;
  assign _0193_ = \aes_top_0.aes_reg_key0_i.en && \aes_top_0.aes_reg_key0_i.wr ;
  assign \aes_top_0.aes_reg_key0_i.wr0 = _0193_ && _0161_;
  assign \aes_top_0.aes_reg_key0_i.wr1 = _0193_ && _0162_;
  assign \aes_top_0.aes_reg_key0_i.wr2 = _0193_ && _0163_;
  assign \aes_top_0.aes_reg_key0_i.wr3 = _0193_ && _0164_;
  assign \aes_top_0.aes_reg_key0_i.wr4 = _0193_ && _0165_;
  assign \aes_top_0.aes_reg_key0_i.wr5 = _0193_ && _0166_;
  assign \aes_top_0.aes_reg_key0_i.wr6 = _0193_ && _0167_;
  assign \aes_top_0.aes_reg_key0_i.wr7 = _0193_ && _0168_;
  assign \aes_top_0.aes_reg_key0_i.wr8 = _0193_ && _0169_;
  assign \aes_top_0.aes_reg_key0_i.wr9 = _0193_ && _0170_;
  assign \aes_top_0.aes_reg_key0_i.wr10 = _0193_ && _0171_;
  assign \aes_top_0.aes_reg_key0_i.wr11 = _0193_ && _0172_;
  assign \aes_top_0.aes_reg_key0_i.wr12 = _0193_ && _0173_;
  assign \aes_top_0.aes_reg_key0_i.wr13 = _0193_ && _0174_;
  assign \aes_top_0.aes_reg_key0_i.wr14 = _0193_ && _0175_;
  assign \aes_top_0.aes_reg_key0_i.wr15 = _0193_ && _0176_;
  always @(posedge clk)
      \aes_top_0.aes_reg_key0_i.reg_out <= _0192_;
  assign _0192_[127:120] = rst ? 8'b00000000 : \aes_top_0.aes_reg_key0_i.reg15_next ;
  assign _0192_[119:112] = rst ? 8'b00000000 : \aes_top_0.aes_reg_key0_i.reg14_next ;
  assign _0192_[111:104] = rst ? 8'b00000000 : \aes_top_0.aes_reg_key0_i.reg13_next ;
  assign _0192_[103:96] = rst ? 8'b00000000 : \aes_top_0.aes_reg_key0_i.reg12_next ;
  assign _0192_[95:88] = rst ? 8'b00000000 : \aes_top_0.aes_reg_key0_i.reg11_next ;
  assign _0192_[87:80] = rst ? 8'b00000000 : \aes_top_0.aes_reg_key0_i.reg10_next ;
  assign _0192_[79:72] = rst ? 8'b00000000 : \aes_top_0.aes_reg_key0_i.reg9_next ;
  assign _0192_[71:64] = rst ? 8'b00000000 : \aes_top_0.aes_reg_key0_i.reg8_next ;
  assign _0192_[63:56] = rst ? 8'b00000000 : \aes_top_0.aes_reg_key0_i.reg7_next ;
  assign _0192_[55:48] = rst ? 8'b00000000 : \aes_top_0.aes_reg_key0_i.reg6_next ;
  assign _0192_[47:40] = rst ? 8'b00000000 : \aes_top_0.aes_reg_key0_i.reg5_next ;
  assign _0192_[39:32] = rst ? 8'b00000000 : \aes_top_0.aes_reg_key0_i.reg4_next ;
  assign _0192_[31:24] = rst ? 8'b00000000 : \aes_top_0.aes_reg_key0_i.reg3_next ;
  assign _0192_[23:16] = rst ? 8'b00000000 : \aes_top_0.aes_reg_key0_i.reg2_next ;
  assign _0192_[15:8] = rst ? 8'b00000000 : \aes_top_0.aes_reg_key0_i.reg1_next ;
  assign _0192_[7:0] = rst ? 8'b00000000 : \aes_top_0.aes_reg_key0_i.reg0_next ;
  assign \aes_top_0.aes_reg_key0_i.reg0_next = \aes_top_0.aes_reg_key0_i.wr0 ? data_in : \aes_top_0.aes_reg_key0_i.reg_out [7:0];
  assign \aes_top_0.aes_reg_key0_i.reg1_next = \aes_top_0.aes_reg_key0_i.wr1 ? data_in : \aes_top_0.aes_reg_key0_i.reg_out [15:8];
  assign \aes_top_0.aes_reg_key0_i.reg2_next = \aes_top_0.aes_reg_key0_i.wr2 ? data_in : \aes_top_0.aes_reg_key0_i.reg_out [23:16];
  assign \aes_top_0.aes_reg_key0_i.reg3_next = \aes_top_0.aes_reg_key0_i.wr3 ? data_in : \aes_top_0.aes_reg_key0_i.reg_out [31:24];
  assign \aes_top_0.aes_reg_key0_i.reg4_next = \aes_top_0.aes_reg_key0_i.wr4 ? data_in : \aes_top_0.aes_reg_key0_i.reg_out [39:32];
  assign \aes_top_0.aes_reg_key0_i.reg5_next = \aes_top_0.aes_reg_key0_i.wr5 ? data_in : \aes_top_0.aes_reg_key0_i.reg_out [47:40];
  assign \aes_top_0.aes_reg_key0_i.reg6_next = \aes_top_0.aes_reg_key0_i.wr6 ? data_in : \aes_top_0.aes_reg_key0_i.reg_out [55:48];
  assign \aes_top_0.aes_reg_key0_i.reg7_next = \aes_top_0.aes_reg_key0_i.wr7 ? data_in : \aes_top_0.aes_reg_key0_i.reg_out [63:56];
  assign \aes_top_0.aes_reg_key0_i.reg8_next = \aes_top_0.aes_reg_key0_i.wr8 ? data_in : \aes_top_0.aes_reg_key0_i.reg_out [71:64];
  assign \aes_top_0.aes_reg_key0_i.reg9_next = \aes_top_0.aes_reg_key0_i.wr9 ? data_in : \aes_top_0.aes_reg_key0_i.reg_out [79:72];
  assign \aes_top_0.aes_reg_key0_i.reg10_next = \aes_top_0.aes_reg_key0_i.wr10 ? data_in : \aes_top_0.aes_reg_key0_i.reg_out [87:80];
  assign \aes_top_0.aes_reg_key0_i.reg11_next = \aes_top_0.aes_reg_key0_i.wr11 ? data_in : \aes_top_0.aes_reg_key0_i.reg_out [95:88];
  assign \aes_top_0.aes_reg_key0_i.reg12_next = \aes_top_0.aes_reg_key0_i.wr12 ? data_in : \aes_top_0.aes_reg_key0_i.reg_out [103:96];
  assign \aes_top_0.aes_reg_key0_i.reg13_next = \aes_top_0.aes_reg_key0_i.wr13 ? data_in : \aes_top_0.aes_reg_key0_i.reg_out [111:104];
  assign \aes_top_0.aes_reg_key0_i.reg14_next = \aes_top_0.aes_reg_key0_i.wr14 ? data_in : \aes_top_0.aes_reg_key0_i.reg_out [119:112];
  assign \aes_top_0.aes_reg_key0_i.reg15_next = \aes_top_0.aes_reg_key0_i.wr15 ? data_in : \aes_top_0.aes_reg_key0_i.reg_out [127:120];
  assign _0194_ = _0175_ ? \aes_top_0.aes_reg_key0_i.reg_out [119:112] : \aes_top_0.aes_reg_key0_i.reg_out [127:120];
  assign _0195_ = _0174_ ? \aes_top_0.aes_reg_key0_i.reg_out [111:104] : _0194_;
  assign _0196_ = _0173_ ? \aes_top_0.aes_reg_key0_i.reg_out [103:96] : _0195_;
  assign _0197_ = _0172_ ? \aes_top_0.aes_reg_key0_i.reg_out [95:88] : _0196_;
  assign _0198_ = _0171_ ? \aes_top_0.aes_reg_key0_i.reg_out [87:80] : _0197_;
  assign _0199_ = _0170_ ? \aes_top_0.aes_reg_key0_i.reg_out [79:72] : _0198_;
  assign _0200_ = _0169_ ? \aes_top_0.aes_reg_key0_i.reg_out [71:64] : _0199_;
  assign _0201_ = _0168_ ? \aes_top_0.aes_reg_key0_i.reg_out [63:56] : _0200_;
  assign _0202_ = _0167_ ? \aes_top_0.aes_reg_key0_i.reg_out [55:48] : _0201_;
  assign _0203_ = _0166_ ? \aes_top_0.aes_reg_key0_i.reg_out [47:40] : _0202_;
  assign _0204_ = _0165_ ? \aes_top_0.aes_reg_key0_i.reg_out [39:32] : _0203_;
  assign _0205_ = _0164_ ? \aes_top_0.aes_reg_key0_i.reg_out [31:24] : _0204_;
  assign _0206_ = _0163_ ? \aes_top_0.aes_reg_key0_i.reg_out [23:16] : _0205_;
  assign _0207_ = _0162_ ? \aes_top_0.aes_reg_key0_i.reg_out [15:8] : _0206_;
  assign \aes_top_0.aes_key0_dataout = _0161_ ? \aes_top_0.aes_reg_key0_i.reg_out [7:0] : _0207_;
  assign _0209_ = ~ addr[0];
  assign _0210_ = \aes_top_0.aes_reg_opaddr_i.en && \aes_top_0.aes_reg_opaddr_i.wr ;
  assign \aes_top_0.aes_reg_opaddr_i.wr0 = _0210_ && _0209_;
  assign \aes_top_0.aes_reg_opaddr_i.wr1 = _0210_ && addr[0];
  always @(posedge clk)
      \aes_top_0.aes_reg_opaddr_i.reg_out <= _0208_;
  assign _0208_[15:8] = rst ? 8'b00000000 : \aes_top_0.aes_reg_opaddr_i.reg1_next ;
  assign _0208_[7:0] = rst ? 8'b00000000 : \aes_top_0.aes_reg_opaddr_i.reg0_next ;
  assign \aes_top_0.aes_reg_opaddr_i.reg0_next = \aes_top_0.aes_reg_opaddr_i.wr0 ? data_in : \aes_top_0.aes_reg_opaddr_i.reg_out [7:0];
  assign \aes_top_0.aes_reg_opaddr_i.reg1_next = \aes_top_0.aes_reg_opaddr_i.wr1 ? data_in : \aes_top_0.aes_reg_opaddr_i.reg_out [15:8];
  assign \aes_top_0.aes_addr_dataout = addr[0] ? \aes_top_0.aes_reg_opaddr_i.reg_out [15:8] : \aes_top_0.aes_reg_opaddr_i.reg_out [7:0];
  assign _0212_ = \aes_top_0.aes_reg_oplen_i.en && \aes_top_0.aes_reg_oplen_i.wr ;
  assign \aes_top_0.aes_reg_oplen_i.wr0 = _0212_ && _0209_;
  assign \aes_top_0.aes_reg_oplen_i.wr1 = _0212_ && addr[0];
  always @(posedge clk)
      \aes_top_0.aes_reg_oplen_i.reg_out <= _0211_;
  assign _0211_[15:8] = rst ? 8'b00000000 : \aes_top_0.aes_reg_oplen_i.reg1_next ;
  assign _0211_[7:0] = rst ? 8'b00000000 : \aes_top_0.aes_reg_oplen_i.reg0_next ;
  assign \aes_top_0.aes_reg_oplen_i.reg0_next = \aes_top_0.aes_reg_oplen_i.wr0 ? data_in : \aes_top_0.aes_reg_oplen_i.reg_out [7:0];
  assign \aes_top_0.aes_reg_oplen_i.reg1_next = \aes_top_0.aes_reg_oplen_i.wr1 ? data_in : \aes_top_0.aes_reg_oplen_i.reg_out [15:8];
  assign \aes_top_0.aes_len_dataout = addr[0] ? \aes_top_0.aes_reg_oplen_i.reg_out [15:8] : \aes_top_0.aes_reg_oplen_i.reg_out [7:0];
  always @(posedge clk)
      \data_fifo.r1 <= _0224_;
  always @(posedge clk)
      \data_fifo.r2 <= _0235_;
  always @(posedge clk)
      \data_fifo.r3 <= _0246_;
  always @(posedge clk)
      \data_fifo.r4 <= _0247_;
  always @(posedge clk)
      \data_fifo.r5 <= _0248_;
  always @(posedge clk)
      \data_fifo.r6 <= _0249_;
  always @(posedge clk)
      \data_fifo.r7 <= _0250_;
  always @(posedge clk)
      \data_fifo.r8 <= _0251_;
  always @(posedge clk)
      \data_fifo.r9 <= _0252_;
  always @(posedge clk)
      \data_fifo.r0 <= _0213_;
  always @(posedge clk)
      \data_fifo.r10 <= _0214_;
  always @(posedge clk)
      \data_fifo.r11 <= _0215_;
  always @(posedge clk)
      \data_fifo.r12 <= _0216_;
  always @(posedge clk)
      \data_fifo.r13 <= _0217_;
  always @(posedge clk)
      \data_fifo.r14 <= _0218_;
  always @(posedge clk)
      \data_fifo.r15 <= _0219_;
  always @(posedge clk)
      \data_fifo.r16 <= _0220_;
  always @(posedge clk)
      \data_fifo.r17 <= _0221_;
  always @(posedge clk)
      \data_fifo.r18 <= _0222_;
  always @(posedge clk)
      \data_fifo.r19 <= _0223_;
  always @(posedge clk)
      \data_fifo.r20 <= _0225_;
  always @(posedge clk)
      \data_fifo.r21 <= _0226_;
  always @(posedge clk)
      \data_fifo.r22 <= _0227_;
  always @(posedge clk)
      \data_fifo.r23 <= _0228_;
  always @(posedge clk)
      \data_fifo.r24 <= _0229_;
  always @(posedge clk)
      \data_fifo.r25 <= _0230_;
  always @(posedge clk)
      \data_fifo.r26 <= _0231_;
  always @(posedge clk)
      \data_fifo.r27 <= _0232_;
  always @(posedge clk)
      \data_fifo.r28 <= _0233_;
  always @(posedge clk)
      \data_fifo.r29 <= _0234_;
  always @(posedge clk)
      \data_fifo.r30 <= _0236_;
  always @(posedge clk)
      \data_fifo.r31 <= _0237_;
  always @(posedge clk)
      \data_fifo.r32 <= _0238_;
  always @(posedge clk)
      \data_fifo.r33 <= _0239_;
  always @(posedge clk)
      \data_fifo.r34 <= _0240_;
  always @(posedge clk)
      \data_fifo.r35 <= _0241_;
  always @(posedge clk)
      \data_fifo.r36 <= _0242_;
  always @(posedge clk)
      \data_fifo.r37 <= _0243_;
  always @(posedge clk)
      \data_fifo.r38 <= _0244_;
  always @(posedge clk)
      \data_fifo.r39 <= _0245_;
  assign _0253_ = \addr_fifo.wr ? \data_fifo.r38 : \data_fifo.r39 ;
  assign _0245_ = rst ? 8'b00000000 : _0253_;
  assign _0254_ = \addr_fifo.wr ? \data_fifo.r37 : \data_fifo.r38 ;
  assign _0244_ = rst ? 8'b00000000 : _0254_;
  assign _0255_ = \addr_fifo.wr ? \data_fifo.r36 : \data_fifo.r37 ;
  assign _0243_ = rst ? 8'b00000000 : _0255_;
  assign _0256_ = \addr_fifo.wr ? \data_fifo.r35 : \data_fifo.r36 ;
  assign _0242_ = rst ? 8'b00000000 : _0256_;
  assign _0257_ = \addr_fifo.wr ? \data_fifo.r34 : \data_fifo.r35 ;
  assign _0241_ = rst ? 8'b00000000 : _0257_;
  assign _0258_ = \addr_fifo.wr ? \data_fifo.r33 : \data_fifo.r34 ;
  assign _0240_ = rst ? 8'b00000000 : _0258_;
  assign _0259_ = \addr_fifo.wr ? \data_fifo.r32 : \data_fifo.r33 ;
  assign _0239_ = rst ? 8'b00000000 : _0259_;
  assign _0260_ = \addr_fifo.wr ? \data_fifo.r31 : \data_fifo.r32 ;
  assign _0238_ = rst ? 8'b00000000 : _0260_;
  assign _0261_ = \addr_fifo.wr ? \data_fifo.r30 : \data_fifo.r31 ;
  assign _0237_ = rst ? 8'b00000000 : _0261_;
  assign _0262_ = \addr_fifo.wr ? \data_fifo.r29 : \data_fifo.r30 ;
  assign _0236_ = rst ? 8'b00000000 : _0262_;
  assign _0263_ = \addr_fifo.wr ? \data_fifo.r28 : \data_fifo.r29 ;
  assign _0234_ = rst ? 8'b00000000 : _0263_;
  assign _0264_ = \addr_fifo.wr ? \data_fifo.r27 : \data_fifo.r28 ;
  assign _0233_ = rst ? 8'b00000000 : _0264_;
  assign _0265_ = \addr_fifo.wr ? \data_fifo.r26 : \data_fifo.r27 ;
  assign _0232_ = rst ? 8'b00000000 : _0265_;
  assign _0266_ = \addr_fifo.wr ? \data_fifo.r25 : \data_fifo.r26 ;
  assign _0231_ = rst ? 8'b00000000 : _0266_;
  assign _0267_ = \addr_fifo.wr ? \data_fifo.r24 : \data_fifo.r25 ;
  assign _0230_ = rst ? 8'b00000000 : _0267_;
  assign _0268_ = \addr_fifo.wr ? \data_fifo.r23 : \data_fifo.r24 ;
  assign _0229_ = rst ? 8'b00000000 : _0268_;
  assign _0269_ = \addr_fifo.wr ? \data_fifo.r22 : \data_fifo.r23 ;
  assign _0228_ = rst ? 8'b00000000 : _0269_;
  assign _0270_ = \addr_fifo.wr ? \data_fifo.r21 : \data_fifo.r22 ;
  assign _0227_ = rst ? 8'b00000000 : _0270_;
  assign _0271_ = \addr_fifo.wr ? \data_fifo.r20 : \data_fifo.r21 ;
  assign _0226_ = rst ? 8'b00000000 : _0271_;
  assign _0272_ = \addr_fifo.wr ? \data_fifo.r19 : \data_fifo.r20 ;
  assign _0225_ = rst ? 8'b00000000 : _0272_;
  assign _0273_ = \addr_fifo.wr ? \data_fifo.r18 : \data_fifo.r19 ;
  assign _0223_ = rst ? 8'b00000000 : _0273_;
  assign _0274_ = \addr_fifo.wr ? \data_fifo.r17 : \data_fifo.r18 ;
  assign _0222_ = rst ? 8'b00000000 : _0274_;
  assign _0275_ = \addr_fifo.wr ? \data_fifo.r16 : \data_fifo.r17 ;
  assign _0221_ = rst ? 8'b00000000 : _0275_;
  assign _0276_ = \addr_fifo.wr ? \data_fifo.r15 : \data_fifo.r16 ;
  assign _0220_ = rst ? 8'b00000000 : _0276_;
  assign _0277_ = \addr_fifo.wr ? \data_fifo.r14 : \data_fifo.r15 ;
  assign _0219_ = rst ? 8'b00000000 : _0277_;
  assign _0278_ = \addr_fifo.wr ? \data_fifo.r13 : \data_fifo.r14 ;
  assign _0218_ = rst ? 8'b00000000 : _0278_;
  assign _0279_ = \addr_fifo.wr ? \data_fifo.r12 : \data_fifo.r13 ;
  assign _0217_ = rst ? 8'b00000000 : _0279_;
  assign _0280_ = \addr_fifo.wr ? \data_fifo.r11 : \data_fifo.r12 ;
  assign _0216_ = rst ? 8'b00000000 : _0280_;
  assign _0281_ = \addr_fifo.wr ? \data_fifo.r10 : \data_fifo.r11 ;
  assign _0215_ = rst ? 8'b00000000 : _0281_;
  assign _0282_ = \addr_fifo.wr ? \data_fifo.r9 : \data_fifo.r10 ;
  assign _0214_ = rst ? 8'b00000000 : _0282_;
  assign _0283_ = \addr_fifo.wr ? \aes_top_0.xram_data_out : \data_fifo.r0 ;
  assign _0213_ = rst ? 8'b00000000 : _0283_;
  assign _0284_ = \addr_fifo.wr ? \data_fifo.r8 : \data_fifo.r9 ;
  assign _0252_ = rst ? 8'b00000000 : _0284_;
  assign _0285_ = \addr_fifo.wr ? \data_fifo.r7 : \data_fifo.r8 ;
  assign _0251_ = rst ? 8'b00000000 : _0285_;
  assign _0286_ = \addr_fifo.wr ? \data_fifo.r6 : \data_fifo.r7 ;
  assign _0250_ = rst ? 8'b00000000 : _0286_;
  assign _0287_ = \addr_fifo.wr ? \data_fifo.r5 : \data_fifo.r6 ;
  assign _0249_ = rst ? 8'b00000000 : _0287_;
  assign _0288_ = \addr_fifo.wr ? \data_fifo.r4 : \data_fifo.r5 ;
  assign _0248_ = rst ? 8'b00000000 : _0288_;
  assign _0289_ = \addr_fifo.wr ? \data_fifo.r3 : \data_fifo.r4 ;
  assign _0247_ = rst ? 8'b00000000 : _0289_;
  assign _0290_ = \addr_fifo.wr ? \data_fifo.r2 : \data_fifo.r3 ;
  assign _0246_ = rst ? 8'b00000000 : _0290_;
  assign _0291_ = \addr_fifo.wr ? \data_fifo.r1 : \data_fifo.r2 ;
  assign _0235_ = rst ? 8'b00000000 : _0291_;
  assign _0292_ = \addr_fifo.wr ? \data_fifo.r0 : \data_fifo.r1 ;
  assign _0224_ = rst ? 8'b00000000 : _0292_;
  always @(posedge clk)
      \wr_fifo.r1 <= _0304_;
  always @(posedge clk)
      \wr_fifo.r2 <= _0315_;
  always @(posedge clk)
      \wr_fifo.r3 <= _0326_;
  always @(posedge clk)
      \wr_fifo.r4 <= _0327_;
  always @(posedge clk)
      \wr_fifo.r5 <= _0328_;
  always @(posedge clk)
      \wr_fifo.r6 <= _0329_;
  always @(posedge clk)
      \wr_fifo.r7 <= _0330_;
  always @(posedge clk)
      \wr_fifo.r8 <= _0331_;
  always @(posedge clk)
      \wr_fifo.r9 <= _0332_;
  always @(posedge clk)
      \wr_fifo.r0 <= _0293_;
  always @(posedge clk)
      \wr_fifo.r10 <= _0294_;
  always @(posedge clk)
      \wr_fifo.r11 <= _0295_;
  always @(posedge clk)
      \wr_fifo.r12 <= _0296_;
  always @(posedge clk)
      \wr_fifo.r13 <= _0297_;
  always @(posedge clk)
      \wr_fifo.r14 <= _0298_;
  always @(posedge clk)
      \wr_fifo.r15 <= _0299_;
  always @(posedge clk)
      \wr_fifo.r16 <= _0300_;
  always @(posedge clk)
      \wr_fifo.r17 <= _0301_;
  always @(posedge clk)
      \wr_fifo.r18 <= _0302_;
  always @(posedge clk)
      \wr_fifo.r19 <= _0303_;
  always @(posedge clk)
      \wr_fifo.r20 <= _0305_;
  always @(posedge clk)
      \wr_fifo.r21 <= _0306_;
  always @(posedge clk)
      \wr_fifo.r22 <= _0307_;
  always @(posedge clk)
      \wr_fifo.r23 <= _0308_;
  always @(posedge clk)
      \wr_fifo.r24 <= _0309_;
  always @(posedge clk)
      \wr_fifo.r25 <= _0310_;
  always @(posedge clk)
      \wr_fifo.r26 <= _0311_;
  always @(posedge clk)
      \wr_fifo.r27 <= _0312_;
  always @(posedge clk)
      \wr_fifo.r28 <= _0313_;
  always @(posedge clk)
      \wr_fifo.r29 <= _0314_;
  always @(posedge clk)
      \wr_fifo.r30 <= _0316_;
  always @(posedge clk)
      \wr_fifo.r31 <= _0317_;
  always @(posedge clk)
      \wr_fifo.r32 <= _0318_;
  always @(posedge clk)
      \wr_fifo.r33 <= _0319_;
  always @(posedge clk)
      \wr_fifo.r34 <= _0320_;
  always @(posedge clk)
      \wr_fifo.r35 <= _0321_;
  always @(posedge clk)
      \wr_fifo.r36 <= _0322_;
  always @(posedge clk)
      \wr_fifo.r37 <= _0323_;
  always @(posedge clk)
      \wr_fifo.r38 <= _0324_;
  always @(posedge clk)
      \wr_fifo.r39 <= _0325_;
  assign _0333_ = \addr_fifo.wr ? \wr_fifo.r38 : \wr_fifo.r39 ;
  assign _0325_ = rst ? 1'b0 : _0333_;
  assign _0334_ = \addr_fifo.wr ? \wr_fifo.r37 : \wr_fifo.r38 ;
  assign _0324_ = rst ? 1'b0 : _0334_;
  assign _0335_ = \addr_fifo.wr ? \wr_fifo.r36 : \wr_fifo.r37 ;
  assign _0323_ = rst ? 1'b0 : _0335_;
  assign _0336_ = \addr_fifo.wr ? \wr_fifo.r35 : \wr_fifo.r36 ;
  assign _0322_ = rst ? 1'b0 : _0336_;
  assign _0337_ = \addr_fifo.wr ? \wr_fifo.r34 : \wr_fifo.r35 ;
  assign _0321_ = rst ? 1'b0 : _0337_;
  assign _0338_ = \addr_fifo.wr ? \wr_fifo.r33 : \wr_fifo.r34 ;
  assign _0320_ = rst ? 1'b0 : _0338_;
  assign _0339_ = \addr_fifo.wr ? \wr_fifo.r32 : \wr_fifo.r33 ;
  assign _0319_ = rst ? 1'b0 : _0339_;
  assign _0340_ = \addr_fifo.wr ? \wr_fifo.r31 : \wr_fifo.r32 ;
  assign _0318_ = rst ? 1'b0 : _0340_;
  assign _0341_ = \addr_fifo.wr ? \wr_fifo.r30 : \wr_fifo.r31 ;
  assign _0317_ = rst ? 1'b0 : _0341_;
  assign _0342_ = \addr_fifo.wr ? \wr_fifo.r29 : \wr_fifo.r30 ;
  assign _0316_ = rst ? 1'b0 : _0342_;
  assign _0343_ = \addr_fifo.wr ? \wr_fifo.r28 : \wr_fifo.r29 ;
  assign _0314_ = rst ? 1'b0 : _0343_;
  assign _0344_ = \addr_fifo.wr ? \wr_fifo.r27 : \wr_fifo.r28 ;
  assign _0313_ = rst ? 1'b0 : _0344_;
  assign _0345_ = \addr_fifo.wr ? \wr_fifo.r26 : \wr_fifo.r27 ;
  assign _0312_ = rst ? 1'b0 : _0345_;
  assign _0346_ = \addr_fifo.wr ? \wr_fifo.r25 : \wr_fifo.r26 ;
  assign _0311_ = rst ? 1'b0 : _0346_;
  assign _0347_ = \addr_fifo.wr ? \wr_fifo.r24 : \wr_fifo.r25 ;
  assign _0310_ = rst ? 1'b0 : _0347_;
  assign _0348_ = \addr_fifo.wr ? \wr_fifo.r23 : \wr_fifo.r24 ;
  assign _0309_ = rst ? 1'b0 : _0348_;
  assign _0349_ = \addr_fifo.wr ? \wr_fifo.r22 : \wr_fifo.r23 ;
  assign _0308_ = rst ? 1'b0 : _0349_;
  assign _0350_ = \addr_fifo.wr ? \wr_fifo.r21 : \wr_fifo.r22 ;
  assign _0307_ = rst ? 1'b0 : _0350_;
  assign _0351_ = \addr_fifo.wr ? \wr_fifo.r20 : \wr_fifo.r21 ;
  assign _0306_ = rst ? 1'b0 : _0351_;
  assign _0352_ = \addr_fifo.wr ? \wr_fifo.r19 : \wr_fifo.r20 ;
  assign _0305_ = rst ? 1'b0 : _0352_;
  assign _0353_ = \addr_fifo.wr ? \wr_fifo.r18 : \wr_fifo.r19 ;
  assign _0303_ = rst ? 1'b0 : _0353_;
  assign _0354_ = \addr_fifo.wr ? \wr_fifo.r17 : \wr_fifo.r18 ;
  assign _0302_ = rst ? 1'b0 : _0354_;
  assign _0355_ = \addr_fifo.wr ? \wr_fifo.r16 : \wr_fifo.r17 ;
  assign _0301_ = rst ? 1'b0 : _0355_;
  assign _0356_ = \addr_fifo.wr ? \wr_fifo.r15 : \wr_fifo.r16 ;
  assign _0300_ = rst ? 1'b0 : _0356_;
  assign _0357_ = \addr_fifo.wr ? \wr_fifo.r14 : \wr_fifo.r15 ;
  assign _0299_ = rst ? 1'b0 : _0357_;
  assign _0358_ = \addr_fifo.wr ? \wr_fifo.r13 : \wr_fifo.r14 ;
  assign _0298_ = rst ? 1'b0 : _0358_;
  assign _0359_ = \addr_fifo.wr ? \wr_fifo.r12 : \wr_fifo.r13 ;
  assign _0297_ = rst ? 1'b0 : _0359_;
  assign _0360_ = \addr_fifo.wr ? \wr_fifo.r11 : \wr_fifo.r12 ;
  assign _0296_ = rst ? 1'b0 : _0360_;
  assign _0361_ = \addr_fifo.wr ? \wr_fifo.r10 : \wr_fifo.r11 ;
  assign _0295_ = rst ? 1'b0 : _0361_;
  assign _0362_ = \addr_fifo.wr ? \wr_fifo.r9 : \wr_fifo.r10 ;
  assign _0294_ = rst ? 1'b0 : _0362_;
  assign _0363_ = \addr_fifo.wr ? 1'b1 : \wr_fifo.r0 ;
  assign _0293_ = rst ? 1'b0 : _0363_;
  assign _0364_ = \addr_fifo.wr ? \wr_fifo.r8 : \wr_fifo.r9 ;
  assign _0332_ = rst ? 1'b0 : _0364_;
  assign _0365_ = \addr_fifo.wr ? \wr_fifo.r7 : \wr_fifo.r8 ;
  assign _0331_ = rst ? 1'b0 : _0365_;
  assign _0366_ = \addr_fifo.wr ? \wr_fifo.r6 : \wr_fifo.r7 ;
  assign _0330_ = rst ? 1'b0 : _0366_;
  assign _0367_ = \addr_fifo.wr ? \wr_fifo.r5 : \wr_fifo.r6 ;
  assign _0329_ = rst ? 1'b0 : _0367_;
  assign _0368_ = \addr_fifo.wr ? \wr_fifo.r4 : \wr_fifo.r5 ;
  assign _0328_ = rst ? 1'b0 : _0368_;
  assign _0369_ = \addr_fifo.wr ? \wr_fifo.r3 : \wr_fifo.r4 ;
  assign _0327_ = rst ? 1'b0 : _0369_;
  assign _0370_ = \addr_fifo.wr ? \wr_fifo.r2 : \wr_fifo.r3 ;
  assign _0326_ = rst ? 1'b0 : _0370_;
  assign _0371_ = \addr_fifo.wr ? \wr_fifo.r1 : \wr_fifo.r2 ;
  assign _0315_ = rst ? 1'b0 : _0371_;
  assign _0372_ = \addr_fifo.wr ? \wr_fifo.r0 : \wr_fifo.r1 ;
  assign _0304_ = rst ? 1'b0 : _0372_;
  aes_128 \aes_top_0.aes_128_i (
    .clk(clk),
    .key(\aes_top_0.aes_reg_key0_i.reg_out ),
    .out(\aes_top_0.aes_out ),
    .state(\aes_top_0.uaes_ctr )
  );
  assign ack = \aes_top_0.ack ;
  assign \addr_fifo.ack = \aes_top_0.xram_ack ;
  assign \addr_fifo.clk = clk;
  assign \addr_fifo.out = \addr_fifo.r39 ;
  assign \addr_fifo.rst = rst;
  assign \addr_fifo.stb = \aes_top_0.xram_ack ;
  assign addr_fifo_out = \addr_fifo.r39 ;
  assign aes_addr = \aes_top_0.aes_reg_opaddr_i.reg_out ;
  assign aes_ctr = \aes_top_0.aes_reg_ctr_i.reg_out ;
  assign aes_key0 = \aes_top_0.aes_reg_key0_i.reg_out ;
  assign aes_len = \aes_top_0.aes_reg_oplen_i.reg_out ;
  assign aes_state = \aes_top_0.aes_reg_state ;
  assign aes_step = \aes_top_0.aes_step ;
  assign \aes_top_0.addr = addr;
  assign \aes_top_0.aes_addr = \aes_top_0.aes_reg_opaddr_i.reg_out ;
  assign \aes_top_0.aes_ctr = \aes_top_0.aes_reg_ctr_i.reg_out ;
  assign \aes_top_0.aes_curr_key = \aes_top_0.aes_reg_key0_i.reg_out ;
  assign \aes_top_0.aes_key0 = \aes_top_0.aes_reg_key0_i.reg_out ;
  assign \aes_top_0.aes_len = \aes_top_0.aes_reg_oplen_i.reg_out ;
  assign \aes_top_0.aes_reg_ctr = \aes_top_0.aes_reg_ctr_i.reg_out ;
  assign \aes_top_0.aes_reg_ctr_i.addr = addr[3:0];
  assign \aes_top_0.aes_reg_ctr_i.clk = clk;
  assign \aes_top_0.aes_reg_ctr_i.data_in = data_in;
  assign \aes_top_0.aes_reg_ctr_i.data_out = \aes_top_0.aes_ctr_dataout ;
  assign \aes_top_0.aes_reg_ctr_i.data_out_mux = \aes_top_0.aes_ctr_dataout ;
  assign \aes_top_0.aes_reg_ctr_i.rst = rst;
  assign \aes_top_0.aes_reg_key0 = \aes_top_0.aes_reg_key0_i.reg_out ;
  assign \aes_top_0.aes_reg_key0_i.addr = addr[3:0];
  assign \aes_top_0.aes_reg_key0_i.clk = clk;
  assign \aes_top_0.aes_reg_key0_i.data_in = data_in;
  assign \aes_top_0.aes_reg_key0_i.data_out = \aes_top_0.aes_key0_dataout ;
  assign \aes_top_0.aes_reg_key0_i.data_out_mux = \aes_top_0.aes_key0_dataout ;
  assign \aes_top_0.aes_reg_key0_i.rst = rst;
  assign \aes_top_0.aes_reg_opaddr = \aes_top_0.aes_reg_opaddr_i.reg_out ;
  assign \aes_top_0.aes_reg_opaddr_i.addr = addr[0];
  assign \aes_top_0.aes_reg_opaddr_i.clk = clk;
  assign \aes_top_0.aes_reg_opaddr_i.data_in = data_in;
  assign \aes_top_0.aes_reg_opaddr_i.data_out = \aes_top_0.aes_addr_dataout ;
  assign \aes_top_0.aes_reg_opaddr_i.data_out_mux = \aes_top_0.aes_addr_dataout ;
  assign \aes_top_0.aes_reg_opaddr_i.rst = rst;
  assign \aes_top_0.aes_reg_oplen = \aes_top_0.aes_reg_oplen_i.reg_out ;
  assign \aes_top_0.aes_reg_oplen_i.addr = addr[0];
  assign \aes_top_0.aes_reg_oplen_i.clk = clk;
  assign \aes_top_0.aes_reg_oplen_i.data_in = data_in;
  assign \aes_top_0.aes_reg_oplen_i.data_out = \aes_top_0.aes_len_dataout ;
  assign \aes_top_0.aes_reg_oplen_i.data_out_mux = \aes_top_0.aes_len_dataout ;
  assign \aes_top_0.aes_reg_oplen_i.rst = rst;
  assign \aes_top_0.aes_reg_state_next_idle = \aes_top_0.reset_byte_counter ;
  assign \aes_top_0.aes_reg_state_next_operate = \aes_top_0.aes_time_enough ;
  assign \aes_top_0.aes_state = \aes_top_0.aes_reg_state ;
  assign \aes_top_0.aes_state_write_data = \addr_fifo.wr ;
  assign \aes_top_0.clk = clk;
  assign \aes_top_0.data_in = data_in;
  assign \aes_top_0.incr_byte_counter = \aes_top_0.xram_ack ;
  assign \aes_top_0.rst = rst;
  assign \aes_top_0.sel_reg_addr = \aes_top_0.aes_reg_opaddr_i.en ;
  assign \aes_top_0.sel_reg_ctr = \aes_top_0.aes_reg_ctr_i.en ;
  assign \aes_top_0.sel_reg_key0 = \aes_top_0.aes_reg_key0_i.en ;
  assign \aes_top_0.sel_reg_len = \aes_top_0.aes_reg_oplen_i.en ;
  assign \aes_top_0.start_op = \aes_top_0.reset_byte_counter ;
  assign \aes_top_0.stb = stb;
  assign \aes_top_0.wr = wr;
  assign \aes_top_0.xram_addr = \addr_fifo.in ;
  assign \aes_top_0.xram_data_in = xram_data_in;
  assign \aes_top_0.xram_stb = \aes_top_0.xram_ack ;
  assign \aes_top_0.xram_wr = \addr_fifo.wr ;
  assign \data_fifo.ack = \aes_top_0.xram_ack ;
  assign \data_fifo.clk = clk;
  assign \data_fifo.in = \aes_top_0.xram_data_out ;
  assign \data_fifo.out = \data_fifo.r39 ;
  assign \data_fifo.rst = rst;
  assign \data_fifo.stb = \aes_top_0.xram_ack ;
  assign \data_fifo.wr = \addr_fifo.wr ;
  assign data_fifo_out = \data_fifo.r39 ;
  assign data_out = \aes_top_0.data_out ;
  assign \wr_fifo.ack = \aes_top_0.xram_ack ;
  assign \wr_fifo.clk = clk;
  assign \wr_fifo.in = \addr_fifo.wr ;
  assign \wr_fifo.out = \wr_fifo.r39 ;
  assign \wr_fifo.rst = rst;
  assign \wr_fifo.stb = \aes_top_0.xram_ack ;
  assign \wr_fifo.wr = \addr_fifo.wr ;
  assign wr_fifo_out = \wr_fifo.r39 ;
  assign xram_ack = \aes_top_0.xram_ack ;
  assign xram_addr = \addr_fifo.in ;
  assign xram_data_out = \aes_top_0.xram_data_out ;
  assign xram_stb = \aes_top_0.xram_ack ;
  assign xram_wr = \addr_fifo.wr ;
endmodule
