module NV_NVDLA_CSC_dl(nvdla_core_clk, nvdla_core_rstn, sg2dl_pvld, sg2dl_pd, sc_state, sg2dl_reuse_rls, sc2cdma_dat_pending_req, cdma2sc_dat_updt, cdma2sc_dat_entries, cdma2sc_dat_slices, sc2cdma_dat_updt, sc2cdma_dat_entries, sc2cdma_dat_slices, sc2buf_dat_rd_en, sc2buf_dat_rd_addr, sc2buf_dat_rd_valid, sc2buf_dat_rd_data, sc2mac_dat_a_pvld, sc2mac_dat_a_mask, sc2mac_dat_a_data0, sc2mac_dat_a_data1, sc2mac_dat_a_data2, sc2mac_dat_a_data3, sc2mac_dat_a_data4, sc2mac_dat_a_data5, sc2mac_dat_a_data6, sc2mac_dat_a_data7, sc2mac_dat_a_data8, sc2mac_dat_a_data9, sc2mac_dat_a_data10, sc2mac_dat_a_data11, sc2mac_dat_a_data12, sc2mac_dat_a_data13, sc2mac_dat_a_data14, sc2mac_dat_a_data15, sc2mac_dat_a_data16, sc2mac_dat_a_data17, sc2mac_dat_a_data18, sc2mac_dat_a_data19, sc2mac_dat_a_data20, sc2mac_dat_a_data21, sc2mac_dat_a_data22, sc2mac_dat_a_data23, sc2mac_dat_a_data24, sc2mac_dat_a_data25, sc2mac_dat_a_data26, sc2mac_dat_a_data27, sc2mac_dat_a_data28, sc2mac_dat_a_data29, sc2mac_dat_a_data30, sc2mac_dat_a_data31, sc2mac_dat_a_data32, sc2mac_dat_a_data33, sc2mac_dat_a_data34, sc2mac_dat_a_data35, sc2mac_dat_a_data36, sc2mac_dat_a_data37, sc2mac_dat_a_data38, sc2mac_dat_a_data39, sc2mac_dat_a_data40, sc2mac_dat_a_data41, sc2mac_dat_a_data42, sc2mac_dat_a_data43, sc2mac_dat_a_data44, sc2mac_dat_a_data45, sc2mac_dat_a_data46, sc2mac_dat_a_data47, sc2mac_dat_a_data48, sc2mac_dat_a_data49, sc2mac_dat_a_data50, sc2mac_dat_a_data51, sc2mac_dat_a_data52, sc2mac_dat_a_data53, sc2mac_dat_a_data54, sc2mac_dat_a_data55, sc2mac_dat_a_data56, sc2mac_dat_a_data57, sc2mac_dat_a_data58, sc2mac_dat_a_data59, sc2mac_dat_a_data60, sc2mac_dat_a_data61, sc2mac_dat_a_data62, sc2mac_dat_a_data63, sc2mac_dat_a_data64, sc2mac_dat_a_data65, sc2mac_dat_a_data66, sc2mac_dat_a_data67, sc2mac_dat_a_data68, sc2mac_dat_a_data69, sc2mac_dat_a_data70, sc2mac_dat_a_data71, sc2mac_dat_a_data72, sc2mac_dat_a_data73, sc2mac_dat_a_data74, sc2mac_dat_a_data75, sc2mac_dat_a_data76, sc2mac_dat_a_data77, sc2mac_dat_a_data78, sc2mac_dat_a_data79, sc2mac_dat_a_data80, sc2mac_dat_a_data81, sc2mac_dat_a_data82, sc2mac_dat_a_data83, sc2mac_dat_a_data84, sc2mac_dat_a_data85, sc2mac_dat_a_data86, sc2mac_dat_a_data87, sc2mac_dat_a_data88, sc2mac_dat_a_data89, sc2mac_dat_a_data90, sc2mac_dat_a_data91, sc2mac_dat_a_data92, sc2mac_dat_a_data93, sc2mac_dat_a_data94, sc2mac_dat_a_data95, sc2mac_dat_a_data96, sc2mac_dat_a_data97, sc2mac_dat_a_data98, sc2mac_dat_a_data99, sc2mac_dat_a_data100, sc2mac_dat_a_data101, sc2mac_dat_a_data102, sc2mac_dat_a_data103, sc2mac_dat_a_data104, sc2mac_dat_a_data105, sc2mac_dat_a_data106, sc2mac_dat_a_data107, sc2mac_dat_a_data108, sc2mac_dat_a_data109, sc2mac_dat_a_data110, sc2mac_dat_a_data111, sc2mac_dat_a_data112, sc2mac_dat_a_data113, sc2mac_dat_a_data114, sc2mac_dat_a_data115, sc2mac_dat_a_data116, sc2mac_dat_a_data117, sc2mac_dat_a_data118, sc2mac_dat_a_data119, sc2mac_dat_a_data120, sc2mac_dat_a_data121, sc2mac_dat_a_data122, sc2mac_dat_a_data123, sc2mac_dat_a_data124, sc2mac_dat_a_data125, sc2mac_dat_a_data126, sc2mac_dat_a_data127, sc2mac_dat_a_pd, sc2mac_dat_b_pvld, sc2mac_dat_b_mask, sc2mac_dat_b_data0, sc2mac_dat_b_data1, sc2mac_dat_b_data2, sc2mac_dat_b_data3, sc2mac_dat_b_data4, sc2mac_dat_b_data5, sc2mac_dat_b_data6, sc2mac_dat_b_data7, sc2mac_dat_b_data8, sc2mac_dat_b_data9, sc2mac_dat_b_data10, sc2mac_dat_b_data11, sc2mac_dat_b_data12, sc2mac_dat_b_data13, sc2mac_dat_b_data14, sc2mac_dat_b_data15, sc2mac_dat_b_data16, sc2mac_dat_b_data17, sc2mac_dat_b_data18, sc2mac_dat_b_data19, sc2mac_dat_b_data20, sc2mac_dat_b_data21, sc2mac_dat_b_data22, sc2mac_dat_b_data23, sc2mac_dat_b_data24, sc2mac_dat_b_data25, sc2mac_dat_b_data26, sc2mac_dat_b_data27, sc2mac_dat_b_data28, sc2mac_dat_b_data29, sc2mac_dat_b_data30, sc2mac_dat_b_data31, sc2mac_dat_b_data32, sc2mac_dat_b_data33, sc2mac_dat_b_data34, sc2mac_dat_b_data35, sc2mac_dat_b_data36, sc2mac_dat_b_data37, sc2mac_dat_b_data38, sc2mac_dat_b_data39, sc2mac_dat_b_data40, sc2mac_dat_b_data41, sc2mac_dat_b_data42, sc2mac_dat_b_data43, sc2mac_dat_b_data44, sc2mac_dat_b_data45, sc2mac_dat_b_data46, sc2mac_dat_b_data47, sc2mac_dat_b_data48, sc2mac_dat_b_data49, sc2mac_dat_b_data50, sc2mac_dat_b_data51, sc2mac_dat_b_data52, sc2mac_dat_b_data53, sc2mac_dat_b_data54, sc2mac_dat_b_data55, sc2mac_dat_b_data56, sc2mac_dat_b_data57, sc2mac_dat_b_data58, sc2mac_dat_b_data59, sc2mac_dat_b_data60, sc2mac_dat_b_data61, sc2mac_dat_b_data62, sc2mac_dat_b_data63, sc2mac_dat_b_data64, sc2mac_dat_b_data65, sc2mac_dat_b_data66, sc2mac_dat_b_data67, sc2mac_dat_b_data68, sc2mac_dat_b_data69, sc2mac_dat_b_data70, sc2mac_dat_b_data71, sc2mac_dat_b_data72, sc2mac_dat_b_data73, sc2mac_dat_b_data74, sc2mac_dat_b_data75, sc2mac_dat_b_data76, sc2mac_dat_b_data77, sc2mac_dat_b_data78, sc2mac_dat_b_data79, sc2mac_dat_b_data80, sc2mac_dat_b_data81, sc2mac_dat_b_data82, sc2mac_dat_b_data83, sc2mac_dat_b_data84, sc2mac_dat_b_data85, sc2mac_dat_b_data86, sc2mac_dat_b_data87, sc2mac_dat_b_data88, sc2mac_dat_b_data89, sc2mac_dat_b_data90, sc2mac_dat_b_data91, sc2mac_dat_b_data92, sc2mac_dat_b_data93, sc2mac_dat_b_data94, sc2mac_dat_b_data95, sc2mac_dat_b_data96, sc2mac_dat_b_data97, sc2mac_dat_b_data98, sc2mac_dat_b_data99, sc2mac_dat_b_data100, sc2mac_dat_b_data101, sc2mac_dat_b_data102, sc2mac_dat_b_data103, sc2mac_dat_b_data104, sc2mac_dat_b_data105, sc2mac_dat_b_data106, sc2mac_dat_b_data107, sc2mac_dat_b_data108, sc2mac_dat_b_data109, sc2mac_dat_b_data110, sc2mac_dat_b_data111, sc2mac_dat_b_data112, sc2mac_dat_b_data113, sc2mac_dat_b_data114, sc2mac_dat_b_data115, sc2mac_dat_b_data116, sc2mac_dat_b_data117, sc2mac_dat_b_data118, sc2mac_dat_b_data119, sc2mac_dat_b_data120, sc2mac_dat_b_data121, sc2mac_dat_b_data122, sc2mac_dat_b_data123, sc2mac_dat_b_data124, sc2mac_dat_b_data125, sc2mac_dat_b_data126, sc2mac_dat_b_data127, sc2mac_dat_b_pd, nvdla_core_ng_clk, nvdla_wg_clk, reg2dp_op_en, reg2dp_conv_mode, reg2dp_batches, reg2dp_proc_precision, reg2dp_datain_format, reg2dp_skip_data_rls, reg2dp_datain_channel_ext, reg2dp_datain_height_ext, reg2dp_datain_width_ext, reg2dp_y_extension, reg2dp_weight_channel_ext, reg2dp_entries, reg2dp_dataout_width, reg2dp_rls_slices, reg2dp_conv_x_stride_ext, reg2dp_conv_y_stride_ext, reg2dp_x_dilation_ext, reg2dp_y_dilation_ext, reg2dp_pad_left, reg2dp_pad_top, reg2dp_pad_value, reg2dp_data_bank, reg2dp_pra_truncate, slcg_wg_en);
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:3816" *)
  wire [4:0] _0000_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:8547" *)
  wire [4:0] _0001_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:11432" *)
  wire [11:0] _0002_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:11493" *)
  wire [11:0] _0003_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:3572" *)
  wire [3:0] _0004_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:3633" *)
  wire [3:0] _0005_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:6880" *)
  wire [11:0] _0006_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:14649" *)
  wire [511:0] _0007_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:14649" *)
  wire [511:0] _0008_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:14699" *)
  wire [511:0] _0009_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:14699" *)
  wire [511:0] _0010_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:14669" *)
  wire [511:0] _0011_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:14659" *)
  wire [511:0] _0012_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:14719" *)
  wire [511:0] _0013_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:14709" *)
  wire [511:0] _0014_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:14679" *)
  wire [511:0] _0015_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:14679" *)
  wire [511:0] _0016_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:14729" *)
  wire [511:0] _0017_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:14729" *)
  wire [511:0] _0018_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:14689" *)
  wire [511:0] _0019_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:14689" *)
  wire [511:0] _0020_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:14739" *)
  wire [511:0] _0021_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:14739" *)
  wire [511:0] _0022_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18172" *)
  wire [7:0] _0023_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18182" *)
  wire [7:0] _0024_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18192" *)
  wire [7:0] _0025_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17042" *)
  wire [7:0] _0026_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17052" *)
  wire [7:0] _0027_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17062" *)
  wire [7:0] _0028_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17072" *)
  wire [7:0] _0029_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17082" *)
  wire [7:0] _0030_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17092" *)
  wire [7:0] _0031_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17102" *)
  wire [7:0] _0032_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17112" *)
  wire [7:0] _0033_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16932" *)
  wire [7:0] _0034_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17122" *)
  wire [7:0] _0035_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17132" *)
  wire [7:0] _0036_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17142" *)
  wire [7:0] _0037_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17152" *)
  wire [7:0] _0038_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17162" *)
  wire [7:0] _0039_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17172" *)
  wire [7:0] _0040_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17182" *)
  wire [7:0] _0041_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17192" *)
  wire [7:0] _0042_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17202" *)
  wire [7:0] _0043_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17212" *)
  wire [7:0] _0044_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16942" *)
  wire [7:0] _0045_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17222" *)
  wire [7:0] _0046_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17232" *)
  wire [7:0] _0047_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17242" *)
  wire [7:0] _0048_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17252" *)
  wire [7:0] _0049_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17262" *)
  wire [7:0] _0050_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17272" *)
  wire [7:0] _0051_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17282" *)
  wire [7:0] _0052_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17292" *)
  wire [7:0] _0053_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17302" *)
  wire [7:0] _0054_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17312" *)
  wire [7:0] _0055_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16952" *)
  wire [7:0] _0056_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17322" *)
  wire [7:0] _0057_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17332" *)
  wire [7:0] _0058_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17342" *)
  wire [7:0] _0059_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17352" *)
  wire [7:0] _0060_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17362" *)
  wire [7:0] _0061_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17372" *)
  wire [7:0] _0062_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17382" *)
  wire [7:0] _0063_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17392" *)
  wire [7:0] _0064_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17402" *)
  wire [7:0] _0065_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17412" *)
  wire [7:0] _0066_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16962" *)
  wire [7:0] _0067_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17422" *)
  wire [7:0] _0068_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17432" *)
  wire [7:0] _0069_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17442" *)
  wire [7:0] _0070_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17452" *)
  wire [7:0] _0071_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17462" *)
  wire [7:0] _0072_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17472" *)
  wire [7:0] _0073_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17482" *)
  wire [7:0] _0074_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17492" *)
  wire [7:0] _0075_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17502" *)
  wire [7:0] _0076_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17512" *)
  wire [7:0] _0077_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16972" *)
  wire [7:0] _0078_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17522" *)
  wire [7:0] _0079_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17532" *)
  wire [7:0] _0080_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17542" *)
  wire [7:0] _0081_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17552" *)
  wire [7:0] _0082_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17562" *)
  wire [7:0] _0083_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17572" *)
  wire [7:0] _0084_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17582" *)
  wire [7:0] _0085_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17592" *)
  wire [7:0] _0086_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17602" *)
  wire [7:0] _0087_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17612" *)
  wire [7:0] _0088_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16982" *)
  wire [7:0] _0089_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17622" *)
  wire [7:0] _0090_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17632" *)
  wire [7:0] _0091_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17642" *)
  wire [7:0] _0092_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17652" *)
  wire [7:0] _0093_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17662" *)
  wire [7:0] _0094_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17672" *)
  wire [7:0] _0095_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17682" *)
  wire [7:0] _0096_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17692" *)
  wire [7:0] _0097_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17702" *)
  wire [7:0] _0098_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17712" *)
  wire [7:0] _0099_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16992" *)
  wire [7:0] _0100_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17722" *)
  wire [7:0] _0101_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17732" *)
  wire [7:0] _0102_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17742" *)
  wire [7:0] _0103_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17752" *)
  wire [7:0] _0104_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17762" *)
  wire [7:0] _0105_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17772" *)
  wire [7:0] _0106_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17782" *)
  wire [7:0] _0107_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17792" *)
  wire [7:0] _0108_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17802" *)
  wire [7:0] _0109_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17812" *)
  wire [7:0] _0110_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17002" *)
  wire [7:0] _0111_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17822" *)
  wire [7:0] _0112_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17832" *)
  wire [7:0] _0113_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17842" *)
  wire [7:0] _0114_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17852" *)
  wire [7:0] _0115_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17862" *)
  wire [7:0] _0116_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17872" *)
  wire [7:0] _0117_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17882" *)
  wire [7:0] _0118_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17892" *)
  wire [7:0] _0119_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17902" *)
  wire [7:0] _0120_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17912" *)
  wire [7:0] _0121_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17012" *)
  wire [7:0] _0122_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16922" *)
  wire [7:0] _0123_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17922" *)
  wire [7:0] _0124_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17932" *)
  wire [7:0] _0125_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17942" *)
  wire [7:0] _0126_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17952" *)
  wire [7:0] _0127_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17962" *)
  wire [7:0] _0128_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17972" *)
  wire [7:0] _0129_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17982" *)
  wire [7:0] _0130_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17992" *)
  wire [7:0] _0131_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18002" *)
  wire [7:0] _0132_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18012" *)
  wire [7:0] _0133_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17022" *)
  wire [7:0] _0134_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18022" *)
  wire [7:0] _0135_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18032" *)
  wire [7:0] _0136_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18042" *)
  wire [7:0] _0137_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18052" *)
  wire [7:0] _0138_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18062" *)
  wire [7:0] _0139_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18072" *)
  wire [7:0] _0140_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18082" *)
  wire [7:0] _0141_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18092" *)
  wire [7:0] _0142_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18102" *)
  wire [7:0] _0143_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18112" *)
  wire [7:0] _0144_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17032" *)
  wire [7:0] _0145_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18122" *)
  wire [7:0] _0146_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18132" *)
  wire [7:0] _0147_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18142" *)
  wire [7:0] _0148_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18152" *)
  wire [7:0] _0149_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18162" *)
  wire [7:0] _0150_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16861" *)
  wire [63:0] _0151_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16800" *)
  wire [63:0] _0152_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16739" *)
  wire [8:0] _0153_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16393" *)
  wire [8:0] _0154_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16461" *)
  wire [8:0] _0155_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16529" *)
  wire [8:0] _0156_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16597" *)
  wire [8:0] _0157_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16665" *)
  wire [8:0] _0158_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:9178" *)
  wire [7:0] _0159_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:12829" *)
  wire [7:0] _0160_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:10676" *)
  wire _0161_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:12707" *)
  wire _0162_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:10737" *)
  wire _0163_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:12768" *)
  wire _0164_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:10859" *)
  wire [1:0] _0165_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:12951" *)
  wire [1:0] _0166_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:10798" *)
  wire _0167_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:12890" *)
  wire _0168_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:10981" *)
  wire [8:0] _0169_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:13134" *)
  wire [8:0] _0170_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:11042" *)
  wire _0171_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:13073" *)
  wire _0172_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:10615" *)
  wire _0173_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:12646" *)
  wire _0174_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:12198" *)
  wire [11:0] _0175_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:12259" *)
  wire [11:0] _0176_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:12320" *)
  wire [11:0] _0177_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:12381" *)
  wire [11:0] _0178_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:10554" *)
  wire [1:0] _0179_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:12585" *)
  wire [1:0] _0180_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:10493" *)
  wire [1:0] _0181_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:12524" *)
  wire [1:0] _0182_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:10920" *)
  wire _0183_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:13012" *)
  wire _0184_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:13352" *)
  wire _0185_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:13549" *)
  wire _0186_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:13746" *)
  wire _0187_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:13943" *)
  wire _0188_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:14140" *)
  wire _0189_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:14337" *)
  wire _0190_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:13413" *)
  wire [1:0] _0191_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:13610" *)
  wire [1:0] _0192_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:13807" *)
  wire [1:0] _0193_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:14004" *)
  wire [1:0] _0194_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:14201" *)
  wire [1:0] _0195_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:14398" *)
  wire [1:0] _0196_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16147" *)
  wire [255:0] _0197_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16157" *)
  wire [255:0] _0198_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16167" *)
  wire [127:0] _0199_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16177" *)
  wire [127:0] _0200_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16187" *)
  wire [127:0] _0201_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16197" *)
  wire [127:0] _0202_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16207" *)
  wire [127:0] _0203_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16217" *)
  wire [127:0] _0204_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16227" *)
  wire [127:0] _0205_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16237" *)
  wire [127:0] _0206_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16247" *)
  wire [127:0] _0207_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16257" *)
  wire [127:0] _0208_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:14770" *)
  wire [26:0] _0209_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:14838" *)
  wire [26:0] _0210_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:14906" *)
  wire [26:0] _0211_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:14974" *)
  wire [26:0] _0212_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:13284" *)
  wire [28:0] _0213_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:13481" *)
  wire [28:0] _0214_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:13678" *)
  wire [28:0] _0215_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:13875" *)
  wire [28:0] _0216_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:14072" *)
  wire [28:0] _0217_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:14269" *)
  wire [28:0] _0218_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18220" *)
  wire [255:0] _0219_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18230" *)
  wire [255:0] _0220_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18240" *)
  wire [255:0] _0221_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18250" *)
  wire [255:0] _0222_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:2413" *)
  wire [3:0] _0223_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:3755" *)
  wire [5:0] _0224_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:9539" *)
  wire [10:0] _0225_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:2657" *)
  wire [10:0] _0226_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:10280" *)
  wire [13:0] _0227_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:10341" *)
  wire [13:0] _0228_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:2596" *)
  wire [12:0] _0229_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:9744" *)
  wire [13:0] _0230_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:9805" *)
  wire [13:0] _0231_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:2474" *)
  wire [13:0] _0232_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:2535" *)
  wire [12:0] _0233_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:9387" *)
  wire [12:0] _0234_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:9448" *)
  wire [12:0] _0235_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:5158" *)
  wire [12:0] _0236_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:7890" *)
  wire [30:0] _0237_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:7958" *)
  wire [30:0] _0238_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:8026" *)
  wire [30:0] _0239_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:8094" *)
  wire [30:0] _0240_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:8162" *)
  wire [30:0] _0241_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18627" *)
  wire [7:0] _0242_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:19627" *)
  wire [7:0] _0243_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:19637" *)
  wire [7:0] _0244_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:19647" *)
  wire [7:0] _0245_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:19657" *)
  wire [7:0] _0246_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:19667" *)
  wire [7:0] _0247_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:19677" *)
  wire [7:0] _0248_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:19687" *)
  wire [7:0] _0249_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:19697" *)
  wire [7:0] _0250_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:19707" *)
  wire [7:0] _0251_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:19717" *)
  wire [7:0] _0252_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18727" *)
  wire [7:0] _0253_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:19727" *)
  wire [7:0] _0254_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:19737" *)
  wire [7:0] _0255_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:19747" *)
  wire [7:0] _0256_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:19757" *)
  wire [7:0] _0257_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:19767" *)
  wire [7:0] _0258_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:19777" *)
  wire [7:0] _0259_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:19787" *)
  wire [7:0] _0260_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:19797" *)
  wire [7:0] _0261_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:19807" *)
  wire [7:0] _0262_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:19817" *)
  wire [7:0] _0263_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18737" *)
  wire [7:0] _0264_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:19827" *)
  wire [7:0] _0265_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:19837" *)
  wire [7:0] _0266_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:19847" *)
  wire [7:0] _0267_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:19857" *)
  wire [7:0] _0268_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:19867" *)
  wire [7:0] _0269_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:19877" *)
  wire [7:0] _0270_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:19887" *)
  wire [7:0] _0271_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:19897" *)
  wire [7:0] _0272_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18747" *)
  wire [7:0] _0273_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18757" *)
  wire [7:0] _0274_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18767" *)
  wire [7:0] _0275_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18777" *)
  wire [7:0] _0276_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18787" *)
  wire [7:0] _0277_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18797" *)
  wire [7:0] _0278_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18807" *)
  wire [7:0] _0279_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18817" *)
  wire [7:0] _0280_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18637" *)
  wire [7:0] _0281_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18827" *)
  wire [7:0] _0282_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18837" *)
  wire [7:0] _0283_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18847" *)
  wire [7:0] _0284_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18857" *)
  wire [7:0] _0285_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18867" *)
  wire [7:0] _0286_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18877" *)
  wire [7:0] _0287_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18887" *)
  wire [7:0] _0288_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18897" *)
  wire [7:0] _0289_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18907" *)
  wire [7:0] _0290_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18917" *)
  wire [7:0] _0291_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18647" *)
  wire [7:0] _0292_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18927" *)
  wire [7:0] _0293_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18937" *)
  wire [7:0] _0294_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18947" *)
  wire [7:0] _0295_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18957" *)
  wire [7:0] _0296_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18967" *)
  wire [7:0] _0297_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18977" *)
  wire [7:0] _0298_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18987" *)
  wire [7:0] _0299_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18997" *)
  wire [7:0] _0300_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:19007" *)
  wire [7:0] _0301_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:19017" *)
  wire [7:0] _0302_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18657" *)
  wire [7:0] _0303_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:19027" *)
  wire [7:0] _0304_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:19037" *)
  wire [7:0] _0305_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:19047" *)
  wire [7:0] _0306_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:19057" *)
  wire [7:0] _0307_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:19067" *)
  wire [7:0] _0308_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:19077" *)
  wire [7:0] _0309_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:19087" *)
  wire [7:0] _0310_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:19097" *)
  wire [7:0] _0311_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:19107" *)
  wire [7:0] _0312_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:19117" *)
  wire [7:0] _0313_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18667" *)
  wire [7:0] _0314_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:19127" *)
  wire [7:0] _0315_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:19137" *)
  wire [7:0] _0316_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:19147" *)
  wire [7:0] _0317_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:19157" *)
  wire [7:0] _0318_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:19167" *)
  wire [7:0] _0319_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:19177" *)
  wire [7:0] _0320_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:19187" *)
  wire [7:0] _0321_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:19197" *)
  wire [7:0] _0322_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:19207" *)
  wire [7:0] _0323_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:19217" *)
  wire [7:0] _0324_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18677" *)
  wire [7:0] _0325_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:19227" *)
  wire [7:0] _0326_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:19237" *)
  wire [7:0] _0327_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:19247" *)
  wire [7:0] _0328_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:19257" *)
  wire [7:0] _0329_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:19267" *)
  wire [7:0] _0330_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:19277" *)
  wire [7:0] _0331_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:19287" *)
  wire [7:0] _0332_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:19297" *)
  wire [7:0] _0333_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:19307" *)
  wire [7:0] _0334_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:19317" *)
  wire [7:0] _0335_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18687" *)
  wire [7:0] _0336_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:19327" *)
  wire [7:0] _0337_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:19337" *)
  wire [7:0] _0338_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:19347" *)
  wire [7:0] _0339_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:19357" *)
  wire [7:0] _0340_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:19367" *)
  wire [7:0] _0341_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:19377" *)
  wire [7:0] _0342_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:19387" *)
  wire [7:0] _0343_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:19397" *)
  wire [7:0] _0344_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:19407" *)
  wire [7:0] _0345_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:19417" *)
  wire [7:0] _0346_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18697" *)
  wire [7:0] _0347_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:19427" *)
  wire [7:0] _0348_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:19437" *)
  wire [7:0] _0349_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:19447" *)
  wire [7:0] _0350_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:19457" *)
  wire [7:0] _0351_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:19467" *)
  wire [7:0] _0352_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:19477" *)
  wire [7:0] _0353_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:19487" *)
  wire [7:0] _0354_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:19497" *)
  wire [7:0] _0355_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:19507" *)
  wire [7:0] _0356_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:19517" *)
  wire [7:0] _0357_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18707" *)
  wire [7:0] _0358_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:19527" *)
  wire [7:0] _0359_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:19537" *)
  wire [7:0] _0360_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:19547" *)
  wire [7:0] _0361_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:19557" *)
  wire [7:0] _0362_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:19567" *)
  wire [7:0] _0363_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:19577" *)
  wire [7:0] _0364_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:19587" *)
  wire [7:0] _0365_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:19597" *)
  wire [7:0] _0366_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:19607" *)
  wire [7:0] _0367_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:19617" *)
  wire [7:0] _0368_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18717" *)
  wire [7:0] _0369_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18566" *)
  wire [8:0] _0370_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18505" *)
  wire [127:0] _0371_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:8234" *)
  wire [30:0] _0372_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:8302" *)
  wire [30:0] _0373_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:8370" *)
  wire [30:0] _0374_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:8438" *)
  wire [30:0] _0375_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:4365" *)
  wire [11:0] _0376_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:4426" *)
  wire [11:0] _0377_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:4487" *)
  wire [11:0] _0378_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:11554" *)
  wire [11:0] _0379_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:4609" *)
  wire [11:0] _0380_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:11615" *)
  wire [11:0] _0381_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:4670" *)
  wire [11:0] _0382_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:11676" *)
  wire [11:0] _0383_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:4731" *)
  wire [11:0] _0384_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:11737" *)
  wire [11:0] _0385_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:4792" *)
  wire [11:0] _0386_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:4548" *)
  wire [11:0] _0387_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:2352" *)
  wire [1:0] _0388_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:2230" *)
  wire [33:0] _0389_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:2291" *)
  wire [22:0] _0390_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:2169" *)
  wire [21:0] _0391_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:5097" *)
  wire [11:0] _0392_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:5036" *)
  wire [11:0] _0393_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:4304" *)
  wire [15:0] _0394_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:4121" *)
  wire [11:0] _0395_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:11164" *)
  wire _0396_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:11103" *)
  wire _0397_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:10049" *)
  wire _0398_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:10110" *)
  wire _0399_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:9988" *)
  wire [15:0] _0400_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:9866" *)
  wire [15:0] _0401_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:9927" *)
  wire [15:0] _0402_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:3999" *)
  wire [6:0] _0403_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:4060" *)
  wire [6:0] _0404_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:3877" *)
  wire [5:0] _0405_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:3938" *)
  wire [6:0] _0406_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:3694" *)
  wire _0407_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:5280" *)
  wire [7:0] _0408_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:5219" *)
  wire [7:0] _0409_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:4914" *)
  wire [11:0] _0410_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:4853" *)
  wire [11:0] _0411_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15266" *)
  wire [7:0] _0412_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15510" *)
  wire [7:0] _0413_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15327" *)
  wire [7:0] _0414_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15571" *)
  wire [7:0] _0415_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15388" *)
  wire [7:0] _0416_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15632" *)
  wire [7:0] _0417_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15449" *)
  wire [7:0] _0418_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15693" *)
  wire [7:0] _0419_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:12449" *)
  wire [11:0] _0420_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:7532" *)
  wire [11:0] _0421_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:7471" *)
  wire [11:0] _0422_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:20181" *)
  wire [7:0] _0423_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21181" *)
  wire [7:0] _0424_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21191" *)
  wire [7:0] _0425_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21201" *)
  wire [7:0] _0426_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21211" *)
  wire [7:0] _0427_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21221" *)
  wire [7:0] _0428_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21231" *)
  wire [7:0] _0429_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21241" *)
  wire [7:0] _0430_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21251" *)
  wire [7:0] _0431_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21261" *)
  wire [7:0] _0432_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21271" *)
  wire [7:0] _0433_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:20281" *)
  wire [7:0] _0434_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21281" *)
  wire [7:0] _0435_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21291" *)
  wire [7:0] _0436_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21301" *)
  wire [7:0] _0437_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21311" *)
  wire [7:0] _0438_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21321" *)
  wire [7:0] _0439_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21331" *)
  wire [7:0] _0440_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21341" *)
  wire [7:0] _0441_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21351" *)
  wire [7:0] _0442_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21361" *)
  wire [7:0] _0443_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21371" *)
  wire [7:0] _0444_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:20291" *)
  wire [7:0] _0445_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21381" *)
  wire [7:0] _0446_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21391" *)
  wire [7:0] _0447_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21401" *)
  wire [7:0] _0448_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21411" *)
  wire [7:0] _0449_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21421" *)
  wire [7:0] _0450_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21431" *)
  wire [7:0] _0451_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21441" *)
  wire [7:0] _0452_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21451" *)
  wire [7:0] _0453_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:20301" *)
  wire [7:0] _0454_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:20311" *)
  wire [7:0] _0455_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:20321" *)
  wire [7:0] _0456_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:20331" *)
  wire [7:0] _0457_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:20341" *)
  wire [7:0] _0458_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:20351" *)
  wire [7:0] _0459_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:20361" *)
  wire [7:0] _0460_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:20371" *)
  wire [7:0] _0461_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:20191" *)
  wire [7:0] _0462_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:20381" *)
  wire [7:0] _0463_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:20391" *)
  wire [7:0] _0464_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:20401" *)
  wire [7:0] _0465_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:20411" *)
  wire [7:0] _0466_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:20421" *)
  wire [7:0] _0467_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:20431" *)
  wire [7:0] _0468_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:20441" *)
  wire [7:0] _0469_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:20451" *)
  wire [7:0] _0470_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:20461" *)
  wire [7:0] _0471_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:20471" *)
  wire [7:0] _0472_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:20201" *)
  wire [7:0] _0473_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:20481" *)
  wire [7:0] _0474_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:20491" *)
  wire [7:0] _0475_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:20501" *)
  wire [7:0] _0476_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:20511" *)
  wire [7:0] _0477_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:20521" *)
  wire [7:0] _0478_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:20531" *)
  wire [7:0] _0479_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:20541" *)
  wire [7:0] _0480_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:20551" *)
  wire [7:0] _0481_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:20561" *)
  wire [7:0] _0482_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:20571" *)
  wire [7:0] _0483_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:20211" *)
  wire [7:0] _0484_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:20581" *)
  wire [7:0] _0485_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:20591" *)
  wire [7:0] _0486_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:20601" *)
  wire [7:0] _0487_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:20611" *)
  wire [7:0] _0488_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:20621" *)
  wire [7:0] _0489_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:20631" *)
  wire [7:0] _0490_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:20641" *)
  wire [7:0] _0491_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:20651" *)
  wire [7:0] _0492_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:20661" *)
  wire [7:0] _0493_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:20671" *)
  wire [7:0] _0494_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:20221" *)
  wire [7:0] _0495_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:20681" *)
  wire [7:0] _0496_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:20691" *)
  wire [7:0] _0497_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:20701" *)
  wire [7:0] _0498_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:20711" *)
  wire [7:0] _0499_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:20721" *)
  wire [7:0] _0500_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:20731" *)
  wire [7:0] _0501_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:20741" *)
  wire [7:0] _0502_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:20751" *)
  wire [7:0] _0503_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:20761" *)
  wire [7:0] _0504_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:20771" *)
  wire [7:0] _0505_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:20231" *)
  wire [7:0] _0506_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:20781" *)
  wire [7:0] _0507_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:20791" *)
  wire [7:0] _0508_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:20801" *)
  wire [7:0] _0509_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:20811" *)
  wire [7:0] _0510_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:20821" *)
  wire [7:0] _0511_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:20831" *)
  wire [7:0] _0512_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:20841" *)
  wire [7:0] _0513_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:20851" *)
  wire [7:0] _0514_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:20861" *)
  wire [7:0] _0515_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:20871" *)
  wire [7:0] _0516_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:20241" *)
  wire [7:0] _0517_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:20881" *)
  wire [7:0] _0518_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:20891" *)
  wire [7:0] _0519_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:20901" *)
  wire [7:0] _0520_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:20911" *)
  wire [7:0] _0521_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:20921" *)
  wire [7:0] _0522_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:20931" *)
  wire [7:0] _0523_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:20941" *)
  wire [7:0] _0524_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:20951" *)
  wire [7:0] _0525_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:20961" *)
  wire [7:0] _0526_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:20971" *)
  wire [7:0] _0527_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:20251" *)
  wire [7:0] _0528_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:20981" *)
  wire [7:0] _0529_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:20991" *)
  wire [7:0] _0530_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21001" *)
  wire [7:0] _0531_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21011" *)
  wire [7:0] _0532_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21021" *)
  wire [7:0] _0533_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21031" *)
  wire [7:0] _0534_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21041" *)
  wire [7:0] _0535_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21051" *)
  wire [7:0] _0536_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21061" *)
  wire [7:0] _0537_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21071" *)
  wire [7:0] _0538_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:20261" *)
  wire [7:0] _0539_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21081" *)
  wire [7:0] _0540_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21091" *)
  wire [7:0] _0541_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21101" *)
  wire [7:0] _0542_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21111" *)
  wire [7:0] _0543_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21121" *)
  wire [7:0] _0544_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21131" *)
  wire [7:0] _0545_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21141" *)
  wire [7:0] _0546_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21151" *)
  wire [7:0] _0547_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21161" *)
  wire [7:0] _0548_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21171" *)
  wire [7:0] _0549_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:20271" *)
  wire [7:0] _0550_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:20059" *)
  wire [127:0] _0551_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:19937" *)
  wire [8:0] _0552_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21461" *)
  wire [7:0] _0553_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:22461" *)
  wire [7:0] _0554_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:22471" *)
  wire [7:0] _0555_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:22481" *)
  wire [7:0] _0556_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:22491" *)
  wire [7:0] _0557_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:22501" *)
  wire [7:0] _0558_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:22511" *)
  wire [7:0] _0559_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:22521" *)
  wire [7:0] _0560_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:22531" *)
  wire [7:0] _0561_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:22541" *)
  wire [7:0] _0562_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:22551" *)
  wire [7:0] _0563_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21561" *)
  wire [7:0] _0564_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:22561" *)
  wire [7:0] _0565_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:22571" *)
  wire [7:0] _0566_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:22581" *)
  wire [7:0] _0567_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:22591" *)
  wire [7:0] _0568_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:22601" *)
  wire [7:0] _0569_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:22611" *)
  wire [7:0] _0570_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:22621" *)
  wire [7:0] _0571_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:22631" *)
  wire [7:0] _0572_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:22641" *)
  wire [7:0] _0573_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:22651" *)
  wire [7:0] _0574_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21571" *)
  wire [7:0] _0575_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:22661" *)
  wire [7:0] _0576_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:22671" *)
  wire [7:0] _0577_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:22681" *)
  wire [7:0] _0578_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:22691" *)
  wire [7:0] _0579_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:22701" *)
  wire [7:0] _0580_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:22711" *)
  wire [7:0] _0581_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:22721" *)
  wire [7:0] _0582_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:22731" *)
  wire [7:0] _0583_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21581" *)
  wire [7:0] _0584_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21591" *)
  wire [7:0] _0585_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21601" *)
  wire [7:0] _0586_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21611" *)
  wire [7:0] _0587_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21621" *)
  wire [7:0] _0588_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21631" *)
  wire [7:0] _0589_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21641" *)
  wire [7:0] _0590_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21651" *)
  wire [7:0] _0591_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21471" *)
  wire [7:0] _0592_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21661" *)
  wire [7:0] _0593_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21671" *)
  wire [7:0] _0594_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21681" *)
  wire [7:0] _0595_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21691" *)
  wire [7:0] _0596_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21701" *)
  wire [7:0] _0597_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21711" *)
  wire [7:0] _0598_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21721" *)
  wire [7:0] _0599_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21731" *)
  wire [7:0] _0600_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21741" *)
  wire [7:0] _0601_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21751" *)
  wire [7:0] _0602_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21481" *)
  wire [7:0] _0603_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21761" *)
  wire [7:0] _0604_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21771" *)
  wire [7:0] _0605_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21781" *)
  wire [7:0] _0606_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21791" *)
  wire [7:0] _0607_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21801" *)
  wire [7:0] _0608_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21811" *)
  wire [7:0] _0609_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21821" *)
  wire [7:0] _0610_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21831" *)
  wire [7:0] _0611_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21841" *)
  wire [7:0] _0612_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21851" *)
  wire [7:0] _0613_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21491" *)
  wire [7:0] _0614_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21861" *)
  wire [7:0] _0615_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21871" *)
  wire [7:0] _0616_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21881" *)
  wire [7:0] _0617_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21891" *)
  wire [7:0] _0618_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21901" *)
  wire [7:0] _0619_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21911" *)
  wire [7:0] _0620_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21921" *)
  wire [7:0] _0621_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21931" *)
  wire [7:0] _0622_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21941" *)
  wire [7:0] _0623_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21951" *)
  wire [7:0] _0624_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21501" *)
  wire [7:0] _0625_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21961" *)
  wire [7:0] _0626_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21971" *)
  wire [7:0] _0627_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21981" *)
  wire [7:0] _0628_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21991" *)
  wire [7:0] _0629_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:22001" *)
  wire [7:0] _0630_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:22011" *)
  wire [7:0] _0631_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:22021" *)
  wire [7:0] _0632_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:22031" *)
  wire [7:0] _0633_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:22041" *)
  wire [7:0] _0634_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:22051" *)
  wire [7:0] _0635_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21511" *)
  wire [7:0] _0636_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:22061" *)
  wire [7:0] _0637_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:22071" *)
  wire [7:0] _0638_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:22081" *)
  wire [7:0] _0639_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:22091" *)
  wire [7:0] _0640_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:22101" *)
  wire [7:0] _0641_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:22111" *)
  wire [7:0] _0642_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:22121" *)
  wire [7:0] _0643_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:22131" *)
  wire [7:0] _0644_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:22141" *)
  wire [7:0] _0645_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:22151" *)
  wire [7:0] _0646_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21521" *)
  wire [7:0] _0647_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:22161" *)
  wire [7:0] _0648_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:22171" *)
  wire [7:0] _0649_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:22181" *)
  wire [7:0] _0650_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:22191" *)
  wire [7:0] _0651_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:22201" *)
  wire [7:0] _0652_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:22211" *)
  wire [7:0] _0653_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:22221" *)
  wire [7:0] _0654_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:22231" *)
  wire [7:0] _0655_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:22241" *)
  wire [7:0] _0656_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:22251" *)
  wire [7:0] _0657_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21531" *)
  wire [7:0] _0658_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:22261" *)
  wire [7:0] _0659_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:22271" *)
  wire [7:0] _0660_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:22281" *)
  wire [7:0] _0661_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:22291" *)
  wire [7:0] _0662_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:22301" *)
  wire [7:0] _0663_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:22311" *)
  wire [7:0] _0664_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:22321" *)
  wire [7:0] _0665_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:22331" *)
  wire [7:0] _0666_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:22341" *)
  wire [7:0] _0667_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:22351" *)
  wire [7:0] _0668_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21541" *)
  wire [7:0] _0669_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:22361" *)
  wire [7:0] _0670_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:22371" *)
  wire [7:0] _0671_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:22381" *)
  wire [7:0] _0672_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:22391" *)
  wire [7:0] _0673_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:22401" *)
  wire [7:0] _0674_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:22411" *)
  wire [7:0] _0675_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:22421" *)
  wire [7:0] _0676_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:22431" *)
  wire [7:0] _0677_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:22441" *)
  wire [7:0] _0678_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:22451" *)
  wire [7:0] _0679_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21551" *)
  wire [7:0] _0680_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:20120" *)
  wire [127:0] _0681_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:19998" *)
  wire [8:0] _0682_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:4975" *)
  wire [11:0] _0683_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:8831" *)
  wire [6:0] _0684_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:3450" *)
  wire [2:0] _0685_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:3511" *)
  wire [2:0] _0686_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:8730" *)
  wire [1:0] _0687_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:2718" *)
  wire [2:0] _0688_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:3328" *)
  wire [2:0] _0689_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:3389" *)
  wire [2:0] _0690_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:2779" *)
  wire [2:0] _0691_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:2840" *)
  wire [1:0] _0692_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:2901" *)
  wire [2:0] _0693_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:2962" *)
  wire [2:0] _0694_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:3023" *)
  wire [2:0] _0695_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:3084" *)
  wire [2:0] _0696_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:3145" *)
  wire [2:0] _0697_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:3206" *)
  wire [2:0] _0698_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:3267" *)
  wire [2:0] _0699_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:11798" *)
  wire [11:0] _0700_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:4182" *)
  wire [5:0] _0701_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:4243" *)
  wire [5:0] _0702_;
  wire [13:0] _0703_;
  wire [11:0] _0704_;
  wire [11:0] _0705_;
  wire [11:0] _0706_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:12157" *)
  wire [12:0] _0707_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:12157" *)
  wire [12:0] _0708_;
  wire [7:0] _0709_;
  wire [7:0] _0710_;
  wire [7:0] _0711_;
  wire [7:0] _0712_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1941" *)
  wire [5:0] _0713_;
  wire [11:0] _0714_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1965" *)
  wire [13:0] _0715_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:2011" *)
  wire [3:0] _0716_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:2018" *)
  wire [5:0] _0717_;
  wire [5:0] _0718_;
  wire [5:0] _0719_;
  wire [5:0] _0720_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:2061" *)
  wire [3:0] _0721_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:2069" *)
  wire [5:0] _0722_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:2077" *)
  wire [5:0] _0723_;
  wire [11:0] _0724_;
  wire [11:0] _0725_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:8539" *)
  (* unused_bits = "5" *)
  wire [5:0] _0726_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:9616" *)
  (* unused_bits = "14" *)
  wire [14:0] _0727_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:9617" *)
  (* unused_bits = "14" *)
  wire [14:0] _0728_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:9656" *)
  (* unused_bits = "16" *)
  wire [16:0] _0729_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:9657" *)
  (* unused_bits = "16" *)
  wire [16:0] _0730_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:9659" *)
  (* unused_bits = "16" *)
  wire [16:0] _0731_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:10244" *)
  wire _0732_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:10245" *)
  wire _0733_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:10256" *)
  wire _0734_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:10264" *)
  wire _0735_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:10264" *)
  wire _0736_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:10417" *)
  wire _0737_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:10448" *)
  wire _0738_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:10448" *)
  wire _0739_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:10455" *)
  wire _0740_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:10464" *)
  wire _0741_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:11047" *)
  wire _0742_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:11047" *)
  wire _0743_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:11330" *)
  wire _0744_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:11342" *)
  wire _0745_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:11351" *)
  wire _0746_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:11391" *)
  wire _0747_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:12194" *)
  wire _0748_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:12195" *)
  wire _0749_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:12196" *)
  wire _0750_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:12197" *)
  wire _0751_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:14552" *)
  wire _0752_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:14553" *)
  wire _0753_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:14553" *)
  wire _0754_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:14554" *)
  wire _0755_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:14555" *)
  wire _0756_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:14555" *)
  wire _0757_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:14556" *)
  wire _0758_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:14557" *)
  wire _0759_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:14558" *)
  wire _0760_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:14560" *)
  wire _0761_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:14564" *)
  wire _0762_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:14581" *)
  wire _0763_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:14584" *)
  wire _0764_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:14587" *)
  wire _0765_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15041" *)
  wire _0766_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15042" *)
  wire _0767_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15043" *)
  wire _0768_;
  wire [11:0] _0769_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15063" *)
  wire [26:0] _0770_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15064" *)
  wire [26:0] _0771_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15176" *)
  wire _0772_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15177" *)
  wire _0773_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15177" *)
  wire _0774_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15178" *)
  wire _0775_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15179" *)
  wire [7:0] _0776_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15192" *)
  wire _0777_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15193" *)
  wire _0778_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15193" *)
  wire _0779_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15194" *)
  wire _0780_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15195" *)
  wire [7:0] _0781_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15208" *)
  wire _0782_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15209" *)
  wire _0783_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15209" *)
  wire _0784_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15210" *)
  wire _0785_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15211" *)
  wire [7:0] _0786_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15224" *)
  wire _0787_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15225" *)
  wire _0788_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15225" *)
  wire _0789_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15226" *)
  wire _0790_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15227" *)
  wire [7:0] _0791_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15239" *)
  wire _0792_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15240" *)
  wire _0793_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15240" *)
  wire _0794_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15241" *)
  wire _0795_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15241" *)
  wire _0796_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15242" *)
  wire _0797_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15242" *)
  wire _0798_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15261" *)
  wire _0799_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15261" *)
  wire _0800_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15261" *)
  wire _0801_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15262" *)
  wire _0802_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15262" *)
  wire _0803_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15262" *)
  wire _0804_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15262" *)
  wire _0805_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15263" *)
  wire _0806_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15263" *)
  wire _0807_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15263" *)
  wire _0808_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15263" *)
  wire _0809_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15264" *)
  wire _0810_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15264" *)
  wire _0811_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15264" *)
  wire _0812_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15264" *)
  wire _0813_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15811" *)
  wire [1023:0] _0814_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15812" *)
  wire [1023:0] _0815_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15813" *)
  wire [1023:0] _0816_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15814" *)
  wire [1023:0] _0817_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15856" *)
  wire [255:0] _0818_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15857" *)
  wire [255:0] _0819_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15858" *)
  wire [255:0] _0820_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15868" *)
  wire [255:0] _0821_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15869" *)
  wire [255:0] _0822_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15870" *)
  wire [255:0] _0823_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15880" *)
  wire [255:0] _0824_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15881" *)
  wire [255:0] _0825_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15882" *)
  wire [255:0] _0826_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15892" *)
  wire [255:0] _0827_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15893" *)
  wire [255:0] _0828_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15894" *)
  wire [255:0] _0829_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15961" *)
  wire _0830_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15961" *)
  wire _0831_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15962" *)
  wire _0832_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15963" *)
  wire _0833_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15964" *)
  wire _0834_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15965" *)
  wire _0835_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15966" *)
  wire _0836_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15981" *)
  wire _0837_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15986" *)
  wire _0838_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16302" *)
  wire [127:0] _0839_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16303" *)
  wire [127:0] _0840_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16312" *)
  wire [63:0] _0841_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16313" *)
  wire [63:0] _0842_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16369" *)
  wire [63:0] _0843_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16370" *)
  wire [127:0] _0844_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16371" *)
  wire [127:0] _0845_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16378" *)
  wire _0846_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16923" *)
  wire _0847_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16933" *)
  wire _0848_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16943" *)
  wire _0849_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16953" *)
  wire _0850_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16963" *)
  wire _0851_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16973" *)
  wire _0852_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16983" *)
  wire _0853_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16993" *)
  wire _0854_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17003" *)
  wire _0855_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17013" *)
  wire _0856_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17023" *)
  wire _0857_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17033" *)
  wire _0858_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17043" *)
  wire _0859_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17053" *)
  wire _0860_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17063" *)
  wire _0861_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17073" *)
  wire _0862_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17083" *)
  wire _0863_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17093" *)
  wire _0864_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17103" *)
  wire _0865_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17113" *)
  wire _0866_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17123" *)
  wire _0867_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17133" *)
  wire _0868_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17143" *)
  wire _0869_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17153" *)
  wire _0870_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17163" *)
  wire _0871_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17173" *)
  wire _0872_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17183" *)
  wire _0873_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17193" *)
  wire _0874_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17203" *)
  wire _0875_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17213" *)
  wire _0876_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17223" *)
  wire _0877_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17233" *)
  wire _0878_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17243" *)
  wire _0879_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17253" *)
  wire _0880_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17263" *)
  wire _0881_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17273" *)
  wire _0882_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17283" *)
  wire _0883_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17293" *)
  wire _0884_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17303" *)
  wire _0885_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17313" *)
  wire _0886_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17323" *)
  wire _0887_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17333" *)
  wire _0888_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17343" *)
  wire _0889_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17353" *)
  wire _0890_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17363" *)
  wire _0891_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17373" *)
  wire _0892_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17383" *)
  wire _0893_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17393" *)
  wire _0894_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17403" *)
  wire _0895_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17413" *)
  wire _0896_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17423" *)
  wire _0897_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17433" *)
  wire _0898_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17443" *)
  wire _0899_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17453" *)
  wire _0900_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17463" *)
  wire _0901_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17473" *)
  wire _0902_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17483" *)
  wire _0903_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17493" *)
  wire _0904_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17503" *)
  wire _0905_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17513" *)
  wire _0906_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17523" *)
  wire _0907_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17533" *)
  wire _0908_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17543" *)
  wire _0909_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17553" *)
  wire _0910_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17563" *)
  wire _0911_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17573" *)
  wire _0912_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17583" *)
  wire _0913_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17593" *)
  wire _0914_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17603" *)
  wire _0915_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17613" *)
  wire _0916_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17623" *)
  wire _0917_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17633" *)
  wire _0918_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17643" *)
  wire _0919_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17653" *)
  wire _0920_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17663" *)
  wire _0921_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17673" *)
  wire _0922_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17683" *)
  wire _0923_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17693" *)
  wire _0924_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17703" *)
  wire _0925_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17713" *)
  wire _0926_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17723" *)
  wire _0927_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17733" *)
  wire _0928_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17743" *)
  wire _0929_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17753" *)
  wire _0930_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17763" *)
  wire _0931_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17773" *)
  wire _0932_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17783" *)
  wire _0933_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17793" *)
  wire _0934_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17803" *)
  wire _0935_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17813" *)
  wire _0936_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17823" *)
  wire _0937_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17833" *)
  wire _0938_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17843" *)
  wire _0939_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17853" *)
  wire _0940_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17863" *)
  wire _0941_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17873" *)
  wire _0942_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17883" *)
  wire _0943_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17893" *)
  wire _0944_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17903" *)
  wire _0945_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17913" *)
  wire _0946_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17923" *)
  wire _0947_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17933" *)
  wire _0948_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17943" *)
  wire _0949_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17953" *)
  wire _0950_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17963" *)
  wire _0951_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17973" *)
  wire _0952_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17983" *)
  wire _0953_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17993" *)
  wire _0954_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18003" *)
  wire _0955_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18013" *)
  wire _0956_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18023" *)
  wire _0957_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18033" *)
  wire _0958_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18043" *)
  wire _0959_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18053" *)
  wire _0960_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18063" *)
  wire _0961_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18073" *)
  wire _0962_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18083" *)
  wire _0963_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18093" *)
  wire _0964_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18103" *)
  wire _0965_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18113" *)
  wire _0966_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18123" *)
  wire _0967_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18133" *)
  wire _0968_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18143" *)
  wire _0969_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18153" *)
  wire _0970_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18163" *)
  wire _0971_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18173" *)
  wire _0972_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18183" *)
  wire _0973_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18193" *)
  wire _0974_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:7446" *)
  wire _0975_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:7446" *)
  wire _0976_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:8505" *)
  wire _0977_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:8506" *)
  wire _0978_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:8507" *)
  wire _0979_;
  wire [12:0] _0980_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:8516" *)
  wire [30:0] _0981_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:8517" *)
  wire [30:0] _0982_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:8728" *)
  wire _0983_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:8807" *)
  wire _0984_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:8829" *)
  wire _0985_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:9100" *)
  wire _0986_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:9100" *)
  wire _0987_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:9348" *)
  wire _0988_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:9377" *)
  wire _0989_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:9655" *)
  wire _0990_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:9655" *)
  wire _0991_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:9655" *)
  wire _0992_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:9656" *)
  wire _0993_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:9657" *)
  wire _0994_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:9658" *)
  wire _0995_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:9669" *)
  wire _0996_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:9678" *)
  wire _0997_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:9678" *)
  wire _0998_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:9678" *)
  wire _0999_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:9687" *)
  wire _1000_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:9687" *)
  wire _1001_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:9696" *)
  wire _1002_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:9696" *)
  wire _1003_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:9696" *)
  wire _1004_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:9706" *)
  wire _1005_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:9706" *)
  wire _1006_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:9706" *)
  wire _1007_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:9706" *)
  wire _1008_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:9732" *)
  wire _1009_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:9733" *)
  wire _1010_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:9733" *)
  wire _1011_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:9733" *)
  wire _1012_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:9734" *)
  wire _1013_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:9735" *)
  wire _1014_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:9740" *)
  wire _1015_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:9743" *)
  wire _1016_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15062" *)
  wire [26:0] _1017_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:8515" *)
  wire [30:0] _1018_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:11388" *)
  (* unused_bits = "12 13" *)
  wire [13:0] _1019_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:2134" *)
  (* unused_bits = "12 13 14 15" *)
  wire [15:0] _1020_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:11407" *)
  wire [14:0] _1021_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:11407" *)
  wire [14:0] _1022_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:11407" *)
  wire [14:0] _1023_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:11421" *)
  wire [14:0] _1024_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:11421" *)
  wire [14:0] _1025_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:10474" *)
  wire _1026_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:12190" *)
  wire _1027_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:12191" *)
  wire _1028_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:12192" *)
  wire _1029_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:12197" *)
  wire _1030_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:12453" *)
  wire _1031_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:14531" *)
  wire _1032_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:14532" *)
  wire _1033_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:14535" *)
  wire _1034_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:14537" *)
  wire _1035_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15241" *)
  wire _1036_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15263" *)
  wire _1037_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15961" *)
  wire _1038_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15963" *)
  wire _1039_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15964" *)
  wire _1040_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15965" *)
  wire _1041_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15966" *)
  wire _1042_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16105" *)
  wire _1043_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16106" *)
  wire _1044_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16122" *)
  wire _1045_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16123" *)
  wire _1046_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16142" *)
  wire _1047_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16278" *)
  wire _1048_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16302" *)
  wire _1049_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16303" *)
  wire _1050_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16312" *)
  wire _1051_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16313" *)
  wire _1052_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18509" *)
  wire _1053_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:19941" *)
  wire _1054_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:2017" *)
  wire _1055_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:2018" *)
  wire _1056_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:2027" *)
  wire _1057_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:2028" *)
  wire _1058_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:2159" *)
  wire _1059_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:6884" *)
  wire _1060_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:8551" *)
  wire _1061_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:8816" *)
  wire _1062_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16276" *)
  wire _1063_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16277" *)
  wire _1064_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:2029" *)
  wire _1065_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:9348" *)
  wire _1066_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:10409" *)
  wire _1067_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:10410" *)
  wire _1068_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:11406" *)
  wire _1069_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:11419" *)
  wire _1070_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15961" *)
  wire _1071_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15961" *)
  wire _1072_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15963" *)
  wire _1073_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:12188" *)
  wire _1074_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15240" *)
  wire _1075_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15262" *)
  wire _1076_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16140" *)
  wire _1077_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:10245" *)
  wire _1078_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:10455" *)
  wire _1079_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:10455" *)
  wire _1080_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:10471" *)
  wire _1081_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:11330" *)
  wire _1082_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:11330" *)
  wire _1083_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:11405" *)
  wire _1084_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:14533" *)
  wire _1085_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:14552" *)
  wire _1086_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:14553" *)
  wire _1087_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:14555" *)
  wire _1088_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:14557" *)
  wire _1089_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:14558" *)
  wire _1090_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:14564" *)
  wire _1091_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15176" *)
  wire _1092_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15178" *)
  wire _1093_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15192" *)
  wire _1094_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15194" *)
  wire _1095_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15208" *)
  wire _1096_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15210" *)
  wire _1097_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15224" *)
  wire _1098_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15226" *)
  wire _1099_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15780" *)
  wire _1100_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15790" *)
  wire _1101_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15980" *)
  wire _1102_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16104" *)
  wire _1103_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16121" *)
  wire _1104_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16121" *)
  wire _1105_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16141" *)
  wire _1106_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16143" *)
  wire _1107_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16145" *)
  wire _1108_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16378" *)
  wire _1109_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16378" *)
  wire _1110_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16379" *)
  wire _1111_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:8807" *)
  wire _1112_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:9100" *)
  wire _1113_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:9100" *)
  wire _1114_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:9100" *)
  wire _1115_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:9656" *)
  wire _1116_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:9658" *)
  wire _1117_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:9669" *)
  wire _1118_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:9678" *)
  wire _1119_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:9733" *)
  wire _1120_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:9734" *)
  wire _1121_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:9735" *)
  wire _1122_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:10244" *)
  wire _1123_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:10256" *)
  wire _1124_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:10410" *)
  wire _1125_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:10410" *)
  wire _1126_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:11330" *)
  wire _1127_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:11391" *)
  wire _1128_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:11405" *)
  wire _1129_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:11405" *)
  wire _1130_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:11419" *)
  wire _1131_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:12179" *)
  wire _1132_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:12188" *)
  wire _1133_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:12194" *)
  wire _1134_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15042" *)
  wire _1135_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15063" *)
  wire [26:0] _1136_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15812" *)
  wire [1023:0] _1137_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15813" *)
  wire [1023:0] _1138_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15857" *)
  wire [255:0] _1139_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15869" *)
  wire [255:0] _1140_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15881" *)
  wire [255:0] _1141_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15893" *)
  wire [255:0] _1142_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15960" *)
  wire _1143_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15960" *)
  wire _1144_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15980" *)
  wire _1145_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15980" *)
  wire _1146_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15986" *)
  wire _1147_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16104" *)
  wire _1148_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16121" *)
  wire _1149_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1940" *)
  wire _1150_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:8506" *)
  wire _1151_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:8516" *)
  wire [30:0] _1152_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:8713" *)
  wire _1153_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:8728" *)
  wire _1154_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:9687" *)
  wire _1155_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:9743" *)
  wire _1156_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:10417" *)
  wire _1157_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:10417" *)
  wire _1158_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:14581" *)
  wire _1159_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:7446" *)
  wire _1160_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:7446" *)
  wire _1161_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:8728" *)
  wire _1162_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:9100" *)
  wire _1163_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:9100" *)
  wire _1164_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:9100" *)
  wire _1165_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16271" *)
  wire [127:0] _1166_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1989" *)
  wire [5:0] _1167_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:10224" *)
  wire [13:0] _1168_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:9608" *)
  wire [13:0] _1169_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:10247" *)
  wire [13:0] _1170_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:10247" *)
  wire [13:0] _1171_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:10440" *)
  wire _1172_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:11343" *)
  wire [12:0] _1173_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:12180" *)
  wire [11:0] _1174_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:12193" *)
  wire [11:0] _1175_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:12193" *)
  wire [11:0] _1176_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:14567" *)
  wire _1177_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:14570" *)
  wire _1178_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:14573" *)
  wire _1179_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:14576" *)
  wire _1180_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:14579" *)
  wire _1181_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:14582" *)
  wire _1182_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:14585" *)
  wire _1183_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:14588" *)
  wire _1184_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15180" *)
  wire [7:0] _1185_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15180" *)
  wire [7:0] _1186_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15180" *)
  wire [7:0] _1187_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15180" *)
  wire [7:0] _1188_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15196" *)
  wire [7:0] _1189_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15196" *)
  wire [7:0] _1190_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15196" *)
  wire [7:0] _1191_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15196" *)
  wire [7:0] _1192_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15212" *)
  wire [7:0] _1193_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15212" *)
  wire [7:0] _1194_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15212" *)
  wire [7:0] _1195_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15212" *)
  wire [7:0] _1196_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15228" *)
  wire [7:0] _1197_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15228" *)
  wire [7:0] _1198_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15228" *)
  wire [7:0] _1199_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15228" *)
  wire [7:0] _1200_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15967" *)
  wire [1023:0] _1201_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15967" *)
  wire [1023:0] _1202_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15967" *)
  wire [1023:0] _1203_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15967" *)
  wire [1023:0] _1204_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15967" *)
  wire [1023:0] _1205_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15967" *)
  wire [1023:0] _1206_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15987" *)
  wire [511:0] _1207_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15987" *)
  wire [511:0] _1208_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15987" *)
  wire [511:0] _1209_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15987" *)
  wire [511:0] _1210_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15987" *)
  wire [511:0] _1211_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15987" *)
  wire [511:0] _1212_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16027" *)
  wire [2047:0] _1213_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16043" *)
  wire [1023:0] _1214_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16043" *)
  wire [1023:0] _1215_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16043" *)
  wire [1023:0] _1216_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16059" *)
  wire [1023:0] _1217_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16059" *)
  wire [1023:0] _1218_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16059" *)
  wire [1023:0] _1219_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16075" *)
  wire [1023:0] _1220_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16075" *)
  wire [1023:0] _1221_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16075" *)
  wire [1023:0] _1222_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16107" *)
  wire [1023:0] _1223_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16107" *)
  wire [1023:0] _1224_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16124" *)
  wire [511:0] _1225_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16124" *)
  wire [511:0] _1226_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16304" *)
  wire [127:0] _1227_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16314" *)
  wire [63:0] _1228_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16371" *)
  wire [127:0] _1229_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18424" *)
  wire [127:0] _1230_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18484" *)
  wire [1023:0] _1231_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18496" *)
  wire [127:0] _1232_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18496" *)
  wire [127:0] _1233_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1999" *)
  wire [2:0] _1234_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:2019" *)
  wire [5:0] _1235_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:2030" *)
  wire [5:0] _1236_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:2030" *)
  wire [7:0] _1237_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:2043" *)
  wire [7:0] _1238_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:6725" *)
  wire [11:0] _1239_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:8539" *)
  wire [5:0] _1240_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:8809" *)
  wire [6:0] _1241_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:8809" *)
  wire [6:0] _1242_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:9089" *)
  wire _1243_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:9101" *)
  wire _1244_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:9369" *)
  wire [12:0] _1245_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:9369" *)
  wire [12:0] _1246_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:9529" *)
  wire [10:0] _1247_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:9608" *)
  wire [13:0] _1248_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:9631" *)
  wire [13:0] _1249_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:9631" *)
  wire [13:0] _1250_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:9659" *)
  wire [16:0] _1251_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:9659" *)
  wire [16:0] _1252_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:9659" *)
  wire [16:0] _1253_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:9659" *)
  wire [16:0] _1254_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:9736" *)
  wire _1255_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:9736" *)
  wire _1256_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:9736" *)
  wire _1257_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:9736" *)
  wire _1258_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:9742" *)
  wire _1259_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:905" *)
  reg [4:0] batch_cmp;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:906" *)
  wire [4:0] batch_cmp_w;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:907" *)
  reg [4:0] batch_cnt;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:908" *)
  wire [4:0] batch_cnt_w;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:909" *)
  reg [11:0] c_bias;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:910" *)
  wire [11:0] c_bias_add;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:911" *)
  reg [11:0] c_bias_d1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:912" *)
  wire c_bias_d1_reg_en;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:913" *)
  wire c_bias_reg_en;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:914" *)
  wire [11:0] c_bias_w;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:915" *)
  wire cbuf_reset;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:327" *)
  input [11:0] cdma2sc_dat_entries;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:328" *)
  input [11:0] cdma2sc_dat_slices;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:326" *)
  input cdma2sc_dat_updt;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:916" *)
  reg [3:0] conv_x_stride;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:917" *)
  wire [3:0] conv_x_stride_w;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:918" *)
  reg [3:0] conv_y_stride;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:919" *)
  wire [3:0] conv_y_stride_w;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:920" *)
  wire dat_conv_req_dummy;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:624" *)
  wire dat_dummy_l0_en;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:625" *)
  wire dat_dummy_l1_en;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:626" *)
  wire dat_dummy_l2_en;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:627" *)
  wire dat_dummy_l3_en;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:923" *)
  wire [11:0] dat_entry_avl_sub;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:929" *)
  reg [11:0] dat_entry_st;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:930" *)
  wire [12:0] dat_entry_st_inc;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:931" *)
  wire [11:0] dat_entry_st_inc_wrap;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:932" *)
  wire [11:0] dat_entry_st_w;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:933" *)
  wire dat_exec_valid;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:934" *)
  reg dat_exec_valid_d1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:935" *)
  reg dat_exec_valid_d2;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:936" *)
  wire dat_img_req_dummy;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:937" *)
  wire dat_img_req_skip;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:628" *)
  wire dat_l0_set;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:938" *)
  reg dat_l0c0_dummy;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:629" *)
  wire dat_l0c0_dummy_w;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:939" *)
  wire dat_l0c0_en;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:940" *)
  reg [511:0] dat_l0c0_hi;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:941" *)
  reg [511:0] dat_l0c0_lo;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:942" *)
  reg dat_l0c1_dummy;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:630" *)
  wire dat_l0c1_dummy_w;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:943" *)
  wire dat_l0c1_en;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:944" *)
  reg [511:0] dat_l0c1_hi;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:945" *)
  reg [511:0] dat_l0c1_lo;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:631" *)
  wire dat_l1_set;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:946" *)
  reg dat_l1c0_dummy;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:632" *)
  wire dat_l1c0_dummy_w;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:947" *)
  wire dat_l1c0_en;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:948" *)
  reg [511:0] dat_l1c0_hi;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:949" *)
  wire dat_l1c0_hi_en;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:950" *)
  reg [511:0] dat_l1c0_lo;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:951" *)
  reg dat_l1c1_dummy;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:633" *)
  wire dat_l1c1_dummy_w;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:952" *)
  wire dat_l1c1_en;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:953" *)
  reg [511:0] dat_l1c1_hi;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:954" *)
  wire dat_l1c1_hi_en;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:955" *)
  reg [511:0] dat_l1c1_lo;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:634" *)
  wire dat_l2_set;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:956" *)
  reg dat_l2c0_dummy;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:635" *)
  wire dat_l2c0_dummy_w;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:957" *)
  wire dat_l2c0_en;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:958" *)
  reg [511:0] dat_l2c0_hi;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:959" *)
  reg [511:0] dat_l2c0_lo;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:960" *)
  reg dat_l2c1_dummy;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:636" *)
  wire dat_l2c1_dummy_w;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:961" *)
  wire dat_l2c1_en;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:962" *)
  reg [511:0] dat_l2c1_hi;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:963" *)
  reg [511:0] dat_l2c1_lo;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:637" *)
  wire dat_l3_set;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:964" *)
  reg dat_l3c0_dummy;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:638" *)
  wire dat_l3c0_dummy_w;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:965" *)
  wire dat_l3c0_en;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:966" *)
  reg [511:0] dat_l3c0_hi;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:967" *)
  reg [511:0] dat_l3c0_lo;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:968" *)
  reg dat_l3c1_dummy;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:639" *)
  wire dat_l3c1_dummy_w;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:969" *)
  wire dat_l3c1_en;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:970" *)
  reg [511:0] dat_l3c1_hi;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:971" *)
  reg [511:0] dat_l3c1_lo;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:972" *)
  reg [1023:0] dat_out_bypass_data;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:640" *)
  wire [1023:0] dat_out_bypass_data_w;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:973" *)
  reg [127:0] dat_out_bypass_mask;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:641" *)
  wire [127:0] dat_out_bypass_mask_w;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:642" *)
  wire dat_out_bypass_p0_vld_w;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:643" *)
  wire dat_out_bypass_p1_vld_w;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:974" *)
  wire [1023:0] dat_out_data;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:975" *)
  reg [8:0] dat_out_flag;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:644" *)
  wire [8:0] dat_out_flag_l0;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:976" *)
  reg [8:0] dat_out_flag_l1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:977" *)
  reg [8:0] dat_out_flag_l2;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:978" *)
  reg [8:0] dat_out_flag_l3;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:979" *)
  reg [8:0] dat_out_flag_l4;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:980" *)
  reg [8:0] dat_out_flag_l5;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:645" *)
  wire [8:0] dat_out_flag_w;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:981" *)
  wire [127:0] dat_out_mask;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:982" *)
  reg dat_out_pvld;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:646" *)
  wire dat_out_pvld_l0;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:983" *)
  reg dat_out_pvld_l1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:984" *)
  reg dat_out_pvld_l2;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:985" *)
  reg dat_out_pvld_l3;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:986" *)
  reg dat_out_pvld_l4;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:987" *)
  reg dat_out_pvld_l5;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:647" *)
  wire dat_out_pvld_w;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:988" *)
  wire [1023:0] dat_out_wg_16b;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:989" *)
  wire [511:0] dat_out_wg_8b;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:990" *)
  wire [1023:0] dat_out_wg_data;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:991" *)
  wire [127:0] dat_out_wg_mask;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:992" *)
  wire [127:0] dat_out_wg_mask_fp16;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:993" *)
  wire [127:0] dat_out_wg_mask_int16;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:994" *)
  wire [63:0] dat_out_wg_mask_int8;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:995" *)
  reg dat_pipe_local_valid;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:996" *)
  wire dat_pipe_local_valid_w;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:648" *)
  wire dat_pipe_valid;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:997" *)
  reg dat_pipe_valid_d1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:998" *)
  reg dat_pipe_valid_d2;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:999" *)
  wire [1023:0] dat_pra_dat;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:649" *)
  wire [255:0] dat_pra_dat_ch0;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:650" *)
  wire [255:0] dat_pra_dat_ch1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:651" *)
  wire [255:0] dat_pra_dat_ch2;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:652" *)
  wire [255:0] dat_pra_dat_ch3;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:653" *)
  wire [11:0] dat_req_addr_last;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1000" *)
  wire [12:0] dat_req_addr_sum;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1001" *)
  wire [11:0] dat_req_addr_w;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1002" *)
  wire [11:0] dat_req_addr_wrap;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:654" *)
  wire [11:0] dat_req_base_d1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:655" *)
  wire [4:0] dat_req_batch_index;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1003" *)
  wire [7:0] dat_req_bytes;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1004" *)
  reg [7:0] dat_req_bytes_d1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1005" *)
  reg [7:0] dat_req_bytes_d2;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1006" *)
  reg dat_req_ch_end_d1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1007" *)
  reg dat_req_ch_end_d2;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1008" *)
  reg dat_req_ch_odd_d1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1009" *)
  reg dat_req_ch_odd_d2;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:656" *)
  wire dat_req_channel_end;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1010" *)
  reg [1:0] dat_req_cur_sub_h_d1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1011" *)
  reg [1:0] dat_req_cur_sub_h_d2;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1012" *)
  wire dat_req_dummy;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1013" *)
  reg dat_req_dummy_d1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1014" *)
  reg dat_req_dummy_d2;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:657" *)
  wire dat_req_exec_dummy;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:658" *)
  wire dat_req_exec_pvld;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:659" *)
  wire [1:0] dat_req_exec_sub_h;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1015" *)
  reg [8:0] dat_req_flag_d1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1016" *)
  reg [8:0] dat_req_flag_d2;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:660" *)
  wire [8:0] dat_req_flag_w;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:661" *)
  wire dat_req_layer_end;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:662" *)
  wire [7:0] dat_req_pipe_bytes;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:663" *)
  wire dat_req_pipe_ch_end;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:664" *)
  wire dat_req_pipe_ch_odd;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:665" *)
  wire [1:0] dat_req_pipe_cur_sub_h;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:666" *)
  wire dat_req_pipe_dummy;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:667" *)
  wire [8:0] dat_req_pipe_flag;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:668" *)
  wire [28:0] dat_req_pipe_pd;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:669" *)
  wire dat_req_pipe_pvld;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:670" *)
  wire dat_req_pipe_rls;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:671" *)
  wire dat_req_pipe_sub_c;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:672" *)
  wire [1:0] dat_req_pipe_sub_h;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:673" *)
  wire [1:0] dat_req_pipe_sub_w;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:674" *)
  wire dat_req_pipe_sub_w_st;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1017" *)
  reg dat_req_rls_d1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1018" *)
  reg dat_req_rls_d2;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1019" *)
  wire dat_req_skip;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:675" *)
  wire dat_req_stripe_end;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:676" *)
  wire dat_req_stripe_st;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1020" *)
  reg dat_req_sub_c_d1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1021" *)
  reg dat_req_sub_c_d2;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1022" *)
  wire dat_req_sub_c_w;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1023" *)
  reg [11:0] dat_req_sub_h_0_addr;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:677" *)
  wire dat_req_sub_h_0_addr_en;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1024" *)
  reg [11:0] dat_req_sub_h_1_addr;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:678" *)
  wire dat_req_sub_h_1_addr_en;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1025" *)
  reg [11:0] dat_req_sub_h_2_addr;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:679" *)
  wire dat_req_sub_h_2_addr_en;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1026" *)
  reg [11:0] dat_req_sub_h_3_addr;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:680" *)
  wire dat_req_sub_h_3_addr_en;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1027" *)
  reg [1:0] dat_req_sub_h_d1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1028" *)
  reg [1:0] dat_req_sub_h_d2;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1029" *)
  reg [1:0] dat_req_sub_w_d1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1030" *)
  reg [1:0] dat_req_sub_w_d2;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1031" *)
  reg dat_req_sub_w_st_d1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1032" *)
  reg dat_req_sub_w_st_d2;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:681" *)
  wire dat_req_sub_w_st_en;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1033" *)
  wire [1:0] dat_req_sub_w_w;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1034" *)
  wire dat_req_valid;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1035" *)
  reg dat_req_valid_d1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1036" *)
  wire dat_rls;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:682" *)
  wire [4:0] dat_rsp_batch_index;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:683" *)
  wire [7:0] dat_rsp_bytes;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:684" *)
  wire dat_rsp_ch_end;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:685" *)
  (* unused_bits = "0" *)
  wire dat_rsp_ch_odd;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:686" *)
  wire dat_rsp_channel_end;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1037" *)
  wire [1023:0] dat_rsp_conv;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1038" *)
  wire [1023:0] dat_rsp_conv_16b;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1039" *)
  wire [511:0] dat_rsp_conv_8b;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1040" *)
  wire [127:0] dat_rsp_cur_h_e2_mask_16b;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1041" *)
  wire [63:0] dat_rsp_cur_h_e2_mask_8b;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1042" *)
  wire [127:0] dat_rsp_cur_h_e4_mask_16b;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1043" *)
  wire [63:0] dat_rsp_cur_h_e4_mask_8b;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1044" *)
  wire [63:0] dat_rsp_cur_h_mask_p1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1045" *)
  wire [31:0] dat_rsp_cur_h_mask_p2;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1046" *)
  wire [31:0] dat_rsp_cur_h_mask_p3;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:687" *)
  wire [1:0] dat_rsp_cur_sub_h;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1047" *)
  wire [1023:0] dat_rsp_data_w;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:688" *)
  wire dat_rsp_exec_dummy;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:689" *)
  wire dat_rsp_exec_dummy_d0;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1048" *)
  reg dat_rsp_exec_dummy_d1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1049" *)
  reg dat_rsp_exec_dummy_d2;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1050" *)
  reg dat_rsp_exec_dummy_d3;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1051" *)
  reg dat_rsp_exec_dummy_d4;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1052" *)
  reg dat_rsp_exec_dummy_d5;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1053" *)
  reg dat_rsp_exec_dummy_d6;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:690" *)
  wire dat_rsp_exec_pvld;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:691" *)
  wire dat_rsp_exec_pvld_d0;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1054" *)
  reg dat_rsp_exec_pvld_d1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1055" *)
  reg dat_rsp_exec_pvld_d2;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1056" *)
  reg dat_rsp_exec_pvld_d3;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1057" *)
  reg dat_rsp_exec_pvld_d4;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1058" *)
  reg dat_rsp_exec_pvld_d5;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1059" *)
  reg dat_rsp_exec_pvld_d6;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:692" *)
  wire [1:0] dat_rsp_exec_sub_h;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:693" *)
  wire [1:0] dat_rsp_exec_sub_h_d0;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1060" *)
  reg [1:0] dat_rsp_exec_sub_h_d1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1061" *)
  reg [1:0] dat_rsp_exec_sub_h_d2;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1062" *)
  reg [1:0] dat_rsp_exec_sub_h_d3;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1063" *)
  reg [1:0] dat_rsp_exec_sub_h_d4;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1064" *)
  reg [1:0] dat_rsp_exec_sub_h_d5;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1065" *)
  reg [1:0] dat_rsp_exec_sub_h_d6;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:694" *)
  wire [8:0] dat_rsp_flag;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1066" *)
  wire [1023:0] dat_rsp_img;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1067" *)
  wire [1023:0] dat_rsp_img_16b;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1068" *)
  wire [511:0] dat_rsp_img_8b;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:695" *)
  wire dat_rsp_l0_block_end;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1069" *)
  wire dat_rsp_l0_ch_odd;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1070" *)
  wire [8:0] dat_rsp_l0_flag;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1071" *)
  wire dat_rsp_l0_pvld;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1072" *)
  wire [1023:0] dat_rsp_l0_sft;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1073" *)
  reg [511:0] dat_rsp_l0_sft_d1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1074" *)
  reg [255:0] dat_rsp_l0_sft_d2;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1075" *)
  reg [255:0] dat_rsp_l0_sft_d3;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1076" *)
  wire [2047:0] dat_rsp_l0_sft_in;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1077" *)
  wire dat_rsp_l0_stripe_end;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1078" *)
  wire dat_rsp_l0_sub_c;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1079" *)
  wire [511:0] dat_rsp_l0c0_hi;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1080" *)
  wire [511:0] dat_rsp_l0c0_lo;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1081" *)
  wire [511:0] dat_rsp_l0c1_hi;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1082" *)
  wire [511:0] dat_rsp_l0c1_lo;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:696" *)
  wire dat_rsp_l1_block_end;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1083" *)
  wire dat_rsp_l1_ch_odd;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1084" *)
  wire [8:0] dat_rsp_l1_flag;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1085" *)
  wire dat_rsp_l1_pvld;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1086" *)
  wire [511:0] dat_rsp_l1_sft;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1087" *)
  reg [255:0] dat_rsp_l1_sft_d2;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1088" *)
  reg [255:0] dat_rsp_l1_sft_d3;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1089" *)
  wire [1023:0] dat_rsp_l1_sft_in;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1090" *)
  wire dat_rsp_l1_stripe_end;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1091" *)
  wire dat_rsp_l1_sub_c;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1092" *)
  wire [511:0] dat_rsp_l1c0_hi;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1093" *)
  wire [511:0] dat_rsp_l1c0_lo;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1094" *)
  wire [511:0] dat_rsp_l1c1_hi;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1095" *)
  wire [511:0] dat_rsp_l1c1_lo;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:697" *)
  wire dat_rsp_l2_block_end;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1096" *)
  wire dat_rsp_l2_ch_odd;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1097" *)
  wire [8:0] dat_rsp_l2_flag;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1098" *)
  wire dat_rsp_l2_pvld;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1099" *)
  wire [255:0] dat_rsp_l2_sft;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1100" *)
  reg [255:0] dat_rsp_l2_sft_d3;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1101" *)
  wire [1023:0] dat_rsp_l2_sft_in;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1102" *)
  wire dat_rsp_l2_stripe_end;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1103" *)
  wire dat_rsp_l2_sub_c;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1104" *)
  wire [511:0] dat_rsp_l2c0_hi;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1105" *)
  wire [511:0] dat_rsp_l2c0_lo;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1106" *)
  wire [511:0] dat_rsp_l2c1_hi;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1107" *)
  wire [511:0] dat_rsp_l2c1_lo;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:698" *)
  wire dat_rsp_l3_block_end;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1108" *)
  wire dat_rsp_l3_ch_odd;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1109" *)
  wire [8:0] dat_rsp_l3_flag;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1110" *)
  wire dat_rsp_l3_pvld;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1111" *)
  wire [255:0] dat_rsp_l3_sft;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1112" *)
  wire [1023:0] dat_rsp_l3_sft_in;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1113" *)
  wire dat_rsp_l3_stripe_end;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1114" *)
  wire dat_rsp_l3_sub_c;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1115" *)
  wire [511:0] dat_rsp_l3c0_hi;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1116" *)
  wire [511:0] dat_rsp_l3c0_lo;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1117" *)
  wire [511:0] dat_rsp_l3c1_hi;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1118" *)
  wire [511:0] dat_rsp_l3c1_lo;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:699" *)
  wire dat_rsp_layer_end;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1119" *)
  wire [127:0] dat_rsp_mask_16b;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1120" *)
  wire [63:0] dat_rsp_mask_8b;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1121" *)
  wire [127:0] dat_rsp_mask_val_fp16;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1122" *)
  wire [127:0] dat_rsp_mask_val_int16;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1123" *)
  wire [63:0] dat_rsp_mask_val_int8;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1124" *)
  wire [127:0] dat_rsp_mask_w;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1125" *)
  wire [127:0] dat_rsp_ori_mask;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1126" *)
  wire dat_rsp_p0_vld_w;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1127" *)
  wire dat_rsp_p1_vld_w;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1128" *)
  wire [511:0] dat_rsp_pad_value;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1129" *)
  (* unused_bits = "3 6" *)
  wire [26:0] dat_rsp_pd;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:700" *)
  wire [26:0] dat_rsp_pd_d0;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1130" *)
  reg [26:0] dat_rsp_pd_d1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1131" *)
  reg [26:0] dat_rsp_pd_d2;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1132" *)
  reg [26:0] dat_rsp_pd_d3;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1133" *)
  reg [26:0] dat_rsp_pd_d4;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:701" *)
  wire [7:0] dat_rsp_pipe_bytes;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:702" *)
  wire dat_rsp_pipe_ch_end;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:703" *)
  wire dat_rsp_pipe_ch_odd;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:704" *)
  wire [1:0] dat_rsp_pipe_cur_sub_h;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:705" *)
  wire dat_rsp_pipe_dummy;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:706" *)
  wire [8:0] dat_rsp_pipe_flag;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:707" *)
  wire [28:0] dat_rsp_pipe_pd;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:708" *)
  wire [28:0] dat_rsp_pipe_pd_d0;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1134" *)
  reg [28:0] dat_rsp_pipe_pd_d1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1135" *)
  reg [28:0] dat_rsp_pipe_pd_d2;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1136" *)
  reg [28:0] dat_rsp_pipe_pd_d3;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1137" *)
  reg [28:0] dat_rsp_pipe_pd_d4;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1138" *)
  reg [28:0] dat_rsp_pipe_pd_d5;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1139" *)
  reg [28:0] dat_rsp_pipe_pd_d6;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:709" *)
  wire dat_rsp_pipe_pvld;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:710" *)
  wire dat_rsp_pipe_pvld_d0;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1140" *)
  reg dat_rsp_pipe_pvld_d1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1141" *)
  reg dat_rsp_pipe_pvld_d2;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1142" *)
  reg dat_rsp_pipe_pvld_d3;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1143" *)
  reg dat_rsp_pipe_pvld_d4;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1144" *)
  reg dat_rsp_pipe_pvld_d5;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1145" *)
  reg dat_rsp_pipe_pvld_d6;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:711" *)
  wire dat_rsp_pipe_rls;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:712" *)
  wire dat_rsp_pipe_sub_c;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:713" *)
  wire [1:0] dat_rsp_pipe_sub_h;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:714" *)
  wire [1:0] dat_rsp_pipe_sub_w;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:715" *)
  wire dat_rsp_pipe_sub_w_st;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1146" *)
  wire dat_rsp_pra_en;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1147" *)
  wire [3:0] dat_rsp_pra_en_d1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1148" *)
  wire dat_rsp_pvld;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:716" *)
  wire dat_rsp_pvld_d0;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1149" *)
  reg dat_rsp_pvld_d1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1150" *)
  reg dat_rsp_pvld_d2;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1151" *)
  reg dat_rsp_pvld_d3;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1152" *)
  reg dat_rsp_pvld_d4;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:717" *)
  wire dat_rsp_rls;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1153" *)
  wire dat_rsp_sft_hi_d1_en;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1154" *)
  wire dat_rsp_sft_hi_d2_en;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1155" *)
  wire dat_rsp_sft_hi_d3_en;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1156" *)
  wire dat_rsp_sft_lo_d1_en;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1157" *)
  wire dat_rsp_sft_lo_d2_en;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1158" *)
  wire dat_rsp_sft_lo_d3_en;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:718" *)
  wire dat_rsp_stripe_end;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:719" *)
  wire dat_rsp_stripe_st;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:720" *)
  wire dat_rsp_sub_c;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:721" *)
  (* unused_bits = "1" *)
  wire [1:0] dat_rsp_sub_h;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:722" *)
  wire [1:0] dat_rsp_sub_w;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1159" *)
  wire [1023:0] dat_rsp_wg;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1160" *)
  wire [255:0] dat_rsp_wg_ch0;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1161" *)
  reg [255:0] dat_rsp_wg_ch0_d1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1162" *)
  wire [255:0] dat_rsp_wg_ch1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1163" *)
  reg [255:0] dat_rsp_wg_ch1_d1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1164" *)
  wire [255:0] dat_rsp_wg_ch2;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1165" *)
  reg [255:0] dat_rsp_wg_ch2_d1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1166" *)
  wire [255:0] dat_rsp_wg_ch3;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1167" *)
  reg [255:0] dat_rsp_wg_ch3_d1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1168" *)
  wire [1023:0] dat_rsp_wg_lb;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1169" *)
  wire [1023:0] dat_rsp_wg_lt;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1170" *)
  wire [1023:0] dat_rsp_wg_rb;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1171" *)
  wire [1023:0] dat_rsp_wg_rt;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1172" *)
  wire dat_rsp_wg_sel_16b;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1173" *)
  wire dat_rsp_wg_sel_8b_hi;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1174" *)
  wire dat_rsp_wg_sel_8b_lo;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1175" *)
  wire dat_rsp_wg_sel_lb;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1176" *)
  wire dat_rsp_wg_sel_lt;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1177" *)
  wire dat_rsp_wg_sel_rb;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1178" *)
  wire dat_rsp_wg_sel_rt;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1183" *)
  wire [2303:0] dat_wg;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:723" *)
  wire [255:0] dat_wg_16b_ch0;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:724" *)
  wire [255:0] dat_wg_16b_ch1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:725" *)
  wire [255:0] dat_wg_16b_ch2;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:726" *)
  wire [255:0] dat_wg_16b_ch3;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:727" *)
  wire [255:0] dat_wg_8b_ch0;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:728" *)
  wire [255:0] dat_wg_8b_ch1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:729" *)
  wire [255:0] dat_wg_8b_ch2;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:730" *)
  wire [255:0] dat_wg_8b_ch3;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:731" *)
  wire [255:0] dat_wg_8b_ch4;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:732" *)
  wire [255:0] dat_wg_8b_ch5;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:733" *)
  wire [255:0] dat_wg_8b_ch6;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:734" *)
  wire [255:0] dat_wg_8b_ch7;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:735" *)
  wire dat_wg_adv;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:736" *)
  wire dat_wg_req_dummy;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1184" *)
  wire dat_wg_req_skip;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1185" *)
  reg [3:0] data_bank;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1186" *)
  wire [3:0] data_bank_w;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1187" *)
  reg [5:0] data_batch;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1188" *)
  wire [5:0] data_batch_w;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1189" *)
  reg [10:0] datain_c_cnt;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1190" *)
  wire [10:0] datain_c_cnt_inc;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1191" *)
  wire datain_c_cnt_reg_en;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1192" *)
  wire [10:0] datain_c_cnt_w;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1193" *)
  reg [10:0] datain_channel_cmp;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1194" *)
  wire [10:0] datain_channel_cmp_w;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1195" *)
  reg [13:0] datain_h_cnt;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1196" *)
  wire [13:0] datain_h_cnt_inc;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1197" *)
  wire datain_h_cnt_reg_en;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1198" *)
  wire [13:0] datain_h_cnt_st;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1199" *)
  wire [13:0] datain_h_cnt_w;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1200" *)
  wire [13:0] datain_h_cur;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1201" *)
  reg [13:0] datain_h_ori;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1202" *)
  wire datain_h_ori_reg_en;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1203" *)
  reg [12:0] datain_height_cmp;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1204" *)
  wire [12:0] datain_height_cmp_w;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1205" *)
  reg [13:0] datain_w_cnt;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1206" *)
  wire [13:0] datain_w_cnt_inc;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1207" *)
  wire datain_w_cnt_reg_en;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1208" *)
  wire [13:0] datain_w_cnt_st;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1209" *)
  wire [13:0] datain_w_cnt_w;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1210" *)
  wire [13:0] datain_w_cur;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1211" *)
  reg [13:0] datain_w_ori;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1212" *)
  wire datain_w_ori_reg_en;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1213" *)
  reg [13:0] datain_width;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1214" *)
  reg [12:0] datain_width_cmp;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1215" *)
  wire [12:0] datain_width_cmp_w;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1216" *)
  wire [13:0] datain_width_w;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:737" *)
  wire [2:0] dataout_w_add;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1217" *)
  reg [12:0] dataout_w_cnt;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1218" *)
  wire [12:0] dataout_w_cnt_inc;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1219" *)
  wire dataout_w_cnt_reg_en;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1220" *)
  wire [12:0] dataout_w_cnt_w;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1221" *)
  wire [12:0] dataout_w_init;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1222" *)
  reg [12:0] dataout_w_ori;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1223" *)
  wire dataout_w_ori_reg_en;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1224" *)
  reg [12:0] dataout_width_cmp;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1225" *)
  wire [12:0] dataout_width_cmp_w;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:867" *)
  wire dl_block_end;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:868" *)
  wire dl_channel_end;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:869" *)
  wire [6:0] dl_channel_size;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:870" *)
  wire [1:0] dl_cur_sub_h;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:871" *)
  wire dl_dat_release;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:872" *)
  wire dl_group_end;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:873" *)
  wire [4:0] dl_h_offset;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1226" *)
  wire [9:0] dl_h_offset_ext;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:874" *)
  wire [30:0] dl_in_pd;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:875" *)
  wire [30:0] dl_in_pd_d0;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1227" *)
  reg [30:0] dl_in_pd_d1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1228" *)
  reg [30:0] dl_in_pd_d2;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1229" *)
  reg [30:0] dl_in_pd_d3;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1230" *)
  reg [30:0] dl_in_pd_d4;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1231" *)
  reg [30:0] dl_in_pd_d5;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:876" *)
  wire dl_in_pvld;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:877" *)
  wire dl_in_pvld_d0;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1232" *)
  reg dl_in_pvld_d1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1233" *)
  reg dl_in_pvld_d2;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1234" *)
  reg dl_in_pvld_d3;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1235" *)
  reg dl_in_pvld_d4;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1236" *)
  reg dl_in_pvld_d5;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:878" *)
  wire dl_layer_end;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1237" *)
  reg [7:0] dl_out_data0;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1238" *)
  reg [7:0] dl_out_data1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1239" *)
  reg [7:0] dl_out_data10;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1240" *)
  reg [7:0] dl_out_data100;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1241" *)
  reg [7:0] dl_out_data101;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1242" *)
  reg [7:0] dl_out_data102;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1243" *)
  reg [7:0] dl_out_data103;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1244" *)
  reg [7:0] dl_out_data104;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1245" *)
  reg [7:0] dl_out_data105;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1246" *)
  reg [7:0] dl_out_data106;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1247" *)
  reg [7:0] dl_out_data107;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1248" *)
  reg [7:0] dl_out_data108;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1249" *)
  reg [7:0] dl_out_data109;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1250" *)
  reg [7:0] dl_out_data11;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1251" *)
  reg [7:0] dl_out_data110;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1252" *)
  reg [7:0] dl_out_data111;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1253" *)
  reg [7:0] dl_out_data112;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1254" *)
  reg [7:0] dl_out_data113;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1255" *)
  reg [7:0] dl_out_data114;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1256" *)
  reg [7:0] dl_out_data115;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1257" *)
  reg [7:0] dl_out_data116;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1258" *)
  reg [7:0] dl_out_data117;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1259" *)
  reg [7:0] dl_out_data118;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1260" *)
  reg [7:0] dl_out_data119;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1261" *)
  reg [7:0] dl_out_data12;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1262" *)
  reg [7:0] dl_out_data120;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1263" *)
  reg [7:0] dl_out_data121;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1264" *)
  reg [7:0] dl_out_data122;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1265" *)
  reg [7:0] dl_out_data123;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1266" *)
  reg [7:0] dl_out_data124;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1267" *)
  reg [7:0] dl_out_data125;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1268" *)
  reg [7:0] dl_out_data126;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1269" *)
  reg [7:0] dl_out_data127;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1270" *)
  reg [7:0] dl_out_data13;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1271" *)
  reg [7:0] dl_out_data14;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1272" *)
  reg [7:0] dl_out_data15;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1273" *)
  reg [7:0] dl_out_data16;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1274" *)
  reg [7:0] dl_out_data17;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1275" *)
  reg [7:0] dl_out_data18;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1276" *)
  reg [7:0] dl_out_data19;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1277" *)
  reg [7:0] dl_out_data2;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1278" *)
  reg [7:0] dl_out_data20;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1279" *)
  reg [7:0] dl_out_data21;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1280" *)
  reg [7:0] dl_out_data22;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1281" *)
  reg [7:0] dl_out_data23;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1282" *)
  reg [7:0] dl_out_data24;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1283" *)
  reg [7:0] dl_out_data25;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1284" *)
  reg [7:0] dl_out_data26;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1285" *)
  reg [7:0] dl_out_data27;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1286" *)
  reg [7:0] dl_out_data28;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1287" *)
  reg [7:0] dl_out_data29;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1288" *)
  reg [7:0] dl_out_data3;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1289" *)
  reg [7:0] dl_out_data30;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1290" *)
  reg [7:0] dl_out_data31;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1291" *)
  reg [7:0] dl_out_data32;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1292" *)
  reg [7:0] dl_out_data33;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1293" *)
  reg [7:0] dl_out_data34;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1294" *)
  reg [7:0] dl_out_data35;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1295" *)
  reg [7:0] dl_out_data36;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1296" *)
  reg [7:0] dl_out_data37;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1297" *)
  reg [7:0] dl_out_data38;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1298" *)
  reg [7:0] dl_out_data39;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1299" *)
  reg [7:0] dl_out_data4;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1300" *)
  reg [7:0] dl_out_data40;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1301" *)
  reg [7:0] dl_out_data41;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1302" *)
  reg [7:0] dl_out_data42;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1303" *)
  reg [7:0] dl_out_data43;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1304" *)
  reg [7:0] dl_out_data44;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1305" *)
  reg [7:0] dl_out_data45;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1306" *)
  reg [7:0] dl_out_data46;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1307" *)
  reg [7:0] dl_out_data47;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1308" *)
  reg [7:0] dl_out_data48;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1309" *)
  reg [7:0] dl_out_data49;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1310" *)
  reg [7:0] dl_out_data5;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1311" *)
  reg [7:0] dl_out_data50;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1312" *)
  reg [7:0] dl_out_data51;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1313" *)
  reg [7:0] dl_out_data52;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1314" *)
  reg [7:0] dl_out_data53;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1315" *)
  reg [7:0] dl_out_data54;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1316" *)
  reg [7:0] dl_out_data55;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1317" *)
  reg [7:0] dl_out_data56;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1318" *)
  reg [7:0] dl_out_data57;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1319" *)
  reg [7:0] dl_out_data58;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1320" *)
  reg [7:0] dl_out_data59;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1321" *)
  reg [7:0] dl_out_data6;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1322" *)
  reg [7:0] dl_out_data60;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1323" *)
  reg [7:0] dl_out_data61;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1324" *)
  reg [7:0] dl_out_data62;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1325" *)
  reg [7:0] dl_out_data63;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1326" *)
  reg [7:0] dl_out_data64;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1327" *)
  reg [7:0] dl_out_data65;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1328" *)
  reg [7:0] dl_out_data66;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1329" *)
  reg [7:0] dl_out_data67;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1330" *)
  reg [7:0] dl_out_data68;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1331" *)
  reg [7:0] dl_out_data69;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1332" *)
  reg [7:0] dl_out_data7;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1333" *)
  reg [7:0] dl_out_data70;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1334" *)
  reg [7:0] dl_out_data71;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1335" *)
  reg [7:0] dl_out_data72;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1336" *)
  reg [7:0] dl_out_data73;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1337" *)
  reg [7:0] dl_out_data74;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1338" *)
  reg [7:0] dl_out_data75;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1339" *)
  reg [7:0] dl_out_data76;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1340" *)
  reg [7:0] dl_out_data77;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1341" *)
  reg [7:0] dl_out_data78;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1342" *)
  reg [7:0] dl_out_data79;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1343" *)
  reg [7:0] dl_out_data8;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1344" *)
  reg [7:0] dl_out_data80;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1345" *)
  reg [7:0] dl_out_data81;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1346" *)
  reg [7:0] dl_out_data82;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1347" *)
  reg [7:0] dl_out_data83;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1348" *)
  reg [7:0] dl_out_data84;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1349" *)
  reg [7:0] dl_out_data85;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1350" *)
  reg [7:0] dl_out_data86;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1351" *)
  reg [7:0] dl_out_data87;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1352" *)
  reg [7:0] dl_out_data88;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1353" *)
  reg [7:0] dl_out_data89;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1354" *)
  reg [7:0] dl_out_data9;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1355" *)
  reg [7:0] dl_out_data90;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1356" *)
  reg [7:0] dl_out_data91;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1357" *)
  reg [7:0] dl_out_data92;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1358" *)
  reg [7:0] dl_out_data93;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1359" *)
  reg [7:0] dl_out_data94;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1360" *)
  reg [7:0] dl_out_data95;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1361" *)
  reg [7:0] dl_out_data96;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1362" *)
  reg [7:0] dl_out_data97;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1363" *)
  reg [7:0] dl_out_data98;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1364" *)
  reg [7:0] dl_out_data99;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1365" *)
  reg [8:0] dl_out_flag;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1366" *)
  reg [127:0] dl_out_mask;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1367" *)
  reg dl_out_pvld;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1368" *)
  wire dl_out_pvld_d1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1369" *)
  wire [30:0] dl_pd;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:879" *)
  wire [30:0] dl_pd_d0;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1370" *)
  reg [30:0] dl_pd_d1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1371" *)
  reg [30:0] dl_pd_d2;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1372" *)
  reg [30:0] dl_pd_d3;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1373" *)
  reg [30:0] dl_pd_d4;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1374" *)
  wire dl_pvld;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:880" *)
  wire dl_pvld_d0;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1375" *)
  reg dl_pvld_d1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1376" *)
  reg dl_pvld_d2;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1377" *)
  reg dl_pvld_d3;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1378" *)
  reg dl_pvld_d4;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:881" *)
  wire [6:0] dl_stripe_length;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:882" *)
  wire [4:0] dl_w_offset;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1379" *)
  wire [9:0] dl_w_offset_ext;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1380" *)
  reg [11:0] entries;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1381" *)
  reg [11:0] entries_batch;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1382" *)
  wire [11:0] entries_batch_w;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1383" *)
  reg [11:0] entries_cmp;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1384" *)
  wire [11:0] entries_single_w;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1385" *)
  wire [11:0] entries_w;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1386" *)
  reg [11:0] h_bias_0_d1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1387" *)
  reg [11:0] h_bias_0_stride;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1388" *)
  wire [11:0] h_bias_0_stride_w;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1389" *)
  wire [11:0] h_bias_0_w;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1390" *)
  reg [11:0] h_bias_1_d1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1391" *)
  reg [11:0] h_bias_1_stride;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1392" *)
  wire [11:0] h_bias_1_stride_w;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1393" *)
  wire [11:0] h_bias_1_w;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1394" *)
  reg [11:0] h_bias_2_d1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1395" *)
  reg [11:0] h_bias_2_stride;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1396" *)
  wire [11:0] h_bias_2_w;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1397" *)
  reg [11:0] h_bias_3_d1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1398" *)
  reg [11:0] h_bias_3_stride;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1399" *)
  wire [11:0] h_bias_3_w;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1400" *)
  wire [11:0] h_bias_d1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:883" *)
  wire [1:0] h_bias_reg_en;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1401" *)
  reg [11:0] h_offset_slice;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1402" *)
  wire [11:0] h_offset_slice_w;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1403" *)
  wire is_batch_end;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1404" *)
  wire is_conv;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1406" *)
  wire is_dat_entry_st_wrap;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1407" *)
  wire is_dat_req_addr_wrap;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1408" *)
  wire is_fp16;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1409" *)
  reg [1:0] is_fp16_d1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1410" *)
  wire is_img;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1411" *)
  reg [33:0] is_img_d1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1412" *)
  wire is_int8;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1413" *)
  reg [22:0] is_int8_d1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1414" *)
  wire is_last_channel;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1415" *)
  wire is_pixel;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1417" *)
  wire is_sg_done;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1418" *)
  wire is_sg_idle;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1421" *)
  wire is_stripe_end;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1422" *)
  wire is_stripe_equal;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1423" *)
  wire is_sub_h_end;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1424" *)
  wire is_w_end;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1425" *)
  wire is_w_end_ahead;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1426" *)
  wire is_winograd;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1427" *)
  reg [21:0] is_winograd_d1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1428" *)
  reg [11:0] last_entries;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1429" *)
  reg [11:0] last_slices;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1430" *)
  wire layer_st;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1431" *)
  reg layer_st_d1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1432" *)
  wire mon_batch_cnt_w;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1433" *)
  wire mon_c_bias_w;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:884" *)
  (* unused_bits = "0 1 2 3" *)
  wire [3:0] mon_dat_out_pra_vld;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:885" *)
  (* unused_bits = "0 1 2 3" *)
  wire [3:0] mon_dat_rsp_pra_rdy;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1447" *)
  wire mon_datain_w_cnt_inc;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1452" *)
  wire mon_entries_w;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1458" *)
  wire [1:0] mon_h_bias_3_w;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1460" *)
  wire mon_pixel_w_cnt_w;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1461" *)
  wire [1:0] mon_pixel_x_init_w;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1468" *)
  wire [1:0] mon_slice_left_w;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1470" *)
  (* unused_bits = "0 1 2" *)
  wire [2:0] mon_sub_h_total_w;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:319" *)
  input nvdla_core_clk;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:598" *)
  input nvdla_core_ng_clk;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:320" *)
  input nvdla_core_rstn;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:599" *)
  input nvdla_wg_clk;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1471" *)
  reg [15:0] pad_value;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1472" *)
  wire pixel_ch_ori_reg_en;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1473" *)
  reg [11:0] pixel_ch_stride;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1474" *)
  wire [11:0] pixel_ch_stride_w;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:886" *)
  wire pixel_force_clr;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1475" *)
  reg pixel_force_clr_d1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:887" *)
  wire pixel_force_fetch;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1476" *)
  reg pixel_force_fetch_d1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1477" *)
  reg pixel_req_ch_odd;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:888" *)
  wire pixel_req_ch_odd_en;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1478" *)
  reg pixel_req_ch_odd_ori;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:889" *)
  wire pixel_req_ch_odd_ori_en;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1479" *)
  wire pixel_req_ch_odd_w;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1480" *)
  reg [15:0] pixel_w_ch_ori;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1481" *)
  reg [15:0] pixel_w_cnt;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1482" *)
  wire pixel_w_cnt_reg_en;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1483" *)
  wire [15:0] pixel_w_cnt_w;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:890" *)
  wire [9:0] pixel_w_cur;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1484" *)
  reg [15:0] pixel_w_ori;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1485" *)
  wire pixel_w_ori_reg_en;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1486" *)
  reg [6:0] pixel_x_add;
  wire [6:0] pixel_x_add_w;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1488" *)
  reg [6:0] pixel_x_byte_stride;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1489" *)
  wire [6:0] pixel_x_byte_stride_w;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1490" *)
  wire [6:0] pixel_x_cnt_add;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1491" *)
  reg [5:0] pixel_x_init;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1492" *)
  reg [6:0] pixel_x_init_offset;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1493" *)
  wire [6:0] pixel_x_init_offset_w;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1494" *)
  wire [5:0] pixel_x_init_w;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1495" *)
  reg pixel_x_stride_odd;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1496" *)
  wire [5:0] pixel_x_stride_w;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1497" *)
  reg [7:0] pra_precision;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:891" *)
  wire [1:0] pra_precision_0;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:892" *)
  wire [1:0] pra_precision_1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:893" *)
  wire [1:0] pra_precision_2;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:894" *)
  wire [1:0] pra_precision_3;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1498" *)
  reg [7:0] pra_truncate;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:895" *)
  wire [1:0] pra_truncate_0;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:896" *)
  wire [1:0] pra_truncate_1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:897" *)
  wire [1:0] pra_truncate_2;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:898" *)
  wire [1:0] pra_truncate_3;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1499" *)
  wire [1:0] pra_truncate_w;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:602" *)
  input [4:0] reg2dp_batches;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:601" *)
  input reg2dp_conv_mode;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:614" *)
  input [2:0] reg2dp_conv_x_stride_ext;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:615" *)
  input [2:0] reg2dp_conv_y_stride_ext;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:621" *)
  input [3:0] reg2dp_data_bank;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:606" *)
  input [12:0] reg2dp_datain_channel_ext;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:604" *)
  input reg2dp_datain_format;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:607" *)
  input [12:0] reg2dp_datain_height_ext;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:608" *)
  input [12:0] reg2dp_datain_width_ext;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:612" *)
  input [12:0] reg2dp_dataout_width;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:611" *)
  input [11:0] reg2dp_entries;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:600" *)
  input reg2dp_op_en;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:618" *)
  input [4:0] reg2dp_pad_left;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:619" *)
  input [4:0] reg2dp_pad_top;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:620" *)
  input [15:0] reg2dp_pad_value;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:622" *)
  input [1:0] reg2dp_pra_truncate;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:603" *)
  input [1:0] reg2dp_proc_precision;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:613" *)
  input [11:0] reg2dp_rls_slices;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:605" *)
  input reg2dp_skip_data_rls;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:610" *)
  input [12:0] reg2dp_weight_channel_ext;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:616" *)
  input [4:0] reg2dp_x_dilation_ext;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:617" *)
  input [4:0] reg2dp_y_dilation_ext;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:609" *)
  input [1:0] reg2dp_y_extension;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1500" *)
  wire reuse_rls;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1501" *)
  reg [11:0] rls_entries;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1502" *)
  reg [11:0] rls_slices;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1503" *)
  wire [11:0] rls_slices_w;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1504" *)
  reg [7:0] rsp_sft_cnt_l0;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1505" *)
  wire rsp_sft_cnt_l0_en;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1506" *)
  wire [7:0] rsp_sft_cnt_l0_inc;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1507" *)
  reg [7:0] rsp_sft_cnt_l0_ori;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1508" *)
  wire rsp_sft_cnt_l0_ori_en;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:899" *)
  wire [7:0] rsp_sft_cnt_l0_sub;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1509" *)
  wire [7:0] rsp_sft_cnt_l0_w;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1510" *)
  reg [7:0] rsp_sft_cnt_l1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1511" *)
  wire rsp_sft_cnt_l1_en;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1512" *)
  wire [7:0] rsp_sft_cnt_l1_inc;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1513" *)
  reg [7:0] rsp_sft_cnt_l1_ori;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1514" *)
  wire rsp_sft_cnt_l1_ori_en;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:900" *)
  wire [7:0] rsp_sft_cnt_l1_sub;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1515" *)
  wire [7:0] rsp_sft_cnt_l1_w;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1516" *)
  reg [7:0] rsp_sft_cnt_l2;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1517" *)
  wire rsp_sft_cnt_l2_en;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1518" *)
  wire [7:0] rsp_sft_cnt_l2_inc;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1519" *)
  reg [7:0] rsp_sft_cnt_l2_ori;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1520" *)
  wire rsp_sft_cnt_l2_ori_en;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:901" *)
  wire [7:0] rsp_sft_cnt_l2_sub;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1521" *)
  wire [7:0] rsp_sft_cnt_l2_w;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1522" *)
  reg [7:0] rsp_sft_cnt_l3;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1523" *)
  wire rsp_sft_cnt_l3_en;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1524" *)
  wire [7:0] rsp_sft_cnt_l3_inc;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1525" *)
  reg [7:0] rsp_sft_cnt_l3_ori;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1526" *)
  wire rsp_sft_cnt_l3_ori_en;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:902" *)
  wire [7:0] rsp_sft_cnt_l3_sub;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1527" *)
  wire [7:0] rsp_sft_cnt_l3_w;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1528" *)
  wire rsp_sft_l1_sel_1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1529" *)
  wire rsp_sft_l1_sel_2;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1530" *)
  wire rsp_sft_l1_sel_3;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1531" *)
  wire rsp_sft_l2_sel_1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1532" *)
  wire rsp_sft_l2_sel_2;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1533" *)
  wire rsp_sft_l2_sel_3;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1534" *)
  wire rsp_sft_l3_sel_1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1535" *)
  wire rsp_sft_l3_sel_2;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1536" *)
  wire rsp_sft_l3_sel_3;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:333" *)
  output [11:0] sc2buf_dat_rd_addr;
  reg [11:0] sc2buf_dat_rd_addr;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:335" *)
  input [1023:0] sc2buf_dat_rd_data;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:332" *)
  output sc2buf_dat_rd_en;
  reg sc2buf_dat_rd_en;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1539" *)
  wire sc2buf_dat_rd_en_w;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:334" *)
  input sc2buf_dat_rd_valid;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:330" *)
  output [11:0] sc2cdma_dat_entries;
  reg [11:0] sc2cdma_dat_entries;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1541" *)
  wire [11:0] sc2cdma_dat_entries_w;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:325" *)
  input sc2cdma_dat_pending_req;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:331" *)
  output [11:0] sc2cdma_dat_slices;
  reg [11:0] sc2cdma_dat_slices;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1543" *)
  wire [11:0] sc2cdma_dat_slices_w;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:329" *)
  output sc2cdma_dat_updt;
  reg sc2cdma_dat_updt;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:338" *)
  output [7:0] sc2mac_dat_a_data0;
  reg [7:0] sc2mac_dat_a_data0;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:339" *)
  output [7:0] sc2mac_dat_a_data1;
  reg [7:0] sc2mac_dat_a_data1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:348" *)
  output [7:0] sc2mac_dat_a_data10;
  reg [7:0] sc2mac_dat_a_data10;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:438" *)
  output [7:0] sc2mac_dat_a_data100;
  reg [7:0] sc2mac_dat_a_data100;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:439" *)
  output [7:0] sc2mac_dat_a_data101;
  reg [7:0] sc2mac_dat_a_data101;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:440" *)
  output [7:0] sc2mac_dat_a_data102;
  reg [7:0] sc2mac_dat_a_data102;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:441" *)
  output [7:0] sc2mac_dat_a_data103;
  reg [7:0] sc2mac_dat_a_data103;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:442" *)
  output [7:0] sc2mac_dat_a_data104;
  reg [7:0] sc2mac_dat_a_data104;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:443" *)
  output [7:0] sc2mac_dat_a_data105;
  reg [7:0] sc2mac_dat_a_data105;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:444" *)
  output [7:0] sc2mac_dat_a_data106;
  reg [7:0] sc2mac_dat_a_data106;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:445" *)
  output [7:0] sc2mac_dat_a_data107;
  reg [7:0] sc2mac_dat_a_data107;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:446" *)
  output [7:0] sc2mac_dat_a_data108;
  reg [7:0] sc2mac_dat_a_data108;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:447" *)
  output [7:0] sc2mac_dat_a_data109;
  reg [7:0] sc2mac_dat_a_data109;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:349" *)
  output [7:0] sc2mac_dat_a_data11;
  reg [7:0] sc2mac_dat_a_data11;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:448" *)
  output [7:0] sc2mac_dat_a_data110;
  reg [7:0] sc2mac_dat_a_data110;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:449" *)
  output [7:0] sc2mac_dat_a_data111;
  reg [7:0] sc2mac_dat_a_data111;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:450" *)
  output [7:0] sc2mac_dat_a_data112;
  reg [7:0] sc2mac_dat_a_data112;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:451" *)
  output [7:0] sc2mac_dat_a_data113;
  reg [7:0] sc2mac_dat_a_data113;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:452" *)
  output [7:0] sc2mac_dat_a_data114;
  reg [7:0] sc2mac_dat_a_data114;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:453" *)
  output [7:0] sc2mac_dat_a_data115;
  reg [7:0] sc2mac_dat_a_data115;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:454" *)
  output [7:0] sc2mac_dat_a_data116;
  reg [7:0] sc2mac_dat_a_data116;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:455" *)
  output [7:0] sc2mac_dat_a_data117;
  reg [7:0] sc2mac_dat_a_data117;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:456" *)
  output [7:0] sc2mac_dat_a_data118;
  reg [7:0] sc2mac_dat_a_data118;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:457" *)
  output [7:0] sc2mac_dat_a_data119;
  reg [7:0] sc2mac_dat_a_data119;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:350" *)
  output [7:0] sc2mac_dat_a_data12;
  reg [7:0] sc2mac_dat_a_data12;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:458" *)
  output [7:0] sc2mac_dat_a_data120;
  reg [7:0] sc2mac_dat_a_data120;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:459" *)
  output [7:0] sc2mac_dat_a_data121;
  reg [7:0] sc2mac_dat_a_data121;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:460" *)
  output [7:0] sc2mac_dat_a_data122;
  reg [7:0] sc2mac_dat_a_data122;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:461" *)
  output [7:0] sc2mac_dat_a_data123;
  reg [7:0] sc2mac_dat_a_data123;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:462" *)
  output [7:0] sc2mac_dat_a_data124;
  reg [7:0] sc2mac_dat_a_data124;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:463" *)
  output [7:0] sc2mac_dat_a_data125;
  reg [7:0] sc2mac_dat_a_data125;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:464" *)
  output [7:0] sc2mac_dat_a_data126;
  reg [7:0] sc2mac_dat_a_data126;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:465" *)
  output [7:0] sc2mac_dat_a_data127;
  reg [7:0] sc2mac_dat_a_data127;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:351" *)
  output [7:0] sc2mac_dat_a_data13;
  reg [7:0] sc2mac_dat_a_data13;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:352" *)
  output [7:0] sc2mac_dat_a_data14;
  reg [7:0] sc2mac_dat_a_data14;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:353" *)
  output [7:0] sc2mac_dat_a_data15;
  reg [7:0] sc2mac_dat_a_data15;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:354" *)
  output [7:0] sc2mac_dat_a_data16;
  reg [7:0] sc2mac_dat_a_data16;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:355" *)
  output [7:0] sc2mac_dat_a_data17;
  reg [7:0] sc2mac_dat_a_data17;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:356" *)
  output [7:0] sc2mac_dat_a_data18;
  reg [7:0] sc2mac_dat_a_data18;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:357" *)
  output [7:0] sc2mac_dat_a_data19;
  reg [7:0] sc2mac_dat_a_data19;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:340" *)
  output [7:0] sc2mac_dat_a_data2;
  reg [7:0] sc2mac_dat_a_data2;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:358" *)
  output [7:0] sc2mac_dat_a_data20;
  reg [7:0] sc2mac_dat_a_data20;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:359" *)
  output [7:0] sc2mac_dat_a_data21;
  reg [7:0] sc2mac_dat_a_data21;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:360" *)
  output [7:0] sc2mac_dat_a_data22;
  reg [7:0] sc2mac_dat_a_data22;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:361" *)
  output [7:0] sc2mac_dat_a_data23;
  reg [7:0] sc2mac_dat_a_data23;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:362" *)
  output [7:0] sc2mac_dat_a_data24;
  reg [7:0] sc2mac_dat_a_data24;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:363" *)
  output [7:0] sc2mac_dat_a_data25;
  reg [7:0] sc2mac_dat_a_data25;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:364" *)
  output [7:0] sc2mac_dat_a_data26;
  reg [7:0] sc2mac_dat_a_data26;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:365" *)
  output [7:0] sc2mac_dat_a_data27;
  reg [7:0] sc2mac_dat_a_data27;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:366" *)
  output [7:0] sc2mac_dat_a_data28;
  reg [7:0] sc2mac_dat_a_data28;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:367" *)
  output [7:0] sc2mac_dat_a_data29;
  reg [7:0] sc2mac_dat_a_data29;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:341" *)
  output [7:0] sc2mac_dat_a_data3;
  reg [7:0] sc2mac_dat_a_data3;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:368" *)
  output [7:0] sc2mac_dat_a_data30;
  reg [7:0] sc2mac_dat_a_data30;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:369" *)
  output [7:0] sc2mac_dat_a_data31;
  reg [7:0] sc2mac_dat_a_data31;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:370" *)
  output [7:0] sc2mac_dat_a_data32;
  reg [7:0] sc2mac_dat_a_data32;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:371" *)
  output [7:0] sc2mac_dat_a_data33;
  reg [7:0] sc2mac_dat_a_data33;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:372" *)
  output [7:0] sc2mac_dat_a_data34;
  reg [7:0] sc2mac_dat_a_data34;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:373" *)
  output [7:0] sc2mac_dat_a_data35;
  reg [7:0] sc2mac_dat_a_data35;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:374" *)
  output [7:0] sc2mac_dat_a_data36;
  reg [7:0] sc2mac_dat_a_data36;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:375" *)
  output [7:0] sc2mac_dat_a_data37;
  reg [7:0] sc2mac_dat_a_data37;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:376" *)
  output [7:0] sc2mac_dat_a_data38;
  reg [7:0] sc2mac_dat_a_data38;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:377" *)
  output [7:0] sc2mac_dat_a_data39;
  reg [7:0] sc2mac_dat_a_data39;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:342" *)
  output [7:0] sc2mac_dat_a_data4;
  reg [7:0] sc2mac_dat_a_data4;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:378" *)
  output [7:0] sc2mac_dat_a_data40;
  reg [7:0] sc2mac_dat_a_data40;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:379" *)
  output [7:0] sc2mac_dat_a_data41;
  reg [7:0] sc2mac_dat_a_data41;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:380" *)
  output [7:0] sc2mac_dat_a_data42;
  reg [7:0] sc2mac_dat_a_data42;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:381" *)
  output [7:0] sc2mac_dat_a_data43;
  reg [7:0] sc2mac_dat_a_data43;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:382" *)
  output [7:0] sc2mac_dat_a_data44;
  reg [7:0] sc2mac_dat_a_data44;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:383" *)
  output [7:0] sc2mac_dat_a_data45;
  reg [7:0] sc2mac_dat_a_data45;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:384" *)
  output [7:0] sc2mac_dat_a_data46;
  reg [7:0] sc2mac_dat_a_data46;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:385" *)
  output [7:0] sc2mac_dat_a_data47;
  reg [7:0] sc2mac_dat_a_data47;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:386" *)
  output [7:0] sc2mac_dat_a_data48;
  reg [7:0] sc2mac_dat_a_data48;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:387" *)
  output [7:0] sc2mac_dat_a_data49;
  reg [7:0] sc2mac_dat_a_data49;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:343" *)
  output [7:0] sc2mac_dat_a_data5;
  reg [7:0] sc2mac_dat_a_data5;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:388" *)
  output [7:0] sc2mac_dat_a_data50;
  reg [7:0] sc2mac_dat_a_data50;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:389" *)
  output [7:0] sc2mac_dat_a_data51;
  reg [7:0] sc2mac_dat_a_data51;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:390" *)
  output [7:0] sc2mac_dat_a_data52;
  reg [7:0] sc2mac_dat_a_data52;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:391" *)
  output [7:0] sc2mac_dat_a_data53;
  reg [7:0] sc2mac_dat_a_data53;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:392" *)
  output [7:0] sc2mac_dat_a_data54;
  reg [7:0] sc2mac_dat_a_data54;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:393" *)
  output [7:0] sc2mac_dat_a_data55;
  reg [7:0] sc2mac_dat_a_data55;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:394" *)
  output [7:0] sc2mac_dat_a_data56;
  reg [7:0] sc2mac_dat_a_data56;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:395" *)
  output [7:0] sc2mac_dat_a_data57;
  reg [7:0] sc2mac_dat_a_data57;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:396" *)
  output [7:0] sc2mac_dat_a_data58;
  reg [7:0] sc2mac_dat_a_data58;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:397" *)
  output [7:0] sc2mac_dat_a_data59;
  reg [7:0] sc2mac_dat_a_data59;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:344" *)
  output [7:0] sc2mac_dat_a_data6;
  reg [7:0] sc2mac_dat_a_data6;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:398" *)
  output [7:0] sc2mac_dat_a_data60;
  reg [7:0] sc2mac_dat_a_data60;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:399" *)
  output [7:0] sc2mac_dat_a_data61;
  reg [7:0] sc2mac_dat_a_data61;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:400" *)
  output [7:0] sc2mac_dat_a_data62;
  reg [7:0] sc2mac_dat_a_data62;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:401" *)
  output [7:0] sc2mac_dat_a_data63;
  reg [7:0] sc2mac_dat_a_data63;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:402" *)
  output [7:0] sc2mac_dat_a_data64;
  reg [7:0] sc2mac_dat_a_data64;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:403" *)
  output [7:0] sc2mac_dat_a_data65;
  reg [7:0] sc2mac_dat_a_data65;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:404" *)
  output [7:0] sc2mac_dat_a_data66;
  reg [7:0] sc2mac_dat_a_data66;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:405" *)
  output [7:0] sc2mac_dat_a_data67;
  reg [7:0] sc2mac_dat_a_data67;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:406" *)
  output [7:0] sc2mac_dat_a_data68;
  reg [7:0] sc2mac_dat_a_data68;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:407" *)
  output [7:0] sc2mac_dat_a_data69;
  reg [7:0] sc2mac_dat_a_data69;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:345" *)
  output [7:0] sc2mac_dat_a_data7;
  reg [7:0] sc2mac_dat_a_data7;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:408" *)
  output [7:0] sc2mac_dat_a_data70;
  reg [7:0] sc2mac_dat_a_data70;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:409" *)
  output [7:0] sc2mac_dat_a_data71;
  reg [7:0] sc2mac_dat_a_data71;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:410" *)
  output [7:0] sc2mac_dat_a_data72;
  reg [7:0] sc2mac_dat_a_data72;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:411" *)
  output [7:0] sc2mac_dat_a_data73;
  reg [7:0] sc2mac_dat_a_data73;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:412" *)
  output [7:0] sc2mac_dat_a_data74;
  reg [7:0] sc2mac_dat_a_data74;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:413" *)
  output [7:0] sc2mac_dat_a_data75;
  reg [7:0] sc2mac_dat_a_data75;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:414" *)
  output [7:0] sc2mac_dat_a_data76;
  reg [7:0] sc2mac_dat_a_data76;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:415" *)
  output [7:0] sc2mac_dat_a_data77;
  reg [7:0] sc2mac_dat_a_data77;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:416" *)
  output [7:0] sc2mac_dat_a_data78;
  reg [7:0] sc2mac_dat_a_data78;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:417" *)
  output [7:0] sc2mac_dat_a_data79;
  reg [7:0] sc2mac_dat_a_data79;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:346" *)
  output [7:0] sc2mac_dat_a_data8;
  reg [7:0] sc2mac_dat_a_data8;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:418" *)
  output [7:0] sc2mac_dat_a_data80;
  reg [7:0] sc2mac_dat_a_data80;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:419" *)
  output [7:0] sc2mac_dat_a_data81;
  reg [7:0] sc2mac_dat_a_data81;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:420" *)
  output [7:0] sc2mac_dat_a_data82;
  reg [7:0] sc2mac_dat_a_data82;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:421" *)
  output [7:0] sc2mac_dat_a_data83;
  reg [7:0] sc2mac_dat_a_data83;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:422" *)
  output [7:0] sc2mac_dat_a_data84;
  reg [7:0] sc2mac_dat_a_data84;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:423" *)
  output [7:0] sc2mac_dat_a_data85;
  reg [7:0] sc2mac_dat_a_data85;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:424" *)
  output [7:0] sc2mac_dat_a_data86;
  reg [7:0] sc2mac_dat_a_data86;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:425" *)
  output [7:0] sc2mac_dat_a_data87;
  reg [7:0] sc2mac_dat_a_data87;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:426" *)
  output [7:0] sc2mac_dat_a_data88;
  reg [7:0] sc2mac_dat_a_data88;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:427" *)
  output [7:0] sc2mac_dat_a_data89;
  reg [7:0] sc2mac_dat_a_data89;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:347" *)
  output [7:0] sc2mac_dat_a_data9;
  reg [7:0] sc2mac_dat_a_data9;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:428" *)
  output [7:0] sc2mac_dat_a_data90;
  reg [7:0] sc2mac_dat_a_data90;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:429" *)
  output [7:0] sc2mac_dat_a_data91;
  reg [7:0] sc2mac_dat_a_data91;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:430" *)
  output [7:0] sc2mac_dat_a_data92;
  reg [7:0] sc2mac_dat_a_data92;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:431" *)
  output [7:0] sc2mac_dat_a_data93;
  reg [7:0] sc2mac_dat_a_data93;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:432" *)
  output [7:0] sc2mac_dat_a_data94;
  reg [7:0] sc2mac_dat_a_data94;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:433" *)
  output [7:0] sc2mac_dat_a_data95;
  reg [7:0] sc2mac_dat_a_data95;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:434" *)
  output [7:0] sc2mac_dat_a_data96;
  reg [7:0] sc2mac_dat_a_data96;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:435" *)
  output [7:0] sc2mac_dat_a_data97;
  reg [7:0] sc2mac_dat_a_data97;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:436" *)
  output [7:0] sc2mac_dat_a_data98;
  reg [7:0] sc2mac_dat_a_data98;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:437" *)
  output [7:0] sc2mac_dat_a_data99;
  reg [7:0] sc2mac_dat_a_data99;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:337" *)
  output [127:0] sc2mac_dat_a_mask;
  reg [127:0] sc2mac_dat_a_mask;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:466" *)
  output [8:0] sc2mac_dat_a_pd;
  reg [8:0] sc2mac_dat_a_pd;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:336" *)
  output sc2mac_dat_a_pvld;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:469" *)
  output [7:0] sc2mac_dat_b_data0;
  reg [7:0] sc2mac_dat_b_data0;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:470" *)
  output [7:0] sc2mac_dat_b_data1;
  reg [7:0] sc2mac_dat_b_data1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:479" *)
  output [7:0] sc2mac_dat_b_data10;
  reg [7:0] sc2mac_dat_b_data10;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:569" *)
  output [7:0] sc2mac_dat_b_data100;
  reg [7:0] sc2mac_dat_b_data100;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:570" *)
  output [7:0] sc2mac_dat_b_data101;
  reg [7:0] sc2mac_dat_b_data101;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:571" *)
  output [7:0] sc2mac_dat_b_data102;
  reg [7:0] sc2mac_dat_b_data102;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:572" *)
  output [7:0] sc2mac_dat_b_data103;
  reg [7:0] sc2mac_dat_b_data103;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:573" *)
  output [7:0] sc2mac_dat_b_data104;
  reg [7:0] sc2mac_dat_b_data104;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:574" *)
  output [7:0] sc2mac_dat_b_data105;
  reg [7:0] sc2mac_dat_b_data105;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:575" *)
  output [7:0] sc2mac_dat_b_data106;
  reg [7:0] sc2mac_dat_b_data106;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:576" *)
  output [7:0] sc2mac_dat_b_data107;
  reg [7:0] sc2mac_dat_b_data107;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:577" *)
  output [7:0] sc2mac_dat_b_data108;
  reg [7:0] sc2mac_dat_b_data108;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:578" *)
  output [7:0] sc2mac_dat_b_data109;
  reg [7:0] sc2mac_dat_b_data109;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:480" *)
  output [7:0] sc2mac_dat_b_data11;
  reg [7:0] sc2mac_dat_b_data11;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:579" *)
  output [7:0] sc2mac_dat_b_data110;
  reg [7:0] sc2mac_dat_b_data110;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:580" *)
  output [7:0] sc2mac_dat_b_data111;
  reg [7:0] sc2mac_dat_b_data111;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:581" *)
  output [7:0] sc2mac_dat_b_data112;
  reg [7:0] sc2mac_dat_b_data112;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:582" *)
  output [7:0] sc2mac_dat_b_data113;
  reg [7:0] sc2mac_dat_b_data113;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:583" *)
  output [7:0] sc2mac_dat_b_data114;
  reg [7:0] sc2mac_dat_b_data114;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:584" *)
  output [7:0] sc2mac_dat_b_data115;
  reg [7:0] sc2mac_dat_b_data115;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:585" *)
  output [7:0] sc2mac_dat_b_data116;
  reg [7:0] sc2mac_dat_b_data116;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:586" *)
  output [7:0] sc2mac_dat_b_data117;
  reg [7:0] sc2mac_dat_b_data117;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:587" *)
  output [7:0] sc2mac_dat_b_data118;
  reg [7:0] sc2mac_dat_b_data118;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:588" *)
  output [7:0] sc2mac_dat_b_data119;
  reg [7:0] sc2mac_dat_b_data119;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:481" *)
  output [7:0] sc2mac_dat_b_data12;
  reg [7:0] sc2mac_dat_b_data12;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:589" *)
  output [7:0] sc2mac_dat_b_data120;
  reg [7:0] sc2mac_dat_b_data120;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:590" *)
  output [7:0] sc2mac_dat_b_data121;
  reg [7:0] sc2mac_dat_b_data121;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:591" *)
  output [7:0] sc2mac_dat_b_data122;
  reg [7:0] sc2mac_dat_b_data122;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:592" *)
  output [7:0] sc2mac_dat_b_data123;
  reg [7:0] sc2mac_dat_b_data123;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:593" *)
  output [7:0] sc2mac_dat_b_data124;
  reg [7:0] sc2mac_dat_b_data124;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:594" *)
  output [7:0] sc2mac_dat_b_data125;
  reg [7:0] sc2mac_dat_b_data125;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:595" *)
  output [7:0] sc2mac_dat_b_data126;
  reg [7:0] sc2mac_dat_b_data126;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:596" *)
  output [7:0] sc2mac_dat_b_data127;
  reg [7:0] sc2mac_dat_b_data127;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:482" *)
  output [7:0] sc2mac_dat_b_data13;
  reg [7:0] sc2mac_dat_b_data13;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:483" *)
  output [7:0] sc2mac_dat_b_data14;
  reg [7:0] sc2mac_dat_b_data14;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:484" *)
  output [7:0] sc2mac_dat_b_data15;
  reg [7:0] sc2mac_dat_b_data15;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:485" *)
  output [7:0] sc2mac_dat_b_data16;
  reg [7:0] sc2mac_dat_b_data16;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:486" *)
  output [7:0] sc2mac_dat_b_data17;
  reg [7:0] sc2mac_dat_b_data17;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:487" *)
  output [7:0] sc2mac_dat_b_data18;
  reg [7:0] sc2mac_dat_b_data18;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:488" *)
  output [7:0] sc2mac_dat_b_data19;
  reg [7:0] sc2mac_dat_b_data19;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:471" *)
  output [7:0] sc2mac_dat_b_data2;
  reg [7:0] sc2mac_dat_b_data2;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:489" *)
  output [7:0] sc2mac_dat_b_data20;
  reg [7:0] sc2mac_dat_b_data20;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:490" *)
  output [7:0] sc2mac_dat_b_data21;
  reg [7:0] sc2mac_dat_b_data21;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:491" *)
  output [7:0] sc2mac_dat_b_data22;
  reg [7:0] sc2mac_dat_b_data22;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:492" *)
  output [7:0] sc2mac_dat_b_data23;
  reg [7:0] sc2mac_dat_b_data23;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:493" *)
  output [7:0] sc2mac_dat_b_data24;
  reg [7:0] sc2mac_dat_b_data24;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:494" *)
  output [7:0] sc2mac_dat_b_data25;
  reg [7:0] sc2mac_dat_b_data25;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:495" *)
  output [7:0] sc2mac_dat_b_data26;
  reg [7:0] sc2mac_dat_b_data26;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:496" *)
  output [7:0] sc2mac_dat_b_data27;
  reg [7:0] sc2mac_dat_b_data27;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:497" *)
  output [7:0] sc2mac_dat_b_data28;
  reg [7:0] sc2mac_dat_b_data28;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:498" *)
  output [7:0] sc2mac_dat_b_data29;
  reg [7:0] sc2mac_dat_b_data29;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:472" *)
  output [7:0] sc2mac_dat_b_data3;
  reg [7:0] sc2mac_dat_b_data3;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:499" *)
  output [7:0] sc2mac_dat_b_data30;
  reg [7:0] sc2mac_dat_b_data30;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:500" *)
  output [7:0] sc2mac_dat_b_data31;
  reg [7:0] sc2mac_dat_b_data31;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:501" *)
  output [7:0] sc2mac_dat_b_data32;
  reg [7:0] sc2mac_dat_b_data32;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:502" *)
  output [7:0] sc2mac_dat_b_data33;
  reg [7:0] sc2mac_dat_b_data33;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:503" *)
  output [7:0] sc2mac_dat_b_data34;
  reg [7:0] sc2mac_dat_b_data34;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:504" *)
  output [7:0] sc2mac_dat_b_data35;
  reg [7:0] sc2mac_dat_b_data35;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:505" *)
  output [7:0] sc2mac_dat_b_data36;
  reg [7:0] sc2mac_dat_b_data36;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:506" *)
  output [7:0] sc2mac_dat_b_data37;
  reg [7:0] sc2mac_dat_b_data37;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:507" *)
  output [7:0] sc2mac_dat_b_data38;
  reg [7:0] sc2mac_dat_b_data38;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:508" *)
  output [7:0] sc2mac_dat_b_data39;
  reg [7:0] sc2mac_dat_b_data39;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:473" *)
  output [7:0] sc2mac_dat_b_data4;
  reg [7:0] sc2mac_dat_b_data4;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:509" *)
  output [7:0] sc2mac_dat_b_data40;
  reg [7:0] sc2mac_dat_b_data40;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:510" *)
  output [7:0] sc2mac_dat_b_data41;
  reg [7:0] sc2mac_dat_b_data41;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:511" *)
  output [7:0] sc2mac_dat_b_data42;
  reg [7:0] sc2mac_dat_b_data42;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:512" *)
  output [7:0] sc2mac_dat_b_data43;
  reg [7:0] sc2mac_dat_b_data43;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:513" *)
  output [7:0] sc2mac_dat_b_data44;
  reg [7:0] sc2mac_dat_b_data44;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:514" *)
  output [7:0] sc2mac_dat_b_data45;
  reg [7:0] sc2mac_dat_b_data45;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:515" *)
  output [7:0] sc2mac_dat_b_data46;
  reg [7:0] sc2mac_dat_b_data46;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:516" *)
  output [7:0] sc2mac_dat_b_data47;
  reg [7:0] sc2mac_dat_b_data47;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:517" *)
  output [7:0] sc2mac_dat_b_data48;
  reg [7:0] sc2mac_dat_b_data48;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:518" *)
  output [7:0] sc2mac_dat_b_data49;
  reg [7:0] sc2mac_dat_b_data49;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:474" *)
  output [7:0] sc2mac_dat_b_data5;
  reg [7:0] sc2mac_dat_b_data5;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:519" *)
  output [7:0] sc2mac_dat_b_data50;
  reg [7:0] sc2mac_dat_b_data50;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:520" *)
  output [7:0] sc2mac_dat_b_data51;
  reg [7:0] sc2mac_dat_b_data51;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:521" *)
  output [7:0] sc2mac_dat_b_data52;
  reg [7:0] sc2mac_dat_b_data52;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:522" *)
  output [7:0] sc2mac_dat_b_data53;
  reg [7:0] sc2mac_dat_b_data53;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:523" *)
  output [7:0] sc2mac_dat_b_data54;
  reg [7:0] sc2mac_dat_b_data54;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:524" *)
  output [7:0] sc2mac_dat_b_data55;
  reg [7:0] sc2mac_dat_b_data55;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:525" *)
  output [7:0] sc2mac_dat_b_data56;
  reg [7:0] sc2mac_dat_b_data56;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:526" *)
  output [7:0] sc2mac_dat_b_data57;
  reg [7:0] sc2mac_dat_b_data57;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:527" *)
  output [7:0] sc2mac_dat_b_data58;
  reg [7:0] sc2mac_dat_b_data58;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:528" *)
  output [7:0] sc2mac_dat_b_data59;
  reg [7:0] sc2mac_dat_b_data59;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:475" *)
  output [7:0] sc2mac_dat_b_data6;
  reg [7:0] sc2mac_dat_b_data6;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:529" *)
  output [7:0] sc2mac_dat_b_data60;
  reg [7:0] sc2mac_dat_b_data60;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:530" *)
  output [7:0] sc2mac_dat_b_data61;
  reg [7:0] sc2mac_dat_b_data61;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:531" *)
  output [7:0] sc2mac_dat_b_data62;
  reg [7:0] sc2mac_dat_b_data62;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:532" *)
  output [7:0] sc2mac_dat_b_data63;
  reg [7:0] sc2mac_dat_b_data63;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:533" *)
  output [7:0] sc2mac_dat_b_data64;
  reg [7:0] sc2mac_dat_b_data64;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:534" *)
  output [7:0] sc2mac_dat_b_data65;
  reg [7:0] sc2mac_dat_b_data65;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:535" *)
  output [7:0] sc2mac_dat_b_data66;
  reg [7:0] sc2mac_dat_b_data66;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:536" *)
  output [7:0] sc2mac_dat_b_data67;
  reg [7:0] sc2mac_dat_b_data67;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:537" *)
  output [7:0] sc2mac_dat_b_data68;
  reg [7:0] sc2mac_dat_b_data68;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:538" *)
  output [7:0] sc2mac_dat_b_data69;
  reg [7:0] sc2mac_dat_b_data69;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:476" *)
  output [7:0] sc2mac_dat_b_data7;
  reg [7:0] sc2mac_dat_b_data7;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:539" *)
  output [7:0] sc2mac_dat_b_data70;
  reg [7:0] sc2mac_dat_b_data70;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:540" *)
  output [7:0] sc2mac_dat_b_data71;
  reg [7:0] sc2mac_dat_b_data71;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:541" *)
  output [7:0] sc2mac_dat_b_data72;
  reg [7:0] sc2mac_dat_b_data72;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:542" *)
  output [7:0] sc2mac_dat_b_data73;
  reg [7:0] sc2mac_dat_b_data73;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:543" *)
  output [7:0] sc2mac_dat_b_data74;
  reg [7:0] sc2mac_dat_b_data74;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:544" *)
  output [7:0] sc2mac_dat_b_data75;
  reg [7:0] sc2mac_dat_b_data75;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:545" *)
  output [7:0] sc2mac_dat_b_data76;
  reg [7:0] sc2mac_dat_b_data76;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:546" *)
  output [7:0] sc2mac_dat_b_data77;
  reg [7:0] sc2mac_dat_b_data77;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:547" *)
  output [7:0] sc2mac_dat_b_data78;
  reg [7:0] sc2mac_dat_b_data78;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:548" *)
  output [7:0] sc2mac_dat_b_data79;
  reg [7:0] sc2mac_dat_b_data79;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:477" *)
  output [7:0] sc2mac_dat_b_data8;
  reg [7:0] sc2mac_dat_b_data8;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:549" *)
  output [7:0] sc2mac_dat_b_data80;
  reg [7:0] sc2mac_dat_b_data80;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:550" *)
  output [7:0] sc2mac_dat_b_data81;
  reg [7:0] sc2mac_dat_b_data81;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:551" *)
  output [7:0] sc2mac_dat_b_data82;
  reg [7:0] sc2mac_dat_b_data82;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:552" *)
  output [7:0] sc2mac_dat_b_data83;
  reg [7:0] sc2mac_dat_b_data83;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:553" *)
  output [7:0] sc2mac_dat_b_data84;
  reg [7:0] sc2mac_dat_b_data84;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:554" *)
  output [7:0] sc2mac_dat_b_data85;
  reg [7:0] sc2mac_dat_b_data85;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:555" *)
  output [7:0] sc2mac_dat_b_data86;
  reg [7:0] sc2mac_dat_b_data86;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:556" *)
  output [7:0] sc2mac_dat_b_data87;
  reg [7:0] sc2mac_dat_b_data87;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:557" *)
  output [7:0] sc2mac_dat_b_data88;
  reg [7:0] sc2mac_dat_b_data88;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:558" *)
  output [7:0] sc2mac_dat_b_data89;
  reg [7:0] sc2mac_dat_b_data89;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:478" *)
  output [7:0] sc2mac_dat_b_data9;
  reg [7:0] sc2mac_dat_b_data9;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:559" *)
  output [7:0] sc2mac_dat_b_data90;
  reg [7:0] sc2mac_dat_b_data90;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:560" *)
  output [7:0] sc2mac_dat_b_data91;
  reg [7:0] sc2mac_dat_b_data91;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:561" *)
  output [7:0] sc2mac_dat_b_data92;
  reg [7:0] sc2mac_dat_b_data92;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:562" *)
  output [7:0] sc2mac_dat_b_data93;
  reg [7:0] sc2mac_dat_b_data93;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:563" *)
  output [7:0] sc2mac_dat_b_data94;
  reg [7:0] sc2mac_dat_b_data94;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:564" *)
  output [7:0] sc2mac_dat_b_data95;
  reg [7:0] sc2mac_dat_b_data95;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:565" *)
  output [7:0] sc2mac_dat_b_data96;
  reg [7:0] sc2mac_dat_b_data96;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:566" *)
  output [7:0] sc2mac_dat_b_data97;
  reg [7:0] sc2mac_dat_b_data97;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:567" *)
  output [7:0] sc2mac_dat_b_data98;
  reg [7:0] sc2mac_dat_b_data98;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:568" *)
  output [7:0] sc2mac_dat_b_data99;
  reg [7:0] sc2mac_dat_b_data99;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:468" *)
  output [127:0] sc2mac_dat_b_mask;
  reg [127:0] sc2mac_dat_b_mask;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:597" *)
  output [8:0] sc2mac_dat_b_pd;
  reg [8:0] sc2mac_dat_b_pd;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:467" *)
  output sc2mac_dat_b_pvld;
  reg sc2mac_dat_b_pvld;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1807" *)
  wire [8:0] sc2mac_dat_pd_w;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:323" *)
  input [1:0] sc_state;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:322" *)
  input [30:0] sg2dl_pd;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:321" *)
  input sg2dl_pvld;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:324" *)
  input sg2dl_reuse_rls;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:623" *)
  output slcg_wg_en;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1808" *)
  reg slcg_wg_en_d1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1809" *)
  reg slcg_wg_en_d2;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1810" *)
  reg slcg_wg_en_d3;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:903" *)
  wire slcg_wg_en_w;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1811" *)
  wire [11:0] slice_entries_w;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1812" *)
  reg [11:0] slice_left;
  wire [11:0] slice_left_w;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1814" *)
  wire [11:0] slices_oprand;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1815" *)
  reg [6:0] stripe_cnt;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1816" *)
  wire [6:0] stripe_cnt_inc;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1817" *)
  wire stripe_cnt_reg_en;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1818" *)
  wire [6:0] stripe_cnt_w;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1819" *)
  reg [2:0] sub_h_cmp_g0;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1820" *)
  reg [2:0] sub_h_cmp_g1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1821" *)
  wire [2:0] sub_h_cmp_w;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1822" *)
  reg [1:0] sub_h_cnt;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1823" *)
  wire [2:0] sub_h_cnt_inc;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1824" *)
  wire sub_h_cnt_reg_en;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1825" *)
  wire [1:0] sub_h_cnt_w;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1826" *)
  reg [2:0] sub_h_total_g0;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1827" *)
  reg [2:0] sub_h_total_g1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1828" *)
  reg [2:0] sub_h_total_g10;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1829" *)
  reg [2:0] sub_h_total_g11;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1830" *)
  reg [1:0] sub_h_total_g2;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1831" *)
  reg [2:0] sub_h_total_g3;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1832" *)
  reg [2:0] sub_h_total_g4;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1833" *)
  reg [2:0] sub_h_total_g5;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1834" *)
  reg [2:0] sub_h_total_g6;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1835" *)
  reg [2:0] sub_h_total_g7;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1836" *)
  reg [2:0] sub_h_total_g8;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1837" *)
  reg [2:0] sub_h_total_g9;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1838" *)
  wire [2:0] sub_h_total_w;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1839" *)
  wire sub_rls;
  wire [13:0] w_bias_16;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1841" *)
  reg [11:0] w_bias_d1;
  wire [13:0] w_bias_int8;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:904" *)
  wire w_bias_reg_en;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1843" *)
  (* unused_bits = "0 1" *)
  wire [13:0] w_bias_w;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1844" *)
  reg [5:0] x_dilate;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1845" *)
  wire [5:0] x_dilate_w;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1846" *)
  reg [5:0] y_dilate;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1847" *)
  wire [5:0] y_dilate_w;
  assign datain_h_cnt_inc = datain_h_cnt + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:10231" *) conv_y_stride;
  assign _0703_ = datain_h_cnt + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:10278" *) dl_h_offset_ext;
  assign datain_h_cur = _0703_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:10278" *) sub_h_cnt;
  assign _0704_ = c_bias + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:11343" *) c_bias_add;
  assign _0705_ = h_bias_0_d1 + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:12149" *) h_bias_1_d1;
  assign _0706_ = _0705_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:12149" *) h_bias_2_d1;
  assign h_bias_d1 = _0706_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:12149" *) h_bias_3_d1;
  assign _0707_ = dat_entry_st + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:12157" *) c_bias_d1;
  assign _0708_ = _0707_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:12157" *) h_bias_d1;
  assign dat_req_addr_sum = _0708_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:12157" *) w_bias_d1;
  assign _0709_ = rsp_sft_cnt_l0 + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15136" *) pixel_x_byte_stride;
  assign _0710_ = rsp_sft_cnt_l1 + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15144" *) pixel_x_byte_stride;
  assign _0711_ = rsp_sft_cnt_l2 + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15152" *) pixel_x_byte_stride;
  assign _0712_ = rsp_sft_cnt_l3 + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15160" *) pixel_x_byte_stride;
  assign data_bank_w = reg2dp_data_bank + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1933" *) 1'b1;
  assign _0713_ = reg2dp_batches + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1941" *) 1'b1;
  assign _0714_ = reg2dp_datain_width_ext[12:2] + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1964" *) 1'b1;
  assign _0715_ = reg2dp_datain_width_ext + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1965" *) 1'b1;
  assign _0716_ = reg2dp_conv_x_stride_ext + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:2011" *) 1'b1;
  assign _0717_ = { conv_x_stride_w, 1'b0 } + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:2018" *) conv_x_stride_w;
  assign _0718_ = { pixel_x_stride_w[4:0], 1'b0 } + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:2027" *) pixel_x_stride_w;
  assign _0719_ = _0718_ + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:2027" *) reg2dp_weight_channel_ext[5:0];
  assign _0720_ = pixel_x_stride_w + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:2028" *) reg2dp_weight_channel_ext[5:0];
  assign pixel_x_init_offset_w = reg2dp_weight_channel_ext[5:0] + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:2035" *) 1'b1;
  assign _0721_ = reg2dp_conv_y_stride_ext + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:2061" *) 1'b1;
  assign _0722_ = reg2dp_x_dilation_ext + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:2069" *) 1'b1;
  assign _0723_ = reg2dp_y_dilation_ext + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:2077" *) 1'b1;
  assign entries_single_w = reg2dp_entries + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:2083" *) 1'b1;
  assign _0724_ = { reg2dp_entries[9:0], 2'b00 } + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:2098" *) 3'b100;
  assign rls_slices_w = reg2dp_rls_slices + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:2125" *) 1'b1;
  assign _0725_ = reg2dp_datain_height_ext[11:0] + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:2133" *) 1'b1;
  assign dat_entry_st_inc = dat_entry_st + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:6702" *) dat_entry_avl_sub;
  assign _0726_[4:0] = batch_cnt + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:8539" *) 1'b1;
  assign sub_h_cnt_inc = sub_h_cnt + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:8706" *) 1'b1;
  assign stripe_cnt_inc = stripe_cnt + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:8796" *) 1'b1;
  assign dataout_w_cnt_inc = dataout_w_cnt + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:9340" *) sub_h_cmp_g1;
  assign datain_c_cnt_inc = datain_c_cnt + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:9514" *) 1'b1;
  assign _0727_[13:0] = datain_w_cnt + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:9616" *) 2'b10;
  assign _0728_[13:0] = datain_w_cnt + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:9617" *) conv_x_stride;
  assign _0729_[15:0] = pixel_w_ch_ori + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:9656" *) pixel_ch_stride;
  assign _0730_[15:0] = pixel_w_ch_ori + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:9657" *) pixel_x_init_offset;
  assign _0731_[15:0] = pixel_w_cnt + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:9659" *) pixel_x_cnt_add;
  assign datain_w_cur = datain_w_cnt + (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:9719" *) dl_w_offset_ext;
  assign _0732_ = is_stripe_end & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:10244" *) dl_pd[28];
  assign _0733_ = is_stripe_end & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:10245" *) _1078_;
  assign _0734_ = dat_exec_valid & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:10256" *) _1124_;
  assign _0735_ = dat_exec_valid & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:10264" *) is_stripe_end;
  assign _0736_ = _0735_ & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:10264" *) dl_pd[27];
  assign _0737_ = _1157_ & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:10417" *) datain_w_cur[1];
  assign dat_wg_req_skip = _0737_ & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:10417" *) _1158_;
  assign _0738_ = is_winograd_d1[5] & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:10448" *) dat_wg_req_skip;
  assign _0739_ = is_img_d1[6] & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:10448" *) dat_img_req_skip;
  assign _0740_ = dat_exec_valid & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:10455" *) _1079_;
  assign dat_req_valid = _0740_ & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:10455" *) _1080_;
  assign _0741_ = is_int8_d1[2] & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:10464" *) datain_c_cnt[0];
  assign dat_req_sub_w_st_en = dat_exec_valid & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:10474" *) _1026_;
  assign dat_req_stripe_end = is_stripe_equal & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:10477" *) dat_pipe_valid;
  assign _0742_ = dl_pd[30] & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:11047" *) is_stripe_equal;
  assign _0743_ = _0742_ & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:11047" *) dat_pipe_valid;
  assign _0744_ = _1082_ & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:11330" *) _1127_;
  assign _0745_ = is_stripe_end & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:11342" *) dl_pd[27];
  assign _0746_ = _0735_ & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:11351" *) dl_pd[26];
  assign _0747_ = dat_exec_valid & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:11391" *) _1128_;
  assign sc2buf_dat_rd_en_w = dat_req_valid_d1 & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:12188" *) _1133_;
  assign _0748_ = _1134_ & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:12194" *) _1027_;
  assign _0749_ = _1134_ & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:12195" *) _1028_;
  assign _0750_ = _1134_ & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:12196" *) _1029_;
  assign _0751_ = _1134_ & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:12197" *) _1030_;
  assign dat_l0c0_en = sc2buf_dat_rd_valid & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:14531" *) _1032_;
  assign dat_l1c0_en = sc2buf_dat_rd_valid & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:14532" *) _1033_;
  assign dat_l1c0_hi_en = dat_l1c0_en & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:14533" *) _1085_;
  assign dat_l2c0_en = sc2buf_dat_rd_valid & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:14535" *) _1034_;
  assign dat_l3c0_en = sc2buf_dat_rd_valid & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:14537" *) _1035_;
  assign _0752_ = dat_wg_adv & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:14552" *) _1086_;
  assign _0753_ = is_img_d1[12] & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:14553" *) dat_l0c0_en;
  assign _0754_ = _0753_ & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:14553" *) _1087_;
  assign _0755_ = dat_wg_adv & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:14554" *) dat_rsp_exec_sub_h_d6[0];
  assign _0756_ = is_img_d1[13] & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:14555" *) dat_l1c0_en;
  assign _0757_ = _0756_ & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:14555" *) _1088_;
  assign _0758_ = is_img_d1[14] & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:14556" *) dat_l1c0_en;
  assign dat_l1c1_hi_en = _0758_ & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:14556" *) _1088_;
  assign _0759_ = is_img_d1[15] & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:14557" *) dat_l2c0_en;
  assign dat_l2c1_en = _0759_ & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:14557" *) _1089_;
  assign _0760_ = is_img_d1[16] & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:14558" *) dat_l3c0_en;
  assign dat_l3c1_en = _0760_ & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:14558" *) _1090_;
  assign _0761_ = dat_rsp_exec_pvld_d6 & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:14560" *) dat_rsp_exec_dummy_d6;
  assign dat_dummy_l0_en = _0761_ & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:14560" *) _1032_;
  assign dat_dummy_l1_en = _0761_ & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:14561" *) _1033_;
  assign dat_dummy_l2_en = _0761_ & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:14562" *) _1034_;
  assign dat_dummy_l3_en = _0761_ & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:14563" *) _1035_;
  assign _0762_ = sc2buf_dat_rd_valid & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:14564" *) is_winograd_d1[11];
  assign dat_wg_adv = _0762_ & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:14564" *) _1091_;
  assign _0763_ = dat_l1_set & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:14581" *) _1159_;
  assign _0764_ = dat_l2_set & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:14584" *) sub_h_total_g2[1];
  assign _0765_ = dat_l3_set & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:14587" *) sub_h_total_g2[1];
  assign _0766_ = sub_h_total_g3[2] & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15041" *) dat_rsp_pvld_d4;
  assign _0767_ = sub_h_total_g3[1] & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15042" *) dat_rsp_pvld_d2;
  assign _0768_ = sub_h_total_g3[0] & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15043" *) dat_rsp_pvld_d1;
  assign { _1017_[26:12], _0769_ } = { sub_h_total_g4[2], sub_h_total_g4[2], sub_h_total_g4[2], sub_h_total_g4[2], sub_h_total_g4[2], sub_h_total_g4[2], sub_h_total_g4[2], sub_h_total_g4[2], sub_h_total_g4[2], sub_h_total_g4[2], sub_h_total_g4[2], sub_h_total_g4[2], sub_h_total_g4[2], sub_h_total_g4[2], sub_h_total_g4[2], sub_h_total_g4[2], sub_h_total_g4[2], sub_h_total_g4[2], sub_h_total_g4[2], sub_h_total_g4[2], sub_h_total_g4[2], sub_h_total_g4[2], sub_h_total_g4[2], sub_h_total_g4[2], sub_h_total_g4[2], sub_h_total_g4[2], sub_h_total_g4[2] } & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15062" *) dat_rsp_pd_d4;
  assign _0770_ = { sub_h_total_g4[1], sub_h_total_g4[1], sub_h_total_g4[1], sub_h_total_g4[1], sub_h_total_g4[1], sub_h_total_g4[1], sub_h_total_g4[1], sub_h_total_g4[1], sub_h_total_g4[1], sub_h_total_g4[1], sub_h_total_g4[1], sub_h_total_g4[1], sub_h_total_g4[1], sub_h_total_g4[1], sub_h_total_g4[1], sub_h_total_g4[1], sub_h_total_g4[1], sub_h_total_g4[1], sub_h_total_g4[1], sub_h_total_g4[1], sub_h_total_g4[1], sub_h_total_g4[1], sub_h_total_g4[1], sub_h_total_g4[1], sub_h_total_g4[1], sub_h_total_g4[1], sub_h_total_g4[1] } & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15063" *) dat_rsp_pd_d2;
  assign _0771_ = { sub_h_total_g4[0], sub_h_total_g4[0], sub_h_total_g4[0], sub_h_total_g4[0], sub_h_total_g4[0], sub_h_total_g4[0], sub_h_total_g4[0], sub_h_total_g4[0], sub_h_total_g4[0], sub_h_total_g4[0], sub_h_total_g4[0], sub_h_total_g4[0], sub_h_total_g4[0], sub_h_total_g4[0], sub_h_total_g4[0], sub_h_total_g4[0], sub_h_total_g4[0], sub_h_total_g4[0], sub_h_total_g4[0], sub_h_total_g4[0], sub_h_total_g4[0], sub_h_total_g4[0], sub_h_total_g4[0], sub_h_total_g4[0], sub_h_total_g4[0], sub_h_total_g4[0], sub_h_total_g4[0] } & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15064" *) dat_rsp_pd_d1;
  assign _0772_ = dat_rsp_pd_d1[24] & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15176" *) _1092_;
  assign _0773_ = dat_rsp_pd_d1[24] & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15177" *) dat_rsp_pd_d1[4];
  assign _0774_ = _0773_ & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15177" *) dat_rsp_pd_d1[6];
  assign _0775_ = _0773_ & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15178" *) _1093_;
  assign _0776_ = rsp_sft_cnt_l0_inc & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15179" *) 7'b1111111;
  assign _0777_ = dat_rsp_pd_d2[24] & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15192" *) _1094_;
  assign _0778_ = dat_rsp_pd_d2[24] & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15193" *) dat_rsp_pd_d2[4];
  assign _0779_ = _0778_ & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15193" *) dat_rsp_pd_d2[6];
  assign _0780_ = _0778_ & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15194" *) _1095_;
  assign _0781_ = rsp_sft_cnt_l1_inc & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15195" *) 7'b1111111;
  assign _0782_ = dat_rsp_pd_d3[24] & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15208" *) _1096_;
  assign _0783_ = dat_rsp_pd_d3[24] & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15209" *) dat_rsp_pd_d3[4];
  assign _0784_ = _0783_ & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15209" *) dat_rsp_pd_d3[6];
  assign _0785_ = _0783_ & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15210" *) _1097_;
  assign _0786_ = rsp_sft_cnt_l2_inc & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15211" *) 7'b1111111;
  assign _0787_ = dat_rsp_pd_d4[24] & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15224" *) _1098_;
  assign _0788_ = dat_rsp_pd_d4[24] & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15225" *) dat_rsp_pd_d4[4];
  assign _0789_ = _0788_ & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15225" *) dat_rsp_pd_d4[6];
  assign _0790_ = _0788_ & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15226" *) _1099_;
  assign _0791_ = rsp_sft_cnt_l3_inc & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15227" *) 7'b1111111;
  assign _0792_ = is_img_d1[17] & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15239" *) dat_rsp_pvld_d1;
  assign _0793_ = is_img_d1[18] & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15240" *) dat_rsp_pvld_d2;
  assign _0794_ = _0793_ & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15240" *) _1075_;
  assign _0795_ = is_img_d1[19] & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15241" *) dat_rsp_pvld_d3;
  assign _0796_ = _0795_ & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15241" *) _1036_;
  assign _0797_ = is_img_d1[20] & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15242" *) dat_rsp_pvld_d4;
  assign _0798_ = _0797_ & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15242" *) _1036_;
  assign _0799_ = is_img_d1[21] & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15261" *) dat_rsp_pvld_d1;
  assign _0800_ = _0799_ & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15261" *) dat_rsp_pd_d1[24];
  assign _0801_ = _0800_ & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15261" *) dat_rsp_pd_d1[4];
  assign _0802_ = is_img_d1[22] & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15262" *) dat_rsp_pvld_d2;
  assign _0803_ = _0802_ & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15262" *) dat_rsp_pd_d2[24];
  assign _0804_ = _0803_ & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15262" *) dat_rsp_pd_d2[4];
  assign _0805_ = _0804_ & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15262" *) _1076_;
  assign _0806_ = is_img_d1[23] & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15263" *) dat_rsp_pvld_d3;
  assign _0807_ = _0806_ & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15263" *) dat_rsp_pd_d3[24];
  assign _0808_ = _0807_ & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15263" *) dat_rsp_pd_d3[4];
  assign _0809_ = _0808_ & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15263" *) _1037_;
  assign _0810_ = is_img_d1[24] & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15264" *) dat_rsp_pvld_d4;
  assign _0811_ = _0810_ & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15264" *) dat_rsp_pd_d4[24];
  assign _0812_ = _0811_ & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15264" *) dat_rsp_pd_d4[4];
  assign _0813_ = _0812_ & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15264" *) _1037_;
  assign dat_rsp_wg_sel_lt = _1100_ & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15780" *) _1038_;
  assign dat_rsp_wg_sel_lb = dat_rsp_pd[2] & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15781" *) _1038_;
  assign dat_rsp_wg_sel_rt = _1100_ & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15782" *) dat_rsp_pd[0];
  assign dat_rsp_wg_sel_rb = dat_rsp_pd[2] & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15783" *) dat_rsp_pd[0];
  assign dat_rsp_wg_sel_8b_lo = is_int8_d1[6] & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15790" *) _1101_;
  assign dat_rsp_wg_sel_8b_hi = is_int8_d1[7] & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15791" *) dat_rsp_pd[4];
  assign _0814_ = { dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt, dat_rsp_wg_sel_lt } & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15811" *) { dat_wg[1535:1280], dat_wg[1151:896], dat_wg[767:512], dat_wg[383:128] };
  assign _0815_ = { dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb, dat_rsp_wg_sel_lb } & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15812" *) { dat_wg[2303:2048], dat_wg[1919:1664], dat_wg[1535:1280], dat_wg[1151:896] };
  assign _0816_ = { dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt, dat_rsp_wg_sel_rt } & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15813" *) { dat_wg[1407:1152], dat_wg[1023:768], dat_wg[639:384], dat_wg[255:0] };
  assign _0817_ = { dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb, dat_rsp_wg_sel_rb } & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15814" *) { dat_wg[2175:1920], dat_wg[1791:1536], dat_wg[1407:1152], dat_wg[1023:768] };
  assign _0818_ = { dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b } & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15856" *) { dat_rsp_wg[975:960], dat_rsp_wg[911:896], dat_rsp_wg[847:832], dat_rsp_wg[783:768], dat_rsp_wg[719:704], dat_rsp_wg[655:640], dat_rsp_wg[591:576], dat_rsp_wg[527:512], dat_rsp_wg[463:448], dat_rsp_wg[399:384], dat_rsp_wg[335:320], dat_rsp_wg[271:256], dat_rsp_wg[207:192], dat_rsp_wg[143:128], dat_rsp_wg[79:64], dat_rsp_wg[15:0] };
  assign _0819_ = { dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo } & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15857" *) { dat_rsp_wg[967], dat_rsp_wg[967], dat_rsp_wg[967], dat_rsp_wg[967], dat_rsp_wg[967], dat_rsp_wg[967], dat_rsp_wg[967], dat_rsp_wg[967], dat_rsp_wg[967:960], dat_rsp_wg[903], dat_rsp_wg[903], dat_rsp_wg[903], dat_rsp_wg[903], dat_rsp_wg[903], dat_rsp_wg[903], dat_rsp_wg[903], dat_rsp_wg[903], dat_rsp_wg[903:896], dat_rsp_wg[839], dat_rsp_wg[839], dat_rsp_wg[839], dat_rsp_wg[839], dat_rsp_wg[839], dat_rsp_wg[839], dat_rsp_wg[839], dat_rsp_wg[839], dat_rsp_wg[839:832], dat_rsp_wg[775], dat_rsp_wg[775], dat_rsp_wg[775], dat_rsp_wg[775], dat_rsp_wg[775], dat_rsp_wg[775], dat_rsp_wg[775], dat_rsp_wg[775], dat_rsp_wg[775:768], dat_rsp_wg[711], dat_rsp_wg[711], dat_rsp_wg[711], dat_rsp_wg[711], dat_rsp_wg[711], dat_rsp_wg[711], dat_rsp_wg[711], dat_rsp_wg[711], dat_rsp_wg[711:704], dat_rsp_wg[647], dat_rsp_wg[647], dat_rsp_wg[647], dat_rsp_wg[647], dat_rsp_wg[647], dat_rsp_wg[647], dat_rsp_wg[647], dat_rsp_wg[647], dat_rsp_wg[647:640], dat_rsp_wg[583], dat_rsp_wg[583], dat_rsp_wg[583], dat_rsp_wg[583], dat_rsp_wg[583], dat_rsp_wg[583], dat_rsp_wg[583], dat_rsp_wg[583], dat_rsp_wg[583:576], dat_rsp_wg[519], dat_rsp_wg[519], dat_rsp_wg[519], dat_rsp_wg[519], dat_rsp_wg[519], dat_rsp_wg[519], dat_rsp_wg[519], dat_rsp_wg[519], dat_rsp_wg[519:512], dat_rsp_wg[455], dat_rsp_wg[455], dat_rsp_wg[455], dat_rsp_wg[455], dat_rsp_wg[455], dat_rsp_wg[455], dat_rsp_wg[455], dat_rsp_wg[455], dat_rsp_wg[455:448], dat_rsp_wg[391], dat_rsp_wg[391], dat_rsp_wg[391], dat_rsp_wg[391], dat_rsp_wg[391], dat_rsp_wg[391], dat_rsp_wg[391], dat_rsp_wg[391], dat_rsp_wg[391:384], dat_rsp_wg[327], dat_rsp_wg[327], dat_rsp_wg[327], dat_rsp_wg[327], dat_rsp_wg[327], dat_rsp_wg[327], dat_rsp_wg[327], dat_rsp_wg[327], dat_rsp_wg[327:320], dat_rsp_wg[263], dat_rsp_wg[263], dat_rsp_wg[263], dat_rsp_wg[263], dat_rsp_wg[263], dat_rsp_wg[263], dat_rsp_wg[263], dat_rsp_wg[263], dat_rsp_wg[263:256], dat_rsp_wg[199], dat_rsp_wg[199], dat_rsp_wg[199], dat_rsp_wg[199], dat_rsp_wg[199], dat_rsp_wg[199], dat_rsp_wg[199], dat_rsp_wg[199], dat_rsp_wg[199:192], dat_rsp_wg[135], dat_rsp_wg[135], dat_rsp_wg[135], dat_rsp_wg[135], dat_rsp_wg[135], dat_rsp_wg[135], dat_rsp_wg[135], dat_rsp_wg[135], dat_rsp_wg[135:128], dat_rsp_wg[71], dat_rsp_wg[71], dat_rsp_wg[71], dat_rsp_wg[71], dat_rsp_wg[71], dat_rsp_wg[71], dat_rsp_wg[71], dat_rsp_wg[71], dat_rsp_wg[71:64], dat_rsp_wg[7], dat_rsp_wg[7], dat_rsp_wg[7], dat_rsp_wg[7], dat_rsp_wg[7], dat_rsp_wg[7], dat_rsp_wg[7], dat_rsp_wg[7], dat_rsp_wg[7:0] };
  assign _0820_ = { dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi } & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15858" *) { dat_rsp_wg[999], dat_rsp_wg[999], dat_rsp_wg[999], dat_rsp_wg[999], dat_rsp_wg[999], dat_rsp_wg[999], dat_rsp_wg[999], dat_rsp_wg[999], dat_rsp_wg[999:992], dat_rsp_wg[935], dat_rsp_wg[935], dat_rsp_wg[935], dat_rsp_wg[935], dat_rsp_wg[935], dat_rsp_wg[935], dat_rsp_wg[935], dat_rsp_wg[935], dat_rsp_wg[935:928], dat_rsp_wg[871], dat_rsp_wg[871], dat_rsp_wg[871], dat_rsp_wg[871], dat_rsp_wg[871], dat_rsp_wg[871], dat_rsp_wg[871], dat_rsp_wg[871], dat_rsp_wg[871:864], dat_rsp_wg[807], dat_rsp_wg[807], dat_rsp_wg[807], dat_rsp_wg[807], dat_rsp_wg[807], dat_rsp_wg[807], dat_rsp_wg[807], dat_rsp_wg[807], dat_rsp_wg[807:800], dat_rsp_wg[743], dat_rsp_wg[743], dat_rsp_wg[743], dat_rsp_wg[743], dat_rsp_wg[743], dat_rsp_wg[743], dat_rsp_wg[743], dat_rsp_wg[743], dat_rsp_wg[743:736], dat_rsp_wg[679], dat_rsp_wg[679], dat_rsp_wg[679], dat_rsp_wg[679], dat_rsp_wg[679], dat_rsp_wg[679], dat_rsp_wg[679], dat_rsp_wg[679], dat_rsp_wg[679:672], dat_rsp_wg[615], dat_rsp_wg[615], dat_rsp_wg[615], dat_rsp_wg[615], dat_rsp_wg[615], dat_rsp_wg[615], dat_rsp_wg[615], dat_rsp_wg[615], dat_rsp_wg[615:608], dat_rsp_wg[551], dat_rsp_wg[551], dat_rsp_wg[551], dat_rsp_wg[551], dat_rsp_wg[551], dat_rsp_wg[551], dat_rsp_wg[551], dat_rsp_wg[551], dat_rsp_wg[551:544], dat_rsp_wg[487], dat_rsp_wg[487], dat_rsp_wg[487], dat_rsp_wg[487], dat_rsp_wg[487], dat_rsp_wg[487], dat_rsp_wg[487], dat_rsp_wg[487], dat_rsp_wg[487:480], dat_rsp_wg[423], dat_rsp_wg[423], dat_rsp_wg[423], dat_rsp_wg[423], dat_rsp_wg[423], dat_rsp_wg[423], dat_rsp_wg[423], dat_rsp_wg[423], dat_rsp_wg[423:416], dat_rsp_wg[359], dat_rsp_wg[359], dat_rsp_wg[359], dat_rsp_wg[359], dat_rsp_wg[359], dat_rsp_wg[359], dat_rsp_wg[359], dat_rsp_wg[359], dat_rsp_wg[359:352], dat_rsp_wg[295], dat_rsp_wg[295], dat_rsp_wg[295], dat_rsp_wg[295], dat_rsp_wg[295], dat_rsp_wg[295], dat_rsp_wg[295], dat_rsp_wg[295], dat_rsp_wg[295:288], dat_rsp_wg[231], dat_rsp_wg[231], dat_rsp_wg[231], dat_rsp_wg[231], dat_rsp_wg[231], dat_rsp_wg[231], dat_rsp_wg[231], dat_rsp_wg[231], dat_rsp_wg[231:224], dat_rsp_wg[167], dat_rsp_wg[167], dat_rsp_wg[167], dat_rsp_wg[167], dat_rsp_wg[167], dat_rsp_wg[167], dat_rsp_wg[167], dat_rsp_wg[167], dat_rsp_wg[167:160], dat_rsp_wg[103], dat_rsp_wg[103], dat_rsp_wg[103], dat_rsp_wg[103], dat_rsp_wg[103], dat_rsp_wg[103], dat_rsp_wg[103], dat_rsp_wg[103], dat_rsp_wg[103:96], dat_rsp_wg[39], dat_rsp_wg[39], dat_rsp_wg[39], dat_rsp_wg[39], dat_rsp_wg[39], dat_rsp_wg[39], dat_rsp_wg[39], dat_rsp_wg[39], dat_rsp_wg[39:32] };
  assign _0821_ = { dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b } & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15868" *) { dat_rsp_wg[991:976], dat_rsp_wg[927:912], dat_rsp_wg[863:848], dat_rsp_wg[799:784], dat_rsp_wg[735:720], dat_rsp_wg[671:656], dat_rsp_wg[607:592], dat_rsp_wg[543:528], dat_rsp_wg[479:464], dat_rsp_wg[415:400], dat_rsp_wg[351:336], dat_rsp_wg[287:272], dat_rsp_wg[223:208], dat_rsp_wg[159:144], dat_rsp_wg[95:80], dat_rsp_wg[31:16] };
  assign _0822_ = { dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo } & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15869" *) { dat_rsp_wg[975], dat_rsp_wg[975], dat_rsp_wg[975], dat_rsp_wg[975], dat_rsp_wg[975], dat_rsp_wg[975], dat_rsp_wg[975], dat_rsp_wg[975], dat_rsp_wg[975:968], dat_rsp_wg[911], dat_rsp_wg[911], dat_rsp_wg[911], dat_rsp_wg[911], dat_rsp_wg[911], dat_rsp_wg[911], dat_rsp_wg[911], dat_rsp_wg[911], dat_rsp_wg[911:904], dat_rsp_wg[847], dat_rsp_wg[847], dat_rsp_wg[847], dat_rsp_wg[847], dat_rsp_wg[847], dat_rsp_wg[847], dat_rsp_wg[847], dat_rsp_wg[847], dat_rsp_wg[847:840], dat_rsp_wg[783], dat_rsp_wg[783], dat_rsp_wg[783], dat_rsp_wg[783], dat_rsp_wg[783], dat_rsp_wg[783], dat_rsp_wg[783], dat_rsp_wg[783], dat_rsp_wg[783:776], dat_rsp_wg[719], dat_rsp_wg[719], dat_rsp_wg[719], dat_rsp_wg[719], dat_rsp_wg[719], dat_rsp_wg[719], dat_rsp_wg[719], dat_rsp_wg[719], dat_rsp_wg[719:712], dat_rsp_wg[655], dat_rsp_wg[655], dat_rsp_wg[655], dat_rsp_wg[655], dat_rsp_wg[655], dat_rsp_wg[655], dat_rsp_wg[655], dat_rsp_wg[655], dat_rsp_wg[655:648], dat_rsp_wg[591], dat_rsp_wg[591], dat_rsp_wg[591], dat_rsp_wg[591], dat_rsp_wg[591], dat_rsp_wg[591], dat_rsp_wg[591], dat_rsp_wg[591], dat_rsp_wg[591:584], dat_rsp_wg[527], dat_rsp_wg[527], dat_rsp_wg[527], dat_rsp_wg[527], dat_rsp_wg[527], dat_rsp_wg[527], dat_rsp_wg[527], dat_rsp_wg[527], dat_rsp_wg[527:520], dat_rsp_wg[463], dat_rsp_wg[463], dat_rsp_wg[463], dat_rsp_wg[463], dat_rsp_wg[463], dat_rsp_wg[463], dat_rsp_wg[463], dat_rsp_wg[463], dat_rsp_wg[463:456], dat_rsp_wg[399], dat_rsp_wg[399], dat_rsp_wg[399], dat_rsp_wg[399], dat_rsp_wg[399], dat_rsp_wg[399], dat_rsp_wg[399], dat_rsp_wg[399], dat_rsp_wg[399:392], dat_rsp_wg[335], dat_rsp_wg[335], dat_rsp_wg[335], dat_rsp_wg[335], dat_rsp_wg[335], dat_rsp_wg[335], dat_rsp_wg[335], dat_rsp_wg[335], dat_rsp_wg[335:328], dat_rsp_wg[271], dat_rsp_wg[271], dat_rsp_wg[271], dat_rsp_wg[271], dat_rsp_wg[271], dat_rsp_wg[271], dat_rsp_wg[271], dat_rsp_wg[271], dat_rsp_wg[271:264], dat_rsp_wg[207], dat_rsp_wg[207], dat_rsp_wg[207], dat_rsp_wg[207], dat_rsp_wg[207], dat_rsp_wg[207], dat_rsp_wg[207], dat_rsp_wg[207], dat_rsp_wg[207:200], dat_rsp_wg[143], dat_rsp_wg[143], dat_rsp_wg[143], dat_rsp_wg[143], dat_rsp_wg[143], dat_rsp_wg[143], dat_rsp_wg[143], dat_rsp_wg[143], dat_rsp_wg[143:136], dat_rsp_wg[79], dat_rsp_wg[79], dat_rsp_wg[79], dat_rsp_wg[79], dat_rsp_wg[79], dat_rsp_wg[79], dat_rsp_wg[79], dat_rsp_wg[79], dat_rsp_wg[79:72], dat_rsp_wg[15], dat_rsp_wg[15], dat_rsp_wg[15], dat_rsp_wg[15], dat_rsp_wg[15], dat_rsp_wg[15], dat_rsp_wg[15], dat_rsp_wg[15], dat_rsp_wg[15:8] };
  assign _0823_ = { dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi } & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15870" *) { dat_rsp_wg[1007], dat_rsp_wg[1007], dat_rsp_wg[1007], dat_rsp_wg[1007], dat_rsp_wg[1007], dat_rsp_wg[1007], dat_rsp_wg[1007], dat_rsp_wg[1007], dat_rsp_wg[1007:1000], dat_rsp_wg[943], dat_rsp_wg[943], dat_rsp_wg[943], dat_rsp_wg[943], dat_rsp_wg[943], dat_rsp_wg[943], dat_rsp_wg[943], dat_rsp_wg[943], dat_rsp_wg[943:936], dat_rsp_wg[879], dat_rsp_wg[879], dat_rsp_wg[879], dat_rsp_wg[879], dat_rsp_wg[879], dat_rsp_wg[879], dat_rsp_wg[879], dat_rsp_wg[879], dat_rsp_wg[879:872], dat_rsp_wg[815], dat_rsp_wg[815], dat_rsp_wg[815], dat_rsp_wg[815], dat_rsp_wg[815], dat_rsp_wg[815], dat_rsp_wg[815], dat_rsp_wg[815], dat_rsp_wg[815:808], dat_rsp_wg[751], dat_rsp_wg[751], dat_rsp_wg[751], dat_rsp_wg[751], dat_rsp_wg[751], dat_rsp_wg[751], dat_rsp_wg[751], dat_rsp_wg[751], dat_rsp_wg[751:744], dat_rsp_wg[687], dat_rsp_wg[687], dat_rsp_wg[687], dat_rsp_wg[687], dat_rsp_wg[687], dat_rsp_wg[687], dat_rsp_wg[687], dat_rsp_wg[687], dat_rsp_wg[687:680], dat_rsp_wg[623], dat_rsp_wg[623], dat_rsp_wg[623], dat_rsp_wg[623], dat_rsp_wg[623], dat_rsp_wg[623], dat_rsp_wg[623], dat_rsp_wg[623], dat_rsp_wg[623:616], dat_rsp_wg[559], dat_rsp_wg[559], dat_rsp_wg[559], dat_rsp_wg[559], dat_rsp_wg[559], dat_rsp_wg[559], dat_rsp_wg[559], dat_rsp_wg[559], dat_rsp_wg[559:552], dat_rsp_wg[495], dat_rsp_wg[495], dat_rsp_wg[495], dat_rsp_wg[495], dat_rsp_wg[495], dat_rsp_wg[495], dat_rsp_wg[495], dat_rsp_wg[495], dat_rsp_wg[495:488], dat_rsp_wg[431], dat_rsp_wg[431], dat_rsp_wg[431], dat_rsp_wg[431], dat_rsp_wg[431], dat_rsp_wg[431], dat_rsp_wg[431], dat_rsp_wg[431], dat_rsp_wg[431:424], dat_rsp_wg[367], dat_rsp_wg[367], dat_rsp_wg[367], dat_rsp_wg[367], dat_rsp_wg[367], dat_rsp_wg[367], dat_rsp_wg[367], dat_rsp_wg[367], dat_rsp_wg[367:360], dat_rsp_wg[303], dat_rsp_wg[303], dat_rsp_wg[303], dat_rsp_wg[303], dat_rsp_wg[303], dat_rsp_wg[303], dat_rsp_wg[303], dat_rsp_wg[303], dat_rsp_wg[303:296], dat_rsp_wg[239], dat_rsp_wg[239], dat_rsp_wg[239], dat_rsp_wg[239], dat_rsp_wg[239], dat_rsp_wg[239], dat_rsp_wg[239], dat_rsp_wg[239], dat_rsp_wg[239:232], dat_rsp_wg[175], dat_rsp_wg[175], dat_rsp_wg[175], dat_rsp_wg[175], dat_rsp_wg[175], dat_rsp_wg[175], dat_rsp_wg[175], dat_rsp_wg[175], dat_rsp_wg[175:168], dat_rsp_wg[111], dat_rsp_wg[111], dat_rsp_wg[111], dat_rsp_wg[111], dat_rsp_wg[111], dat_rsp_wg[111], dat_rsp_wg[111], dat_rsp_wg[111], dat_rsp_wg[111:104], dat_rsp_wg[47], dat_rsp_wg[47], dat_rsp_wg[47], dat_rsp_wg[47], dat_rsp_wg[47], dat_rsp_wg[47], dat_rsp_wg[47], dat_rsp_wg[47], dat_rsp_wg[47:40] };
  assign _0824_ = { dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b } & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15880" *) { dat_rsp_wg[1007:992], dat_rsp_wg[943:928], dat_rsp_wg[879:864], dat_rsp_wg[815:800], dat_rsp_wg[751:736], dat_rsp_wg[687:672], dat_rsp_wg[623:608], dat_rsp_wg[559:544], dat_rsp_wg[495:480], dat_rsp_wg[431:416], dat_rsp_wg[367:352], dat_rsp_wg[303:288], dat_rsp_wg[239:224], dat_rsp_wg[175:160], dat_rsp_wg[111:96], dat_rsp_wg[47:32] };
  assign _0825_ = { dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo } & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15881" *) { dat_rsp_wg[983], dat_rsp_wg[983], dat_rsp_wg[983], dat_rsp_wg[983], dat_rsp_wg[983], dat_rsp_wg[983], dat_rsp_wg[983], dat_rsp_wg[983], dat_rsp_wg[983:976], dat_rsp_wg[919], dat_rsp_wg[919], dat_rsp_wg[919], dat_rsp_wg[919], dat_rsp_wg[919], dat_rsp_wg[919], dat_rsp_wg[919], dat_rsp_wg[919], dat_rsp_wg[919:912], dat_rsp_wg[855], dat_rsp_wg[855], dat_rsp_wg[855], dat_rsp_wg[855], dat_rsp_wg[855], dat_rsp_wg[855], dat_rsp_wg[855], dat_rsp_wg[855], dat_rsp_wg[855:848], dat_rsp_wg[791], dat_rsp_wg[791], dat_rsp_wg[791], dat_rsp_wg[791], dat_rsp_wg[791], dat_rsp_wg[791], dat_rsp_wg[791], dat_rsp_wg[791], dat_rsp_wg[791:784], dat_rsp_wg[727], dat_rsp_wg[727], dat_rsp_wg[727], dat_rsp_wg[727], dat_rsp_wg[727], dat_rsp_wg[727], dat_rsp_wg[727], dat_rsp_wg[727], dat_rsp_wg[727:720], dat_rsp_wg[663], dat_rsp_wg[663], dat_rsp_wg[663], dat_rsp_wg[663], dat_rsp_wg[663], dat_rsp_wg[663], dat_rsp_wg[663], dat_rsp_wg[663], dat_rsp_wg[663:656], dat_rsp_wg[599], dat_rsp_wg[599], dat_rsp_wg[599], dat_rsp_wg[599], dat_rsp_wg[599], dat_rsp_wg[599], dat_rsp_wg[599], dat_rsp_wg[599], dat_rsp_wg[599:592], dat_rsp_wg[535], dat_rsp_wg[535], dat_rsp_wg[535], dat_rsp_wg[535], dat_rsp_wg[535], dat_rsp_wg[535], dat_rsp_wg[535], dat_rsp_wg[535], dat_rsp_wg[535:528], dat_rsp_wg[471], dat_rsp_wg[471], dat_rsp_wg[471], dat_rsp_wg[471], dat_rsp_wg[471], dat_rsp_wg[471], dat_rsp_wg[471], dat_rsp_wg[471], dat_rsp_wg[471:464], dat_rsp_wg[407], dat_rsp_wg[407], dat_rsp_wg[407], dat_rsp_wg[407], dat_rsp_wg[407], dat_rsp_wg[407], dat_rsp_wg[407], dat_rsp_wg[407], dat_rsp_wg[407:400], dat_rsp_wg[343], dat_rsp_wg[343], dat_rsp_wg[343], dat_rsp_wg[343], dat_rsp_wg[343], dat_rsp_wg[343], dat_rsp_wg[343], dat_rsp_wg[343], dat_rsp_wg[343:336], dat_rsp_wg[279], dat_rsp_wg[279], dat_rsp_wg[279], dat_rsp_wg[279], dat_rsp_wg[279], dat_rsp_wg[279], dat_rsp_wg[279], dat_rsp_wg[279], dat_rsp_wg[279:272], dat_rsp_wg[215], dat_rsp_wg[215], dat_rsp_wg[215], dat_rsp_wg[215], dat_rsp_wg[215], dat_rsp_wg[215], dat_rsp_wg[215], dat_rsp_wg[215], dat_rsp_wg[215:208], dat_rsp_wg[151], dat_rsp_wg[151], dat_rsp_wg[151], dat_rsp_wg[151], dat_rsp_wg[151], dat_rsp_wg[151], dat_rsp_wg[151], dat_rsp_wg[151], dat_rsp_wg[151:144], dat_rsp_wg[87], dat_rsp_wg[87], dat_rsp_wg[87], dat_rsp_wg[87], dat_rsp_wg[87], dat_rsp_wg[87], dat_rsp_wg[87], dat_rsp_wg[87], dat_rsp_wg[87:80], dat_rsp_wg[23], dat_rsp_wg[23], dat_rsp_wg[23], dat_rsp_wg[23], dat_rsp_wg[23], dat_rsp_wg[23], dat_rsp_wg[23], dat_rsp_wg[23], dat_rsp_wg[23:16] };
  assign _0826_ = { dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi } & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15882" *) { dat_rsp_wg[1015], dat_rsp_wg[1015], dat_rsp_wg[1015], dat_rsp_wg[1015], dat_rsp_wg[1015], dat_rsp_wg[1015], dat_rsp_wg[1015], dat_rsp_wg[1015], dat_rsp_wg[1015:1008], dat_rsp_wg[951], dat_rsp_wg[951], dat_rsp_wg[951], dat_rsp_wg[951], dat_rsp_wg[951], dat_rsp_wg[951], dat_rsp_wg[951], dat_rsp_wg[951], dat_rsp_wg[951:944], dat_rsp_wg[887], dat_rsp_wg[887], dat_rsp_wg[887], dat_rsp_wg[887], dat_rsp_wg[887], dat_rsp_wg[887], dat_rsp_wg[887], dat_rsp_wg[887], dat_rsp_wg[887:880], dat_rsp_wg[823], dat_rsp_wg[823], dat_rsp_wg[823], dat_rsp_wg[823], dat_rsp_wg[823], dat_rsp_wg[823], dat_rsp_wg[823], dat_rsp_wg[823], dat_rsp_wg[823:816], dat_rsp_wg[759], dat_rsp_wg[759], dat_rsp_wg[759], dat_rsp_wg[759], dat_rsp_wg[759], dat_rsp_wg[759], dat_rsp_wg[759], dat_rsp_wg[759], dat_rsp_wg[759:752], dat_rsp_wg[695], dat_rsp_wg[695], dat_rsp_wg[695], dat_rsp_wg[695], dat_rsp_wg[695], dat_rsp_wg[695], dat_rsp_wg[695], dat_rsp_wg[695], dat_rsp_wg[695:688], dat_rsp_wg[631], dat_rsp_wg[631], dat_rsp_wg[631], dat_rsp_wg[631], dat_rsp_wg[631], dat_rsp_wg[631], dat_rsp_wg[631], dat_rsp_wg[631], dat_rsp_wg[631:624], dat_rsp_wg[567], dat_rsp_wg[567], dat_rsp_wg[567], dat_rsp_wg[567], dat_rsp_wg[567], dat_rsp_wg[567], dat_rsp_wg[567], dat_rsp_wg[567], dat_rsp_wg[567:560], dat_rsp_wg[503], dat_rsp_wg[503], dat_rsp_wg[503], dat_rsp_wg[503], dat_rsp_wg[503], dat_rsp_wg[503], dat_rsp_wg[503], dat_rsp_wg[503], dat_rsp_wg[503:496], dat_rsp_wg[439], dat_rsp_wg[439], dat_rsp_wg[439], dat_rsp_wg[439], dat_rsp_wg[439], dat_rsp_wg[439], dat_rsp_wg[439], dat_rsp_wg[439], dat_rsp_wg[439:432], dat_rsp_wg[375], dat_rsp_wg[375], dat_rsp_wg[375], dat_rsp_wg[375], dat_rsp_wg[375], dat_rsp_wg[375], dat_rsp_wg[375], dat_rsp_wg[375], dat_rsp_wg[375:368], dat_rsp_wg[311], dat_rsp_wg[311], dat_rsp_wg[311], dat_rsp_wg[311], dat_rsp_wg[311], dat_rsp_wg[311], dat_rsp_wg[311], dat_rsp_wg[311], dat_rsp_wg[311:304], dat_rsp_wg[247], dat_rsp_wg[247], dat_rsp_wg[247], dat_rsp_wg[247], dat_rsp_wg[247], dat_rsp_wg[247], dat_rsp_wg[247], dat_rsp_wg[247], dat_rsp_wg[247:240], dat_rsp_wg[183], dat_rsp_wg[183], dat_rsp_wg[183], dat_rsp_wg[183], dat_rsp_wg[183], dat_rsp_wg[183], dat_rsp_wg[183], dat_rsp_wg[183], dat_rsp_wg[183:176], dat_rsp_wg[119], dat_rsp_wg[119], dat_rsp_wg[119], dat_rsp_wg[119], dat_rsp_wg[119], dat_rsp_wg[119], dat_rsp_wg[119], dat_rsp_wg[119], dat_rsp_wg[119:112], dat_rsp_wg[55], dat_rsp_wg[55], dat_rsp_wg[55], dat_rsp_wg[55], dat_rsp_wg[55], dat_rsp_wg[55], dat_rsp_wg[55], dat_rsp_wg[55], dat_rsp_wg[55:48] };
  assign _0827_ = { dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b, dat_rsp_wg_sel_16b } & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15892" *) { dat_rsp_wg[1023:1008], dat_rsp_wg[959:944], dat_rsp_wg[895:880], dat_rsp_wg[831:816], dat_rsp_wg[767:752], dat_rsp_wg[703:688], dat_rsp_wg[639:624], dat_rsp_wg[575:560], dat_rsp_wg[511:496], dat_rsp_wg[447:432], dat_rsp_wg[383:368], dat_rsp_wg[319:304], dat_rsp_wg[255:240], dat_rsp_wg[191:176], dat_rsp_wg[127:112], dat_rsp_wg[63:48] };
  assign _0828_ = { dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo, dat_rsp_wg_sel_8b_lo } & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15893" *) { dat_rsp_wg[991], dat_rsp_wg[991], dat_rsp_wg[991], dat_rsp_wg[991], dat_rsp_wg[991], dat_rsp_wg[991], dat_rsp_wg[991], dat_rsp_wg[991], dat_rsp_wg[991:984], dat_rsp_wg[927], dat_rsp_wg[927], dat_rsp_wg[927], dat_rsp_wg[927], dat_rsp_wg[927], dat_rsp_wg[927], dat_rsp_wg[927], dat_rsp_wg[927], dat_rsp_wg[927:920], dat_rsp_wg[863], dat_rsp_wg[863], dat_rsp_wg[863], dat_rsp_wg[863], dat_rsp_wg[863], dat_rsp_wg[863], dat_rsp_wg[863], dat_rsp_wg[863], dat_rsp_wg[863:856], dat_rsp_wg[799], dat_rsp_wg[799], dat_rsp_wg[799], dat_rsp_wg[799], dat_rsp_wg[799], dat_rsp_wg[799], dat_rsp_wg[799], dat_rsp_wg[799], dat_rsp_wg[799:792], dat_rsp_wg[735], dat_rsp_wg[735], dat_rsp_wg[735], dat_rsp_wg[735], dat_rsp_wg[735], dat_rsp_wg[735], dat_rsp_wg[735], dat_rsp_wg[735], dat_rsp_wg[735:728], dat_rsp_wg[671], dat_rsp_wg[671], dat_rsp_wg[671], dat_rsp_wg[671], dat_rsp_wg[671], dat_rsp_wg[671], dat_rsp_wg[671], dat_rsp_wg[671], dat_rsp_wg[671:664], dat_rsp_wg[607], dat_rsp_wg[607], dat_rsp_wg[607], dat_rsp_wg[607], dat_rsp_wg[607], dat_rsp_wg[607], dat_rsp_wg[607], dat_rsp_wg[607], dat_rsp_wg[607:600], dat_rsp_wg[543], dat_rsp_wg[543], dat_rsp_wg[543], dat_rsp_wg[543], dat_rsp_wg[543], dat_rsp_wg[543], dat_rsp_wg[543], dat_rsp_wg[543], dat_rsp_wg[543:536], dat_rsp_wg[479], dat_rsp_wg[479], dat_rsp_wg[479], dat_rsp_wg[479], dat_rsp_wg[479], dat_rsp_wg[479], dat_rsp_wg[479], dat_rsp_wg[479], dat_rsp_wg[479:472], dat_rsp_wg[415], dat_rsp_wg[415], dat_rsp_wg[415], dat_rsp_wg[415], dat_rsp_wg[415], dat_rsp_wg[415], dat_rsp_wg[415], dat_rsp_wg[415], dat_rsp_wg[415:408], dat_rsp_wg[351], dat_rsp_wg[351], dat_rsp_wg[351], dat_rsp_wg[351], dat_rsp_wg[351], dat_rsp_wg[351], dat_rsp_wg[351], dat_rsp_wg[351], dat_rsp_wg[351:344], dat_rsp_wg[287], dat_rsp_wg[287], dat_rsp_wg[287], dat_rsp_wg[287], dat_rsp_wg[287], dat_rsp_wg[287], dat_rsp_wg[287], dat_rsp_wg[287], dat_rsp_wg[287:280], dat_rsp_wg[223], dat_rsp_wg[223], dat_rsp_wg[223], dat_rsp_wg[223], dat_rsp_wg[223], dat_rsp_wg[223], dat_rsp_wg[223], dat_rsp_wg[223], dat_rsp_wg[223:216], dat_rsp_wg[159], dat_rsp_wg[159], dat_rsp_wg[159], dat_rsp_wg[159], dat_rsp_wg[159], dat_rsp_wg[159], dat_rsp_wg[159], dat_rsp_wg[159], dat_rsp_wg[159:152], dat_rsp_wg[95], dat_rsp_wg[95], dat_rsp_wg[95], dat_rsp_wg[95], dat_rsp_wg[95], dat_rsp_wg[95], dat_rsp_wg[95], dat_rsp_wg[95], dat_rsp_wg[95:88], dat_rsp_wg[31], dat_rsp_wg[31], dat_rsp_wg[31], dat_rsp_wg[31], dat_rsp_wg[31], dat_rsp_wg[31], dat_rsp_wg[31], dat_rsp_wg[31], dat_rsp_wg[31:24] };
  assign _0829_ = { dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi, dat_rsp_wg_sel_8b_hi } & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15894" *) { dat_rsp_wg[1023], dat_rsp_wg[1023], dat_rsp_wg[1023], dat_rsp_wg[1023], dat_rsp_wg[1023], dat_rsp_wg[1023], dat_rsp_wg[1023], dat_rsp_wg[1023], dat_rsp_wg[1023:1016], dat_rsp_wg[959], dat_rsp_wg[959], dat_rsp_wg[959], dat_rsp_wg[959], dat_rsp_wg[959], dat_rsp_wg[959], dat_rsp_wg[959], dat_rsp_wg[959], dat_rsp_wg[959:952], dat_rsp_wg[895], dat_rsp_wg[895], dat_rsp_wg[895], dat_rsp_wg[895], dat_rsp_wg[895], dat_rsp_wg[895], dat_rsp_wg[895], dat_rsp_wg[895], dat_rsp_wg[895:888], dat_rsp_wg[831], dat_rsp_wg[831], dat_rsp_wg[831], dat_rsp_wg[831], dat_rsp_wg[831], dat_rsp_wg[831], dat_rsp_wg[831], dat_rsp_wg[831], dat_rsp_wg[831:824], dat_rsp_wg[767], dat_rsp_wg[767], dat_rsp_wg[767], dat_rsp_wg[767], dat_rsp_wg[767], dat_rsp_wg[767], dat_rsp_wg[767], dat_rsp_wg[767], dat_rsp_wg[767:760], dat_rsp_wg[703], dat_rsp_wg[703], dat_rsp_wg[703], dat_rsp_wg[703], dat_rsp_wg[703], dat_rsp_wg[703], dat_rsp_wg[703], dat_rsp_wg[703], dat_rsp_wg[703:696], dat_rsp_wg[639], dat_rsp_wg[639], dat_rsp_wg[639], dat_rsp_wg[639], dat_rsp_wg[639], dat_rsp_wg[639], dat_rsp_wg[639], dat_rsp_wg[639], dat_rsp_wg[639:632], dat_rsp_wg[575], dat_rsp_wg[575], dat_rsp_wg[575], dat_rsp_wg[575], dat_rsp_wg[575], dat_rsp_wg[575], dat_rsp_wg[575], dat_rsp_wg[575], dat_rsp_wg[575:568], dat_rsp_wg[511], dat_rsp_wg[511], dat_rsp_wg[511], dat_rsp_wg[511], dat_rsp_wg[511], dat_rsp_wg[511], dat_rsp_wg[511], dat_rsp_wg[511], dat_rsp_wg[511:504], dat_rsp_wg[447], dat_rsp_wg[447], dat_rsp_wg[447], dat_rsp_wg[447], dat_rsp_wg[447], dat_rsp_wg[447], dat_rsp_wg[447], dat_rsp_wg[447], dat_rsp_wg[447:440], dat_rsp_wg[383], dat_rsp_wg[383], dat_rsp_wg[383], dat_rsp_wg[383], dat_rsp_wg[383], dat_rsp_wg[383], dat_rsp_wg[383], dat_rsp_wg[383], dat_rsp_wg[383:376], dat_rsp_wg[319], dat_rsp_wg[319], dat_rsp_wg[319], dat_rsp_wg[319], dat_rsp_wg[319], dat_rsp_wg[319], dat_rsp_wg[319], dat_rsp_wg[319], dat_rsp_wg[319:312], dat_rsp_wg[255], dat_rsp_wg[255], dat_rsp_wg[255], dat_rsp_wg[255], dat_rsp_wg[255], dat_rsp_wg[255], dat_rsp_wg[255], dat_rsp_wg[255], dat_rsp_wg[255:248], dat_rsp_wg[191], dat_rsp_wg[191], dat_rsp_wg[191], dat_rsp_wg[191], dat_rsp_wg[191], dat_rsp_wg[191], dat_rsp_wg[191], dat_rsp_wg[191], dat_rsp_wg[191:184], dat_rsp_wg[127], dat_rsp_wg[127], dat_rsp_wg[127], dat_rsp_wg[127], dat_rsp_wg[127], dat_rsp_wg[127], dat_rsp_wg[127], dat_rsp_wg[127], dat_rsp_wg[127:120], dat_rsp_wg[63], dat_rsp_wg[63], dat_rsp_wg[63], dat_rsp_wg[63], dat_rsp_wg[63], dat_rsp_wg[63], dat_rsp_wg[63], dat_rsp_wg[63], dat_rsp_wg[63:56] };
  assign _0830_ = _1072_ & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15961" *) _1071_;
  assign _0831_ = _0830_ & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15961" *) _1038_;
  assign _0832_ = _0830_ & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15962" *) dat_rsp_pd[0];
  assign _0833_ = _1073_ & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15963" *) _1039_;
  assign _0834_ = _1073_ & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15964" *) _1040_;
  assign _0835_ = _1073_ & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15965" *) _1041_;
  assign _0836_ = _1073_ & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15966" *) _1042_;
  assign _0837_ = _1073_ & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15981" *) dat_rsp_pd[4];
  assign _0838_ = dat_rsp_pd[0] & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15986" *) dat_rsp_pd[5];
  assign dat_rsp_sft_lo_d1_en = dat_rsp_pvld_d1 & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16140" *) _1077_;
  assign dat_rsp_sft_hi_d1_en = dat_rsp_sft_lo_d1_en & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16141" *) _1106_;
  assign dat_rsp_sft_lo_d2_en = dat_rsp_pvld_d2 & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16142" *) _1047_;
  assign dat_rsp_sft_hi_d2_en = dat_rsp_sft_lo_d2_en & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16143" *) _1107_;
  assign dat_rsp_sft_lo_d3_en = dat_rsp_pvld_d3 & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16144" *) _1047_;
  assign dat_rsp_sft_hi_d3_en = dat_rsp_sft_lo_d3_en & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16145" *) _1108_;
  assign _0839_ = { dat_rsp_ori_mask[31:0], dat_rsp_ori_mask[31:0], dat_rsp_ori_mask[31:0], dat_rsp_ori_mask[31:0] } & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16302" *) { dat_rsp_cur_h_mask_p3, dat_rsp_cur_h_mask_p2, dat_rsp_cur_h_mask_p1[31:0], 32'b11111111111111111111111111111111 };
  assign _0840_ = { dat_rsp_ori_mask[63:0], dat_rsp_ori_mask[63:0] } & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16303" *) { dat_rsp_cur_h_mask_p1, 64'b1111111111111111111111111111111111111111111111111111111111111111 };
  assign _0841_ = { dat_rsp_ori_mask[15:0], dat_rsp_ori_mask[15:0], dat_rsp_ori_mask[15:0], dat_rsp_ori_mask[15:0] } & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16312" *) { dat_rsp_cur_h_mask_p3[15:0], dat_rsp_cur_h_mask_p2[15:0], dat_rsp_cur_h_mask_p1[15:0], 16'b1111111111111111 };
  assign _0842_ = { dat_rsp_ori_mask[31:0], dat_rsp_ori_mask[31:0] } & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16313" *) { dat_rsp_cur_h_mask_p1[31:0], 32'b11111111111111111111111111111111 };
  assign _0843_ = dat_rsp_mask_8b & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16369" *) dat_rsp_mask_val_int8;
  assign _0844_ = dat_rsp_mask_16b & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16370" *) { dat_rsp_mask_val_fp16[127], dat_rsp_mask_val_fp16[127], dat_rsp_mask_val_fp16[125], dat_rsp_mask_val_fp16[125], dat_rsp_mask_val_fp16[123], dat_rsp_mask_val_fp16[123], dat_rsp_mask_val_fp16[121], dat_rsp_mask_val_fp16[121], dat_rsp_mask_val_fp16[119], dat_rsp_mask_val_fp16[119], dat_rsp_mask_val_fp16[117], dat_rsp_mask_val_fp16[117], dat_rsp_mask_val_fp16[115], dat_rsp_mask_val_fp16[115], dat_rsp_mask_val_fp16[113], dat_rsp_mask_val_fp16[113], dat_rsp_mask_val_fp16[111], dat_rsp_mask_val_fp16[111], dat_rsp_mask_val_fp16[109], dat_rsp_mask_val_fp16[109], dat_rsp_mask_val_fp16[107], dat_rsp_mask_val_fp16[107], dat_rsp_mask_val_fp16[105], dat_rsp_mask_val_fp16[105], dat_rsp_mask_val_fp16[103], dat_rsp_mask_val_fp16[103], dat_rsp_mask_val_fp16[101], dat_rsp_mask_val_fp16[101], dat_rsp_mask_val_fp16[99], dat_rsp_mask_val_fp16[99], dat_rsp_mask_val_fp16[97], dat_rsp_mask_val_fp16[97], dat_rsp_mask_val_fp16[95], dat_rsp_mask_val_fp16[95], dat_rsp_mask_val_fp16[93], dat_rsp_mask_val_fp16[93], dat_rsp_mask_val_fp16[91], dat_rsp_mask_val_fp16[91], dat_rsp_mask_val_fp16[89], dat_rsp_mask_val_fp16[89], dat_rsp_mask_val_fp16[87], dat_rsp_mask_val_fp16[87], dat_rsp_mask_val_fp16[85], dat_rsp_mask_val_fp16[85], dat_rsp_mask_val_fp16[83], dat_rsp_mask_val_fp16[83], dat_rsp_mask_val_fp16[81], dat_rsp_mask_val_fp16[81], dat_rsp_mask_val_fp16[79], dat_rsp_mask_val_fp16[79], dat_rsp_mask_val_fp16[77], dat_rsp_mask_val_fp16[77], dat_rsp_mask_val_fp16[75], dat_rsp_mask_val_fp16[75], dat_rsp_mask_val_fp16[73], dat_rsp_mask_val_fp16[73], dat_rsp_mask_val_fp16[71], dat_rsp_mask_val_fp16[71], dat_rsp_mask_val_fp16[69], dat_rsp_mask_val_fp16[69], dat_rsp_mask_val_fp16[67], dat_rsp_mask_val_fp16[67], dat_rsp_mask_val_fp16[65], dat_rsp_mask_val_fp16[65], dat_rsp_mask_val_fp16[63], dat_rsp_mask_val_fp16[63], dat_rsp_mask_val_fp16[61], dat_rsp_mask_val_fp16[61], dat_rsp_mask_val_fp16[59], dat_rsp_mask_val_fp16[59], dat_rsp_mask_val_fp16[57], dat_rsp_mask_val_fp16[57], dat_rsp_mask_val_fp16[55], dat_rsp_mask_val_fp16[55], dat_rsp_mask_val_fp16[53], dat_rsp_mask_val_fp16[53], dat_rsp_mask_val_fp16[51], dat_rsp_mask_val_fp16[51], dat_rsp_mask_val_fp16[49], dat_rsp_mask_val_fp16[49], dat_rsp_mask_val_fp16[47], dat_rsp_mask_val_fp16[47], dat_rsp_mask_val_fp16[45], dat_rsp_mask_val_fp16[45], dat_rsp_mask_val_fp16[43], dat_rsp_mask_val_fp16[43], dat_rsp_mask_val_fp16[41], dat_rsp_mask_val_fp16[41], dat_rsp_mask_val_fp16[39], dat_rsp_mask_val_fp16[39], dat_rsp_mask_val_fp16[37], dat_rsp_mask_val_fp16[37], dat_rsp_mask_val_fp16[35], dat_rsp_mask_val_fp16[35], dat_rsp_mask_val_fp16[33], dat_rsp_mask_val_fp16[33], dat_rsp_mask_val_fp16[31], dat_rsp_mask_val_fp16[31], dat_rsp_mask_val_fp16[29], dat_rsp_mask_val_fp16[29], dat_rsp_mask_val_fp16[27], dat_rsp_mask_val_fp16[27], dat_rsp_mask_val_fp16[25], dat_rsp_mask_val_fp16[25], dat_rsp_mask_val_fp16[23], dat_rsp_mask_val_fp16[23], dat_rsp_mask_val_fp16[21], dat_rsp_mask_val_fp16[21], dat_rsp_mask_val_fp16[19], dat_rsp_mask_val_fp16[19], dat_rsp_mask_val_fp16[17], dat_rsp_mask_val_fp16[17], dat_rsp_mask_val_fp16[15], dat_rsp_mask_val_fp16[15], dat_rsp_mask_val_fp16[13], dat_rsp_mask_val_fp16[13], dat_rsp_mask_val_fp16[11], dat_rsp_mask_val_fp16[11], dat_rsp_mask_val_fp16[9], dat_rsp_mask_val_fp16[9], dat_rsp_mask_val_fp16[7], dat_rsp_mask_val_fp16[7], dat_rsp_mask_val_fp16[5], dat_rsp_mask_val_fp16[5], dat_rsp_mask_val_fp16[3], dat_rsp_mask_val_fp16[3], dat_rsp_mask_val_fp16[1], dat_rsp_mask_val_fp16[1] };
  assign _0845_ = dat_rsp_mask_16b & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16371" *) { dat_rsp_mask_val_int16[127], dat_rsp_mask_val_int16[127], dat_rsp_mask_val_int16[125], dat_rsp_mask_val_int16[125], dat_rsp_mask_val_int16[123], dat_rsp_mask_val_int16[123], dat_rsp_mask_val_int16[121], dat_rsp_mask_val_int16[121], dat_rsp_mask_val_int16[119], dat_rsp_mask_val_int16[119], dat_rsp_mask_val_int16[117], dat_rsp_mask_val_int16[117], dat_rsp_mask_val_int16[115], dat_rsp_mask_val_int16[115], dat_rsp_mask_val_int16[113], dat_rsp_mask_val_int16[113], dat_rsp_mask_val_int16[111], dat_rsp_mask_val_int16[111], dat_rsp_mask_val_int16[109], dat_rsp_mask_val_int16[109], dat_rsp_mask_val_int16[107], dat_rsp_mask_val_int16[107], dat_rsp_mask_val_int16[105], dat_rsp_mask_val_int16[105], dat_rsp_mask_val_int16[103], dat_rsp_mask_val_int16[103], dat_rsp_mask_val_int16[101], dat_rsp_mask_val_int16[101], dat_rsp_mask_val_int16[99], dat_rsp_mask_val_int16[99], dat_rsp_mask_val_int16[97], dat_rsp_mask_val_int16[97], dat_rsp_mask_val_int16[95], dat_rsp_mask_val_int16[95], dat_rsp_mask_val_int16[93], dat_rsp_mask_val_int16[93], dat_rsp_mask_val_int16[91], dat_rsp_mask_val_int16[91], dat_rsp_mask_val_int16[89], dat_rsp_mask_val_int16[89], dat_rsp_mask_val_int16[87], dat_rsp_mask_val_int16[87], dat_rsp_mask_val_int16[85], dat_rsp_mask_val_int16[85], dat_rsp_mask_val_int16[83], dat_rsp_mask_val_int16[83], dat_rsp_mask_val_int16[81], dat_rsp_mask_val_int16[81], dat_rsp_mask_val_int16[79], dat_rsp_mask_val_int16[79], dat_rsp_mask_val_int16[77], dat_rsp_mask_val_int16[77], dat_rsp_mask_val_int16[75], dat_rsp_mask_val_int16[75], dat_rsp_mask_val_int16[73], dat_rsp_mask_val_int16[73], dat_rsp_mask_val_int16[71], dat_rsp_mask_val_int16[71], dat_rsp_mask_val_int16[69], dat_rsp_mask_val_int16[69], dat_rsp_mask_val_int16[67], dat_rsp_mask_val_int16[67], dat_rsp_mask_val_int16[65], dat_rsp_mask_val_int16[65], dat_rsp_mask_val_int16[63], dat_rsp_mask_val_int16[63], dat_rsp_mask_val_int16[61], dat_rsp_mask_val_int16[61], dat_rsp_mask_val_int16[59], dat_rsp_mask_val_int16[59], dat_rsp_mask_val_int16[57], dat_rsp_mask_val_int16[57], dat_rsp_mask_val_int16[55], dat_rsp_mask_val_int16[55], dat_rsp_mask_val_int16[53], dat_rsp_mask_val_int16[53], dat_rsp_mask_val_int16[51], dat_rsp_mask_val_int16[51], dat_rsp_mask_val_int16[49], dat_rsp_mask_val_int16[49], dat_rsp_mask_val_int16[47], dat_rsp_mask_val_int16[47], dat_rsp_mask_val_int16[45], dat_rsp_mask_val_int16[45], dat_rsp_mask_val_int16[43], dat_rsp_mask_val_int16[43], dat_rsp_mask_val_int16[41], dat_rsp_mask_val_int16[41], dat_rsp_mask_val_int16[39], dat_rsp_mask_val_int16[39], dat_rsp_mask_val_int16[37], dat_rsp_mask_val_int16[37], dat_rsp_mask_val_int16[35], dat_rsp_mask_val_int16[35], dat_rsp_mask_val_int16[33], dat_rsp_mask_val_int16[33], dat_rsp_mask_val_int16[31], dat_rsp_mask_val_int16[31], dat_rsp_mask_val_int16[29], dat_rsp_mask_val_int16[29], dat_rsp_mask_val_int16[27], dat_rsp_mask_val_int16[27], dat_rsp_mask_val_int16[25], dat_rsp_mask_val_int16[25], dat_rsp_mask_val_int16[23], dat_rsp_mask_val_int16[23], dat_rsp_mask_val_int16[21], dat_rsp_mask_val_int16[21], dat_rsp_mask_val_int16[19], dat_rsp_mask_val_int16[19], dat_rsp_mask_val_int16[17], dat_rsp_mask_val_int16[17], dat_rsp_mask_val_int16[15], dat_rsp_mask_val_int16[15], dat_rsp_mask_val_int16[13], dat_rsp_mask_val_int16[13], dat_rsp_mask_val_int16[11], dat_rsp_mask_val_int16[11], dat_rsp_mask_val_int16[9], dat_rsp_mask_val_int16[9], dat_rsp_mask_val_int16[7], dat_rsp_mask_val_int16[7], dat_rsp_mask_val_int16[5], dat_rsp_mask_val_int16[5], dat_rsp_mask_val_int16[3], dat_rsp_mask_val_int16[3], dat_rsp_mask_val_int16[1], dat_rsp_mask_val_int16[1] };
  assign _0846_ = _1109_ & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16378" *) dat_rsp_pvld;
  assign dat_out_bypass_p1_vld_w = _0846_ & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16378" *) _1110_;
  assign dat_out_bypass_p0_vld_w = dat_rsp_pvld & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16379" *) _1111_;
  assign _0847_ = dat_out_bypass_p0_vld_w & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16923" *) dat_out_bypass_mask_w[0];
  assign _0848_ = dat_out_bypass_p0_vld_w & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16933" *) dat_out_bypass_mask_w[1];
  assign _0849_ = dat_out_bypass_p0_vld_w & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16943" *) dat_out_bypass_mask_w[2];
  assign _0850_ = dat_out_bypass_p0_vld_w & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16953" *) dat_out_bypass_mask_w[3];
  assign _0851_ = dat_out_bypass_p0_vld_w & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16963" *) dat_out_bypass_mask_w[4];
  assign _0852_ = dat_out_bypass_p0_vld_w & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16973" *) dat_out_bypass_mask_w[5];
  assign _0853_ = dat_out_bypass_p0_vld_w & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16983" *) dat_out_bypass_mask_w[6];
  assign _0854_ = dat_out_bypass_p0_vld_w & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16993" *) dat_out_bypass_mask_w[7];
  assign _0855_ = dat_out_bypass_p0_vld_w & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17003" *) dat_out_bypass_mask_w[8];
  assign _0856_ = dat_out_bypass_p0_vld_w & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17013" *) dat_out_bypass_mask_w[9];
  assign _0857_ = dat_out_bypass_p0_vld_w & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17023" *) dat_out_bypass_mask_w[10];
  assign _0858_ = dat_out_bypass_p0_vld_w & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17033" *) dat_out_bypass_mask_w[11];
  assign _0859_ = dat_out_bypass_p0_vld_w & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17043" *) dat_out_bypass_mask_w[12];
  assign _0860_ = dat_out_bypass_p0_vld_w & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17053" *) dat_out_bypass_mask_w[13];
  assign _0861_ = dat_out_bypass_p0_vld_w & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17063" *) dat_out_bypass_mask_w[14];
  assign _0862_ = dat_out_bypass_p0_vld_w & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17073" *) dat_out_bypass_mask_w[15];
  assign _0863_ = dat_out_bypass_p0_vld_w & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17083" *) dat_out_bypass_mask_w[16];
  assign _0864_ = dat_out_bypass_p0_vld_w & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17093" *) dat_out_bypass_mask_w[17];
  assign _0865_ = dat_out_bypass_p0_vld_w & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17103" *) dat_out_bypass_mask_w[18];
  assign _0866_ = dat_out_bypass_p0_vld_w & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17113" *) dat_out_bypass_mask_w[19];
  assign _0867_ = dat_out_bypass_p0_vld_w & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17123" *) dat_out_bypass_mask_w[20];
  assign _0868_ = dat_out_bypass_p0_vld_w & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17133" *) dat_out_bypass_mask_w[21];
  assign _0869_ = dat_out_bypass_p0_vld_w & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17143" *) dat_out_bypass_mask_w[22];
  assign _0870_ = dat_out_bypass_p0_vld_w & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17153" *) dat_out_bypass_mask_w[23];
  assign _0871_ = dat_out_bypass_p0_vld_w & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17163" *) dat_out_bypass_mask_w[24];
  assign _0872_ = dat_out_bypass_p0_vld_w & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17173" *) dat_out_bypass_mask_w[25];
  assign _0873_ = dat_out_bypass_p0_vld_w & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17183" *) dat_out_bypass_mask_w[26];
  assign _0874_ = dat_out_bypass_p0_vld_w & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17193" *) dat_out_bypass_mask_w[27];
  assign _0875_ = dat_out_bypass_p0_vld_w & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17203" *) dat_out_bypass_mask_w[28];
  assign _0876_ = dat_out_bypass_p0_vld_w & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17213" *) dat_out_bypass_mask_w[29];
  assign _0877_ = dat_out_bypass_p0_vld_w & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17223" *) dat_out_bypass_mask_w[30];
  assign _0878_ = dat_out_bypass_p0_vld_w & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17233" *) dat_out_bypass_mask_w[31];
  assign _0879_ = dat_out_bypass_p0_vld_w & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17243" *) dat_out_bypass_mask_w[32];
  assign _0880_ = dat_out_bypass_p0_vld_w & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17253" *) dat_out_bypass_mask_w[33];
  assign _0881_ = dat_out_bypass_p0_vld_w & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17263" *) dat_out_bypass_mask_w[34];
  assign _0882_ = dat_out_bypass_p0_vld_w & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17273" *) dat_out_bypass_mask_w[35];
  assign _0883_ = dat_out_bypass_p0_vld_w & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17283" *) dat_out_bypass_mask_w[36];
  assign _0884_ = dat_out_bypass_p0_vld_w & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17293" *) dat_out_bypass_mask_w[37];
  assign _0885_ = dat_out_bypass_p0_vld_w & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17303" *) dat_out_bypass_mask_w[38];
  assign _0886_ = dat_out_bypass_p0_vld_w & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17313" *) dat_out_bypass_mask_w[39];
  assign _0887_ = dat_out_bypass_p0_vld_w & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17323" *) dat_out_bypass_mask_w[40];
  assign _0888_ = dat_out_bypass_p0_vld_w & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17333" *) dat_out_bypass_mask_w[41];
  assign _0889_ = dat_out_bypass_p0_vld_w & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17343" *) dat_out_bypass_mask_w[42];
  assign _0890_ = dat_out_bypass_p0_vld_w & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17353" *) dat_out_bypass_mask_w[43];
  assign _0891_ = dat_out_bypass_p0_vld_w & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17363" *) dat_out_bypass_mask_w[44];
  assign _0892_ = dat_out_bypass_p0_vld_w & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17373" *) dat_out_bypass_mask_w[45];
  assign _0893_ = dat_out_bypass_p0_vld_w & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17383" *) dat_out_bypass_mask_w[46];
  assign _0894_ = dat_out_bypass_p0_vld_w & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17393" *) dat_out_bypass_mask_w[47];
  assign _0895_ = dat_out_bypass_p0_vld_w & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17403" *) dat_out_bypass_mask_w[48];
  assign _0896_ = dat_out_bypass_p0_vld_w & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17413" *) dat_out_bypass_mask_w[49];
  assign _0897_ = dat_out_bypass_p0_vld_w & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17423" *) dat_out_bypass_mask_w[50];
  assign _0898_ = dat_out_bypass_p0_vld_w & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17433" *) dat_out_bypass_mask_w[51];
  assign _0899_ = dat_out_bypass_p0_vld_w & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17443" *) dat_out_bypass_mask_w[52];
  assign _0900_ = dat_out_bypass_p0_vld_w & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17453" *) dat_out_bypass_mask_w[53];
  assign _0901_ = dat_out_bypass_p0_vld_w & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17463" *) dat_out_bypass_mask_w[54];
  assign _0902_ = dat_out_bypass_p0_vld_w & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17473" *) dat_out_bypass_mask_w[55];
  assign _0903_ = dat_out_bypass_p0_vld_w & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17483" *) dat_out_bypass_mask_w[56];
  assign _0904_ = dat_out_bypass_p0_vld_w & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17493" *) dat_out_bypass_mask_w[57];
  assign _0905_ = dat_out_bypass_p0_vld_w & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17503" *) dat_out_bypass_mask_w[58];
  assign _0906_ = dat_out_bypass_p0_vld_w & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17513" *) dat_out_bypass_mask_w[59];
  assign _0907_ = dat_out_bypass_p0_vld_w & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17523" *) dat_out_bypass_mask_w[60];
  assign _0908_ = dat_out_bypass_p0_vld_w & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17533" *) dat_out_bypass_mask_w[61];
  assign _0909_ = dat_out_bypass_p0_vld_w & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17543" *) dat_out_bypass_mask_w[62];
  assign _0910_ = dat_out_bypass_p0_vld_w & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17553" *) dat_out_bypass_mask_w[63];
  assign _0911_ = dat_out_bypass_p1_vld_w & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17563" *) dat_out_bypass_mask_w[64];
  assign _0912_ = dat_out_bypass_p1_vld_w & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17573" *) dat_out_bypass_mask_w[65];
  assign _0913_ = dat_out_bypass_p1_vld_w & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17583" *) dat_out_bypass_mask_w[66];
  assign _0914_ = dat_out_bypass_p1_vld_w & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17593" *) dat_out_bypass_mask_w[67];
  assign _0915_ = dat_out_bypass_p1_vld_w & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17603" *) dat_out_bypass_mask_w[68];
  assign _0916_ = dat_out_bypass_p1_vld_w & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17613" *) dat_out_bypass_mask_w[69];
  assign _0917_ = dat_out_bypass_p1_vld_w & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17623" *) dat_out_bypass_mask_w[70];
  assign _0918_ = dat_out_bypass_p1_vld_w & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17633" *) dat_out_bypass_mask_w[71];
  assign _0919_ = dat_out_bypass_p1_vld_w & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17643" *) dat_out_bypass_mask_w[72];
  assign _0920_ = dat_out_bypass_p1_vld_w & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17653" *) dat_out_bypass_mask_w[73];
  assign _0921_ = dat_out_bypass_p1_vld_w & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17663" *) dat_out_bypass_mask_w[74];
  assign _0922_ = dat_out_bypass_p1_vld_w & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17673" *) dat_out_bypass_mask_w[75];
  assign _0923_ = dat_out_bypass_p1_vld_w & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17683" *) dat_out_bypass_mask_w[76];
  assign _0924_ = dat_out_bypass_p1_vld_w & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17693" *) dat_out_bypass_mask_w[77];
  assign _0925_ = dat_out_bypass_p1_vld_w & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17703" *) dat_out_bypass_mask_w[78];
  assign _0926_ = dat_out_bypass_p1_vld_w & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17713" *) dat_out_bypass_mask_w[79];
  assign _0927_ = dat_out_bypass_p1_vld_w & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17723" *) dat_out_bypass_mask_w[80];
  assign _0928_ = dat_out_bypass_p1_vld_w & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17733" *) dat_out_bypass_mask_w[81];
  assign _0929_ = dat_out_bypass_p1_vld_w & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17743" *) dat_out_bypass_mask_w[82];
  assign _0930_ = dat_out_bypass_p1_vld_w & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17753" *) dat_out_bypass_mask_w[83];
  assign _0931_ = dat_out_bypass_p1_vld_w & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17763" *) dat_out_bypass_mask_w[84];
  assign _0932_ = dat_out_bypass_p1_vld_w & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17773" *) dat_out_bypass_mask_w[85];
  assign _0933_ = dat_out_bypass_p1_vld_w & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17783" *) dat_out_bypass_mask_w[86];
  assign _0934_ = dat_out_bypass_p1_vld_w & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17793" *) dat_out_bypass_mask_w[87];
  assign _0935_ = dat_out_bypass_p1_vld_w & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17803" *) dat_out_bypass_mask_w[88];
  assign _0936_ = dat_out_bypass_p1_vld_w & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17813" *) dat_out_bypass_mask_w[89];
  assign _0937_ = dat_out_bypass_p1_vld_w & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17823" *) dat_out_bypass_mask_w[90];
  assign _0938_ = dat_out_bypass_p1_vld_w & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17833" *) dat_out_bypass_mask_w[91];
  assign _0939_ = dat_out_bypass_p1_vld_w & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17843" *) dat_out_bypass_mask_w[92];
  assign _0940_ = dat_out_bypass_p1_vld_w & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17853" *) dat_out_bypass_mask_w[93];
  assign _0941_ = dat_out_bypass_p1_vld_w & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17863" *) dat_out_bypass_mask_w[94];
  assign _0942_ = dat_out_bypass_p1_vld_w & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17873" *) dat_out_bypass_mask_w[95];
  assign _0943_ = dat_out_bypass_p1_vld_w & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17883" *) dat_out_bypass_mask_w[96];
  assign _0944_ = dat_out_bypass_p1_vld_w & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17893" *) dat_out_bypass_mask_w[97];
  assign _0945_ = dat_out_bypass_p1_vld_w & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17903" *) dat_out_bypass_mask_w[98];
  assign _0946_ = dat_out_bypass_p1_vld_w & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17913" *) dat_out_bypass_mask_w[99];
  assign _0947_ = dat_out_bypass_p1_vld_w & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17923" *) dat_out_bypass_mask_w[100];
  assign _0948_ = dat_out_bypass_p1_vld_w & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17933" *) dat_out_bypass_mask_w[101];
  assign _0949_ = dat_out_bypass_p1_vld_w & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17943" *) dat_out_bypass_mask_w[102];
  assign _0950_ = dat_out_bypass_p1_vld_w & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17953" *) dat_out_bypass_mask_w[103];
  assign _0951_ = dat_out_bypass_p1_vld_w & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17963" *) dat_out_bypass_mask_w[104];
  assign _0952_ = dat_out_bypass_p1_vld_w & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17973" *) dat_out_bypass_mask_w[105];
  assign _0953_ = dat_out_bypass_p1_vld_w & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17983" *) dat_out_bypass_mask_w[106];
  assign _0954_ = dat_out_bypass_p1_vld_w & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17993" *) dat_out_bypass_mask_w[107];
  assign _0955_ = dat_out_bypass_p1_vld_w & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18003" *) dat_out_bypass_mask_w[108];
  assign _0956_ = dat_out_bypass_p1_vld_w & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18013" *) dat_out_bypass_mask_w[109];
  assign _0957_ = dat_out_bypass_p1_vld_w & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18023" *) dat_out_bypass_mask_w[110];
  assign _0958_ = dat_out_bypass_p1_vld_w & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18033" *) dat_out_bypass_mask_w[111];
  assign _0959_ = dat_out_bypass_p1_vld_w & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18043" *) dat_out_bypass_mask_w[112];
  assign _0960_ = dat_out_bypass_p1_vld_w & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18053" *) dat_out_bypass_mask_w[113];
  assign _0961_ = dat_out_bypass_p1_vld_w & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18063" *) dat_out_bypass_mask_w[114];
  assign _0962_ = dat_out_bypass_p1_vld_w & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18073" *) dat_out_bypass_mask_w[115];
  assign _0963_ = dat_out_bypass_p1_vld_w & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18083" *) dat_out_bypass_mask_w[116];
  assign _0964_ = dat_out_bypass_p1_vld_w & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18093" *) dat_out_bypass_mask_w[117];
  assign _0965_ = dat_out_bypass_p1_vld_w & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18103" *) dat_out_bypass_mask_w[118];
  assign _0966_ = dat_out_bypass_p1_vld_w & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18113" *) dat_out_bypass_mask_w[119];
  assign _0967_ = dat_out_bypass_p1_vld_w & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18123" *) dat_out_bypass_mask_w[120];
  assign _0968_ = dat_out_bypass_p1_vld_w & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18133" *) dat_out_bypass_mask_w[121];
  assign _0969_ = dat_out_bypass_p1_vld_w & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18143" *) dat_out_bypass_mask_w[122];
  assign _0970_ = dat_out_bypass_p1_vld_w & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18153" *) dat_out_bypass_mask_w[123];
  assign _0971_ = dat_out_bypass_p1_vld_w & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18163" *) dat_out_bypass_mask_w[124];
  assign _0972_ = dat_out_bypass_p1_vld_w & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18173" *) dat_out_bypass_mask_w[125];
  assign _0973_ = dat_out_bypass_p1_vld_w & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18183" *) dat_out_bypass_mask_w[126];
  assign _0974_ = dat_out_bypass_p1_vld_w & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18193" *) dat_out_bypass_mask_w[127];
  assign dat_rsp_pra_en = dat_rsp_pvld & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18209" *) is_winograd_d1[19];
  assign layer_st = reg2dp_op_en & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1906" *) is_sg_idle;
  assign is_img = is_conv & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1927" *) reg2dp_datain_format;
  assign slcg_wg_en_w = reg2dp_op_en & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:6613" *) reg2dp_conv_mode;
  assign sub_rls = dat_rsp_pvld & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:7433" *) dat_rsp_pd[17];
  assign _0975_ = sg2dl_reuse_rls & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:7446" *) _1160_;
  assign _0976_ = sub_rls & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:7446" *) _1161_;
  assign _0977_ = sub_h_total_g0[2] & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:8505" *) dl_pvld_d1;
  assign _0978_ = sub_h_total_g0[1] & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:8506" *) dl_pvld_d3;
  assign _0979_ = sub_h_total_g0[0] & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:8507" *) dl_pvld_d4;
  assign { _1018_[30:13], _0980_ } = { sub_h_total_g1[2], sub_h_total_g1[2], sub_h_total_g1[2], sub_h_total_g1[2], sub_h_total_g1[2], sub_h_total_g1[2], sub_h_total_g1[2], sub_h_total_g1[2], sub_h_total_g1[2], sub_h_total_g1[2], sub_h_total_g1[2], sub_h_total_g1[2], sub_h_total_g1[2], sub_h_total_g1[2], sub_h_total_g1[2], sub_h_total_g1[2], sub_h_total_g1[2], sub_h_total_g1[2], sub_h_total_g1[2], sub_h_total_g1[2], sub_h_total_g1[2], sub_h_total_g1[2], sub_h_total_g1[2], sub_h_total_g1[2], sub_h_total_g1[2], sub_h_total_g1[2], sub_h_total_g1[2], sub_h_total_g1[2], sub_h_total_g1[2], sub_h_total_g1[2], sub_h_total_g1[2] } & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:8515" *) dl_pd_d1;
  assign _0981_ = { sub_h_total_g1[1], sub_h_total_g1[1], sub_h_total_g1[1], sub_h_total_g1[1], sub_h_total_g1[1], sub_h_total_g1[1], sub_h_total_g1[1], sub_h_total_g1[1], sub_h_total_g1[1], sub_h_total_g1[1], sub_h_total_g1[1], sub_h_total_g1[1], sub_h_total_g1[1], sub_h_total_g1[1], sub_h_total_g1[1], sub_h_total_g1[1], sub_h_total_g1[1], sub_h_total_g1[1], sub_h_total_g1[1], sub_h_total_g1[1], sub_h_total_g1[1], sub_h_total_g1[1], sub_h_total_g1[1], sub_h_total_g1[1], sub_h_total_g1[1], sub_h_total_g1[1], sub_h_total_g1[1], sub_h_total_g1[1], sub_h_total_g1[1], sub_h_total_g1[1], sub_h_total_g1[1] } & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:8516" *) dl_pd_d3;
  assign _0982_ = { sub_h_total_g1[0], sub_h_total_g1[0], sub_h_total_g1[0], sub_h_total_g1[0], sub_h_total_g1[0], sub_h_total_g1[0], sub_h_total_g1[0], sub_h_total_g1[0], sub_h_total_g1[0], sub_h_total_g1[0], sub_h_total_g1[0], sub_h_total_g1[0], sub_h_total_g1[0], sub_h_total_g1[0], sub_h_total_g1[0], sub_h_total_g1[0], sub_h_total_g1[0], sub_h_total_g1[0], sub_h_total_g1[0], sub_h_total_g1[0], sub_h_total_g1[0], sub_h_total_g1[0], sub_h_total_g1[0], sub_h_total_g1[0], sub_h_total_g1[0], sub_h_total_g1[0], sub_h_total_g1[0], sub_h_total_g1[0], sub_h_total_g1[0], sub_h_total_g1[0], sub_h_total_g1[0] } & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:8517" *) dl_pd_d4;
  assign _0983_ = _1154_ & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:8728" *) dat_exec_valid;
  assign _0984_ = is_stripe_equal & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:8807" *) _1112_;
  assign is_stripe_equal = is_batch_end & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:8816" *) _1062_;
  assign is_stripe_end = is_stripe_equal & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:8822" *) is_sub_h_end;
  assign _0985_ = dat_exec_valid & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:8829" *) is_batch_end;
  assign _0986_ = _1113_ & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:9100" *) _1114_;
  assign _0987_ = _0986_ & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:9100" *) _1115_;
  assign _0988_ = is_batch_end & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:9348" *) is_sub_h_end;
  assign is_w_end = _0988_ & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:9348" *) _1066_;
  assign is_w_end_ahead = is_batch_end & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:9355" *) _1066_;
  assign _0989_ = _0985_ & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:9377" *) is_sub_h_end;
  assign _0990_ = is_stripe_end & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:9655" *) dl_pd[26];
  assign _0991_ = _0990_ & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:9655" *) dl_pd[27];
  assign _0992_ = _0991_ & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:9655" *) is_w_end;
  assign _0993_ = _0991_ & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:9656" *) _1116_;
  assign _0994_ = _0990_ & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:9657" *) _1078_;
  assign _0995_ = is_stripe_end & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:9658" *) _1117_;
  assign _0996_ = _0989_ & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:9669" *) _1118_;
  assign _0997_ = dat_exec_valid & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:9678" *) _1119_;
  assign _0998_ = _0997_ & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:9678" *) is_stripe_end;
  assign _0999_ = _0998_ & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:9678" *) dl_pd[27];
  assign _1000_ = dat_exec_valid & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:9687" *) is_img_d1[2];
  assign _1001_ = _1000_ & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:9687" *) _1155_;
  assign _1002_ = dat_exec_valid & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:9696" *) is_img_d1[3];
  assign _1003_ = _1002_ & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:9696" *) is_stripe_end;
  assign _1004_ = _1003_ & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:9696" *) dl_pd[26];
  assign _1005_ = dat_exec_valid & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:9706" *) is_img_d1[4];
  assign _1006_ = _1005_ & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:9706" *) is_stripe_end;
  assign _1007_ = _1006_ & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:9706" *) dl_pd[26];
  assign _1008_ = _1007_ & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:9706" *) dl_pd[27];
  assign _1009_ = dl_pd[27] & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:9732" *) is_w_end_ahead;
  assign _1010_ = is_int8_d1[1] & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:9733" *) dl_pd[27];
  assign _1011_ = _1010_ & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:9733" *) _1116_;
  assign _1012_ = _1011_ & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:9733" *) pixel_x_stride_odd;
  assign _1013_ = _1011_ & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:9734" *) _1121_;
  assign _1014_ = is_int8_d1[1] & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:9735" *) _1078_;
  assign _1015_ = is_img_d1[0] & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:9740" *) dat_req_stripe_st;
  assign _1016_ = is_img_d1[0] & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:9743" *) is_sub_h_end;
  assign pixel_force_clr = _1016_ & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:9743" *) _1156_;
  assign _1026_ = ! (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:10474" *) sub_h_cnt;
  assign _1027_ = ! (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:12190" *) dat_req_sub_h_d1;
  assign _1028_ = dat_req_sub_h_d1 == (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:12191" *) 1'b1;
  assign _1029_ = dat_req_sub_h_d1 == (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:12192" *) 2'b10;
  assign _1030_ = dat_req_sub_h_d1 == (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:12197" *) 2'b11;
  assign _1032_ = ! (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:14531" *) dat_rsp_exec_sub_h_d6;
  assign _1033_ = dat_rsp_exec_sub_h_d6 == (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:14532" *) 1'b1;
  assign _1034_ = dat_rsp_exec_sub_h_d6 == (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:14535" *) 2'b10;
  assign _1035_ = dat_rsp_exec_sub_h_d6 == (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:14537" *) 2'b11;
  assign _1036_ = sub_h_total_g5 == (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15241" *) 3'b100;
  assign _1037_ = sub_h_total_g6 == (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15263" *) 3'b100;
  assign _1038_ = ~ (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15961" *) dat_rsp_pd[0];
  assign _1039_ = ! (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15963" *) dat_rsp_pd[1:0];
  assign _1040_ = dat_rsp_pd[1:0] == (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15964" *) 1'b1;
  assign _1041_ = dat_rsp_pd[1:0] == (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15965" *) 2'b10;
  assign _1042_ = dat_rsp_pd[1:0] == (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15966" *) 2'b11;
  assign rsp_sft_l1_sel_3 = rsp_sft_cnt_l1[7:6] == (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15999" *) 2'b11;
  assign rsp_sft_l1_sel_2 = rsp_sft_cnt_l1[7:6] == (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16000" *) 2'b10;
  assign rsp_sft_l1_sel_1 = rsp_sft_cnt_l1[7:6] == (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16001" *) 1'b1;
  assign rsp_sft_l2_sel_3 = rsp_sft_cnt_l2[7:6] == (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16006" *) 2'b11;
  assign rsp_sft_l2_sel_2 = rsp_sft_cnt_l2[7:6] == (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16007" *) 2'b10;
  assign rsp_sft_l2_sel_1 = rsp_sft_cnt_l2[7:6] == (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16008" *) 1'b1;
  assign rsp_sft_l3_sel_3 = rsp_sft_cnt_l3[7:6] == (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16013" *) 2'b11;
  assign rsp_sft_l3_sel_2 = rsp_sft_cnt_l3[7:6] == (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16014" *) 2'b10;
  assign rsp_sft_l3_sel_1 = rsp_sft_cnt_l3[7:6] == (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16015" *) 1'b1;
  assign _1043_ = sub_h_total_g7 == (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16105" *) 3'b100;
  assign _1044_ = sub_h_total_g7 == (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16106" *) 2'b10;
  assign _1045_ = sub_h_total_g8 == (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16122" *) 3'b100;
  assign _1046_ = sub_h_total_g8 == (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16123" *) 2'b10;
  assign _1047_ = sub_h_total_g9 == (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16142" *) 3'b100;
  assign _1048_ = dat_rsp_pd[16:15] == (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16278" *) 2'b11;
  assign _1049_ = sub_h_total_g10 == (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16302" *) 3'b100;
  assign _1050_ = sub_h_total_g10 == (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16303" *) 2'b10;
  assign _1051_ = sub_h_total_g11 == (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16312" *) 3'b100;
  assign _1052_ = sub_h_total_g11 == (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16313" *) 2'b10;
  assign is_sg_idle = ! (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1880" *) sc_state;
  assign is_sg_done = sc_state == (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1890" *) 2'b11;
  assign is_conv = ~ (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1921" *) reg2dp_conv_mode;
  assign is_int8 = ! (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1953" *) reg2dp_proc_precision;
  assign is_fp16 = reg2dp_proc_precision == (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1958" *) 2'b10;
  assign _1055_ = reg2dp_datain_channel_ext[1:0] == (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:2017" *) 2'b11;
  assign _1056_ = reg2dp_datain_channel_ext[1:0] == (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:2018" *) 2'b10;
  assign _1057_ = reg2dp_y_extension == (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:2027" *) 2'b10;
  assign _1058_ = reg2dp_y_extension == (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:2028" *) 1'b1;
  assign _1059_ = reg2dp_pra_truncate == (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:2159" *) 2'b11;
  assign is_batch_end = batch_cnt == (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:8545" *) batch_cmp;
  assign is_sub_h_end = sub_h_cnt_inc == (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:8720" *) sub_h_cmp_g0;
  assign _1062_ = stripe_cnt_inc == (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:8816" *) dl_pd[23:17];
  assign is_last_channel = datain_c_cnt == (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:9520" *) datain_channel_cmp;
  assign is_dat_req_addr_wrap = dat_req_addr_sum >= (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:12163" *) { data_bank, 8'b00000000 };
  assign _1063_ = dat_rsp_pd[16:15] >= (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16276" *) 1'b1;
  assign _1064_ = dat_rsp_pd[16:15] >= (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16277" *) 2'b10;
  assign _1065_ = reg2dp_weight_channel_ext >= (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:2029" *) 6'b111111;
  assign is_dat_entry_st_wrap = dat_entry_st_inc >= (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:6715" *) { data_bank, 8'b00000000 };
  assign _1066_ = dataout_w_cnt >= (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:9348" *) dataout_width_cmp;
  assign _1067_ = datain_w_cur > (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:10409" *) datain_width_cmp;
  assign _1068_ = datain_h_cur > (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:10410" *) datain_height_cmp;
  assign dat_img_req_skip = w_bias_w[13:2] > (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:10429" *) entries_cmp;
  assign _1069_ = dat_req_bytes > (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:11406" *) 6'b100000;
  assign _1070_ = dat_req_bytes > (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:11419" *) 7'b1000000;
  assign _1071_ = dat_rsp_pd[14:7] > (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15961" *) 6'b100000;
  assign _1072_ = dat_rsp_pd[14:7] <= (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15961" *) 7'b1000000;
  assign _1073_ = dat_rsp_pd[14:7] <= (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15963" *) 6'b100000;
  assign dl_h_offset_ext = dl_pd[9:5] * (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:10270" *) y_dilate;
  assign h_bias_0_w = datain_h_cnt[11:0] * (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:11365" *) h_bias_0_stride;
  assign h_bias_1_w = dl_pd[9:5] * (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:11372" *) h_bias_1_stride;
  assign h_bias_2_w = batch_cnt * (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:11379" *) h_bias_2_stride;
  assign _1019_[11:0] = sub_h_cnt * (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:11388" *) h_bias_3_stride;
  assign entries_batch_w = entries_single_w * (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:2090" *) data_batch_w;
  assign h_offset_slice_w = data_batch_w * (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:2105" *) y_dilate_w;
  assign h_bias_0_stride_w = entries * (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:2112" *) data_batch;
  assign h_bias_1_stride_w = entries * (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:2119" *) h_offset_slice;
  assign slice_entries_w = entries_batch * (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:2149" *) slices_oprand;
  assign dl_w_offset_ext = dl_pd[4:0] * (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:9712" *) x_dilate;
  assign c_bias_d1_reg_en = c_bias != (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:11357" *) c_bias_d1;
  assign _1074_ = dat_req_addr_last != (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:12188" *) dat_req_addr_w;
  assign _1075_ = sub_h_total_g5 != (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15240" *) 1'b1;
  assign _1076_ = sub_h_total_g6 != (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15262" *) 1'b1;
  assign _1077_ = sub_h_total_g9 != (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16140" *) 1'b1;
  assign _1078_ = ~ (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:10245" *) dl_pd[27];
  assign _1079_ = ~ (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:10455" *) dat_req_dummy;
  assign _1080_ = ~ (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:10455" *) dat_req_skip;
  assign _1081_ = ~ (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:10471" *) datain_w_cur[1];
  assign _1082_ = ~ (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:11330" *) is_img_d1[8];
  assign _1083_ = ~ (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:11330" *) is_int8_d1[3];
  assign _1084_ = ~ (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:11405" *) is_last_channel;
  assign _1085_ = ~ (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:14533" *) is_winograd_d1[10];
  assign _1086_ = ~ (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:14552" *) dat_rsp_exec_sub_h_d6[0];
  assign _1087_ = ~ (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:14553" *) dat_l0c0_dummy;
  assign _1088_ = ~ (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:14555" *) dat_l1c0_dummy;
  assign _1089_ = ~ (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:14557" *) dat_l2c0_dummy;
  assign _1090_ = ~ (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:14558" *) dat_l3c0_dummy;
  assign _1091_ = ~ (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:14564" *) dat_rsp_pipe_pd_d6[18];
  assign _1092_ = ~ (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15176" *) dat_rsp_pd_d1[4];
  assign _1093_ = ~ (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15178" *) dat_rsp_pd_d1[6];
  assign _1094_ = ~ (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15192" *) dat_rsp_pd_d2[4];
  assign _1095_ = ~ (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15194" *) dat_rsp_pd_d2[6];
  assign _1096_ = ~ (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15208" *) dat_rsp_pd_d3[4];
  assign _1097_ = ~ (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15210" *) dat_rsp_pd_d3[6];
  assign _1098_ = ~ (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15224" *) dat_rsp_pd_d4[4];
  assign _1099_ = ~ (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15226" *) dat_rsp_pd_d4[6];
  assign _1100_ = ~ (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15780" *) dat_rsp_pd[2];
  assign dat_rsp_wg_sel_16b = ~ (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15789" *) is_int8_d1[5];
  assign _1101_ = ~ (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15790" *) dat_rsp_pd[4];
  assign _1102_ = ~ (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15980" *) is_int8_d1[10];
  assign _1103_ = ~ (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16104" *) is_img_d1[31];
  assign _1104_ = ~ (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16121" *) is_img_d1[32];
  assign _1105_ = ~ (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16121" *) is_int8_d1[12];
  assign _1106_ = ~ (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16141" *) is_int8_d1[14];
  assign _1107_ = ~ (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16143" *) is_int8_d1[15];
  assign _1108_ = ~ (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16145" *) is_int8_d1[16];
  assign dat_rsp_ori_mask = ~ (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16271" *) _1166_;
  assign _1109_ = ~ (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16378" *) is_int8_d1[18];
  assign _1110_ = ~ (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16378" *) is_winograd_d1[15];
  assign _1111_ = ~ (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16379" *) is_winograd_d1[16];
  assign _1112_ = ~ (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:8807" *) is_sub_h_end;
  assign _1113_ = ~ (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:9100" *) _1163_;
  assign _1114_ = ~ (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:9100" *) _1164_;
  assign _1115_ = ~ (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:9100" *) _1165_;
  assign _1116_ = ~ (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:9656" *) is_w_end;
  assign _1117_ = ~ (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:9658" *) dl_pd[26];
  assign _1118_ = ~ (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:9669" *) is_img_d1[0];
  assign _1119_ = ~ (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:9678" *) is_img_d1[1];
  assign _1120_ = ~ (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:9733" *) pixel_req_ch_odd_ori;
  assign _1121_ = ~ (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:9734" *) pixel_x_stride_odd;
  assign _1122_ = ~ (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:9735" *) pixel_req_ch_odd;
  assign _1123_ = layer_st | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:10244" *) _0732_;
  assign _1124_ = _0733_ | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:10256" *) is_w_end;
  assign datain_h_cnt_reg_en = layer_st | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:10256" *) _0734_;
  assign datain_h_ori_reg_en = layer_st | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:10264" *) _0736_;
  assign _1125_ = datain_w_cur[13] | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:10410" *) _1067_;
  assign _1126_ = _1125_ | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:10410" *) datain_h_cur[13];
  assign dat_conv_req_dummy = _1126_ | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:10410" *) _1068_;
  assign dat_img_req_dummy = datain_h_cur[13] | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:10423" *) _1068_;
  assign dat_req_skip = _0738_ | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:10448" *) _0739_;
  assign _1127_ = _1083_ | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:11330" *) datain_c_cnt[0];
  assign c_bias_reg_en = layer_st | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:11351" *) _0746_;
  assign _1128_ = is_winograd_d1[7] | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:11391" *) is_img_d1[9];
  assign h_bias_reg_en[1] = layer_st | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:11391" *) _0747_;
  assign _1129_ = _1084_ | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:11405" *) datain_c_cnt[0];
  assign _1130_ = _1129_ | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:11405" *) is_winograd_d1[8];
  assign _1131_ = _1070_ | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:11419" *) is_winograd_d1[9];
  assign _1132_ = layer_st | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:12179" *) dat_req_dummy_d1;
  assign _1133_ = _1074_ | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:12188" *) pixel_force_fetch_d1;
  assign _1134_ = dat_req_valid_d1 | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:12194" *) dat_req_dummy_d1;
  assign dat_req_sub_h_0_addr_en = layer_st | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:12194" *) _0748_;
  assign dat_req_sub_h_1_addr_en = layer_st | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:12195" *) _0749_;
  assign dat_req_sub_h_2_addr_en = layer_st | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:12196" *) _0750_;
  assign dat_req_sub_h_3_addr_en = layer_st | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:12197" *) _0751_;
  assign _1031_ = layer_st | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:12453" *) sc2buf_dat_rd_en_w;
  assign dat_l0c1_en = _0752_ | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:14553" *) _0754_;
  assign dat_l1c1_en = _0755_ | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:14555" *) _0757_;
  assign dat_l0_set = dat_l0c0_en | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:14589" *) dat_dummy_l0_en;
  assign dat_l1_set = dat_l1c0_en | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:14590" *) dat_dummy_l1_en;
  assign dat_l2_set = dat_l2c0_en | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:14591" *) dat_dummy_l2_en;
  assign dat_l3_set = dat_l3c0_en | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:14592" *) dat_dummy_l3_en;
  assign _1135_ = _0766_ | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15042" *) _0767_;
  assign dat_rsp_pvld = _1135_ | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15043" *) _0768_;
  assign _1136_ = { _1017_[26:12], _0769_ } | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15063" *) _0770_;
  assign dat_rsp_pd = _1136_ | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15064" *) _0771_;
  assign rsp_sft_cnt_l0_en = layer_st | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15239" *) _0792_;
  assign rsp_sft_cnt_l1_en = layer_st | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15240" *) _0794_;
  assign rsp_sft_cnt_l2_en = layer_st | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15241" *) _0796_;
  assign rsp_sft_cnt_l3_en = layer_st | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15242" *) _0798_;
  assign rsp_sft_cnt_l0_ori_en = layer_st | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15261" *) _0801_;
  assign rsp_sft_cnt_l1_ori_en = layer_st | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15262" *) _0805_;
  assign rsp_sft_cnt_l2_ori_en = layer_st | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15263" *) _0809_;
  assign rsp_sft_cnt_l3_ori_en = layer_st | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15264" *) _0813_;
  assign _1137_ = _0814_ | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15812" *) _0815_;
  assign _1138_ = _1137_ | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15813" *) _0816_;
  assign dat_rsp_wg = _1138_ | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15814" *) _0817_;
  assign _1139_ = _0818_ | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15857" *) _0819_;
  assign dat_rsp_wg_ch0 = _1139_ | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15858" *) _0820_;
  assign _1140_ = _0821_ | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15869" *) _0822_;
  assign dat_rsp_wg_ch1 = _1140_ | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15870" *) _0823_;
  assign _1141_ = _0824_ | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15881" *) _0825_;
  assign dat_rsp_wg_ch2 = _1141_ | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15882" *) _0826_;
  assign _1142_ = _0827_ | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15893" *) _0828_;
  assign dat_rsp_wg_ch3 = _1142_ | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15894" *) _0829_;
  assign _1143_ = is_int8_d1[9] | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15960" *) is_winograd_d1[13];
  assign _1144_ = _1143_ | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15960" *) is_img_d1[25];
  assign _1145_ = _1102_ | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15980" *) is_winograd_d1[14];
  assign _1146_ = _1145_ | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15980" *) is_img_d1[26];
  assign _1147_ = dat_rsp_pd[4] | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15986" *) _0838_;
  assign dat_rsp_conv = dat_rsp_conv_16b | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15993" *) { dat_rsp_conv_8b, dat_rsp_conv_8b };
  assign _1148_ = _1103_ | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16104" *) is_int8_d1[11];
  assign _1149_ = _1104_ | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16121" *) _1105_;
  assign _1053_ = dat_out_pvld | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18509" *) dl_out_pvld;
  assign _1150_ = reg2dp_conv_mode | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1940" *) is_img;
  assign _1054_ = dl_out_pvld | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:19941" *) sc2mac_dat_b_pvld;
  assign _1060_ = sc2cdma_dat_pending_req | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:6884" *) dat_rls;
  assign dat_rls = _0975_ | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:7446" *) _0976_;
  assign _1151_ = _0977_ | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:8506" *) _0978_;
  assign dat_req_stripe_st = _1151_ | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:8507" *) _0979_;
  assign _1152_ = { _1018_[30:13], _0980_ } | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:8516" *) _0981_;
  assign dl_pd = _1152_ | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:8517" *) _0982_;
  assign _1061_ = layer_st | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:8551" *) dat_exec_valid;
  assign _1153_ = layer_st | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:8713" *) is_sub_h_end;
  assign _1154_ = is_winograd_d1[2] | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:8728" *) _1162_;
  assign sub_h_cnt_reg_en = layer_st | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:8728" *) _0983_;
  assign stripe_cnt_reg_en = layer_st | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:8829" *) _0985_;
  assign dat_pipe_valid = dat_req_stripe_st | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:9091" *) dat_pipe_local_valid;
  assign dataout_w_cnt_reg_en = layer_st | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:9377" *) _0989_;
  assign datain_w_cnt_reg_en = layer_st | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:9669" *) _0996_;
  assign datain_w_ori_reg_en = layer_st | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:9678" *) _0999_;
  assign _1155_ = is_sub_h_end | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:9687" *) is_w_end;
  assign pixel_w_cnt_reg_en = layer_st_d1 | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:9687" *) _1001_;
  assign pixel_req_ch_odd_en = layer_st_d1 | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:9696" *) _1004_;
  assign pixel_ch_ori_reg_en = layer_st_d1 | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:9706" *) _1008_;
  assign _1156_ = pixel_force_fetch | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:9743" *) pixel_force_fetch_d1;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_b_data127 <= _0583_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_b_data126 <= _0582_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_b_data125 <= _0581_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_b_data124 <= _0580_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_b_data123 <= _0579_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_b_data122 <= _0578_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_b_data121 <= _0577_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_b_data120 <= _0576_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_b_data119 <= _0574_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_b_data118 <= _0573_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_b_data117 <= _0572_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_b_data116 <= _0571_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_b_data115 <= _0570_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_b_data114 <= _0569_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_b_data113 <= _0568_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_b_data112 <= _0567_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_b_data111 <= _0566_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_b_data110 <= _0565_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_b_data109 <= _0563_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_b_data108 <= _0562_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_b_data107 <= _0561_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_b_data106 <= _0560_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_b_data105 <= _0559_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_b_data104 <= _0558_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_b_data103 <= _0557_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_b_data102 <= _0556_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_b_data101 <= _0555_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_b_data100 <= _0554_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_b_data99 <= _0679_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_b_data98 <= _0678_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_b_data97 <= _0677_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_b_data96 <= _0676_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_b_data95 <= _0675_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_b_data94 <= _0674_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_b_data93 <= _0673_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_b_data92 <= _0672_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_b_data91 <= _0671_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_b_data90 <= _0670_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_b_data89 <= _0668_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_b_data88 <= _0667_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_b_data87 <= _0666_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_b_data86 <= _0665_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_b_data85 <= _0664_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_b_data84 <= _0663_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_b_data83 <= _0662_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_b_data82 <= _0661_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_b_data81 <= _0660_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_b_data80 <= _0659_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_b_data79 <= _0657_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_b_data78 <= _0656_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_b_data77 <= _0655_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_b_data76 <= _0654_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_b_data75 <= _0653_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_b_data74 <= _0652_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_b_data73 <= _0651_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_b_data72 <= _0650_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_b_data71 <= _0649_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_b_data70 <= _0648_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_b_data69 <= _0646_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_b_data68 <= _0645_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_b_data67 <= _0644_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_b_data66 <= _0643_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_b_data65 <= _0642_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_b_data64 <= _0641_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_b_data63 <= _0640_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_b_data62 <= _0639_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_b_data61 <= _0638_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_b_data60 <= _0637_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_b_data59 <= _0635_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_b_data58 <= _0634_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_b_data57 <= _0633_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_b_data56 <= _0632_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_b_data55 <= _0631_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_b_data54 <= _0630_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_b_data53 <= _0629_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_b_data52 <= _0628_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_b_data51 <= _0627_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_b_data50 <= _0626_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_b_data49 <= _0624_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_b_data48 <= _0623_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_b_data47 <= _0622_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_b_data46 <= _0621_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_b_data45 <= _0620_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_b_data44 <= _0619_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_b_data43 <= _0618_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_b_data42 <= _0617_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_b_data41 <= _0616_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_b_data40 <= _0615_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_b_data39 <= _0613_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_b_data38 <= _0612_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_b_data37 <= _0611_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_b_data36 <= _0610_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_b_data35 <= _0609_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_b_data34 <= _0608_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_b_data33 <= _0607_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_b_data32 <= _0606_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_b_data31 <= _0605_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_b_data30 <= _0604_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_b_data29 <= _0602_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_b_data28 <= _0601_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_b_data27 <= _0600_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_b_data26 <= _0599_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_b_data25 <= _0598_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_b_data24 <= _0597_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_b_data23 <= _0596_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_b_data22 <= _0595_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_b_data21 <= _0594_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_b_data20 <= _0593_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_b_data19 <= _0591_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_b_data18 <= _0590_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_b_data17 <= _0589_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_b_data16 <= _0588_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_b_data15 <= _0587_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_b_data14 <= _0586_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_b_data13 <= _0585_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_b_data12 <= _0584_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_b_data11 <= _0575_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_b_data10 <= _0564_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_b_data9 <= _0680_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_b_data8 <= _0669_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_b_data7 <= _0658_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_b_data6 <= _0647_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_b_data5 <= _0636_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_b_data4 <= _0625_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_b_data3 <= _0614_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_b_data2 <= _0603_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_b_data1 <= _0592_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_b_data0 <= _0553_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_a_data127 <= _0453_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_a_data126 <= _0452_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_a_data125 <= _0451_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_a_data124 <= _0450_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_a_data123 <= _0449_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_a_data122 <= _0448_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_a_data121 <= _0447_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_a_data120 <= _0446_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_a_data119 <= _0444_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_a_data118 <= _0443_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_a_data117 <= _0442_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_a_data116 <= _0441_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_a_data115 <= _0440_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_a_data114 <= _0439_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_a_data113 <= _0438_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_a_data112 <= _0437_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_a_data111 <= _0436_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_a_data110 <= _0435_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_a_data109 <= _0433_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_a_data108 <= _0432_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_a_data107 <= _0431_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_a_data106 <= _0430_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_a_data105 <= _0429_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_a_data104 <= _0428_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_a_data103 <= _0427_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_a_data102 <= _0426_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_a_data101 <= _0425_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_a_data100 <= _0424_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_a_data99 <= _0549_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_a_data98 <= _0548_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_a_data97 <= _0547_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_a_data96 <= _0546_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_a_data95 <= _0545_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_a_data94 <= _0544_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_a_data93 <= _0543_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_a_data92 <= _0542_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_a_data91 <= _0541_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_a_data90 <= _0540_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_a_data89 <= _0538_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_a_data88 <= _0537_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_a_data87 <= _0536_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_a_data86 <= _0535_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_a_data85 <= _0534_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_a_data84 <= _0533_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_a_data83 <= _0532_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_a_data82 <= _0531_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_a_data81 <= _0530_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_a_data80 <= _0529_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_a_data79 <= _0527_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_a_data78 <= _0526_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_a_data77 <= _0525_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_a_data76 <= _0524_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_a_data75 <= _0523_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_a_data74 <= _0522_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_a_data73 <= _0521_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_a_data72 <= _0520_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_a_data71 <= _0519_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_a_data70 <= _0518_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_a_data69 <= _0516_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_a_data68 <= _0515_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_a_data67 <= _0514_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_a_data66 <= _0513_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_a_data65 <= _0512_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_a_data64 <= _0511_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_a_data63 <= _0510_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_a_data62 <= _0509_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_a_data61 <= _0508_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_a_data60 <= _0507_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_a_data59 <= _0505_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_a_data58 <= _0504_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_a_data57 <= _0503_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_a_data56 <= _0502_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_a_data55 <= _0501_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_a_data54 <= _0500_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_a_data53 <= _0499_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_a_data52 <= _0498_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_a_data51 <= _0497_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_a_data50 <= _0496_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_a_data49 <= _0494_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_a_data48 <= _0493_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_a_data47 <= _0492_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_a_data46 <= _0491_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_a_data45 <= _0490_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_a_data44 <= _0489_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_a_data43 <= _0488_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_a_data42 <= _0487_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_a_data41 <= _0486_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_a_data40 <= _0485_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_a_data39 <= _0483_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_a_data38 <= _0482_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_a_data37 <= _0481_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_a_data36 <= _0480_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_a_data35 <= _0479_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_a_data34 <= _0478_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_a_data33 <= _0477_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_a_data32 <= _0476_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_a_data31 <= _0475_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_a_data30 <= _0474_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_a_data29 <= _0472_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_a_data28 <= _0471_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_a_data27 <= _0470_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_a_data26 <= _0469_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_a_data25 <= _0468_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_a_data24 <= _0467_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_a_data23 <= _0466_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_a_data22 <= _0465_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_a_data21 <= _0464_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_a_data20 <= _0463_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_a_data19 <= _0461_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_a_data18 <= _0460_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_a_data17 <= _0459_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_a_data16 <= _0458_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_a_data15 <= _0457_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_a_data14 <= _0456_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_a_data13 <= _0455_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_a_data12 <= _0454_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_a_data11 <= _0445_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_a_data10 <= _0434_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_a_data9 <= _0550_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_a_data8 <= _0539_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_a_data7 <= _0528_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_a_data6 <= _0517_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_a_data5 <= _0506_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_a_data4 <= _0495_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_a_data3 <= _0484_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_a_data2 <= _0473_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_a_data1 <= _0462_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_a_data0 <= _0423_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      sc2mac_dat_b_mask <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    else
      sc2mac_dat_b_mask <= _0681_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      sc2mac_dat_a_mask <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    else
      sc2mac_dat_a_mask <= _0551_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      sc2mac_dat_b_pd <= 9'b000000000;
    else
      sc2mac_dat_b_pd <= _0682_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      sc2mac_dat_a_pd <= 9'b000000000;
    else
      sc2mac_dat_a_pd <= _0552_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      sc2mac_dat_b_pvld <= 1'b0;
    else
      sc2mac_dat_b_pvld <= dl_out_pvld;
  always @(posedge nvdla_core_clk)
      dl_out_data127 <= _0272_;
  always @(posedge nvdla_core_clk)
      dl_out_data126 <= _0271_;
  always @(posedge nvdla_core_clk)
      dl_out_data125 <= _0270_;
  always @(posedge nvdla_core_clk)
      dl_out_data124 <= _0269_;
  always @(posedge nvdla_core_clk)
      dl_out_data123 <= _0268_;
  always @(posedge nvdla_core_clk)
      dl_out_data122 <= _0267_;
  always @(posedge nvdla_core_clk)
      dl_out_data121 <= _0266_;
  always @(posedge nvdla_core_clk)
      dl_out_data120 <= _0265_;
  always @(posedge nvdla_core_clk)
      dl_out_data119 <= _0263_;
  always @(posedge nvdla_core_clk)
      dl_out_data118 <= _0262_;
  always @(posedge nvdla_core_clk)
      dl_out_data117 <= _0261_;
  always @(posedge nvdla_core_clk)
      dl_out_data116 <= _0260_;
  always @(posedge nvdla_core_clk)
      dl_out_data115 <= _0259_;
  always @(posedge nvdla_core_clk)
      dl_out_data114 <= _0258_;
  always @(posedge nvdla_core_clk)
      dl_out_data113 <= _0257_;
  always @(posedge nvdla_core_clk)
      dl_out_data112 <= _0256_;
  always @(posedge nvdla_core_clk)
      dl_out_data111 <= _0255_;
  always @(posedge nvdla_core_clk)
      dl_out_data110 <= _0254_;
  always @(posedge nvdla_core_clk)
      dl_out_data109 <= _0252_;
  always @(posedge nvdla_core_clk)
      dl_out_data108 <= _0251_;
  always @(posedge nvdla_core_clk)
      dl_out_data107 <= _0250_;
  always @(posedge nvdla_core_clk)
      dl_out_data106 <= _0249_;
  always @(posedge nvdla_core_clk)
      dl_out_data105 <= _0248_;
  always @(posedge nvdla_core_clk)
      dl_out_data104 <= _0247_;
  always @(posedge nvdla_core_clk)
      dl_out_data103 <= _0246_;
  always @(posedge nvdla_core_clk)
      dl_out_data102 <= _0245_;
  always @(posedge nvdla_core_clk)
      dl_out_data101 <= _0244_;
  always @(posedge nvdla_core_clk)
      dl_out_data100 <= _0243_;
  always @(posedge nvdla_core_clk)
      dl_out_data99 <= _0368_;
  always @(posedge nvdla_core_clk)
      dl_out_data98 <= _0367_;
  always @(posedge nvdla_core_clk)
      dl_out_data97 <= _0366_;
  always @(posedge nvdla_core_clk)
      dl_out_data96 <= _0365_;
  always @(posedge nvdla_core_clk)
      dl_out_data95 <= _0364_;
  always @(posedge nvdla_core_clk)
      dl_out_data94 <= _0363_;
  always @(posedge nvdla_core_clk)
      dl_out_data93 <= _0362_;
  always @(posedge nvdla_core_clk)
      dl_out_data92 <= _0361_;
  always @(posedge nvdla_core_clk)
      dl_out_data91 <= _0360_;
  always @(posedge nvdla_core_clk)
      dl_out_data90 <= _0359_;
  always @(posedge nvdla_core_clk)
      dl_out_data89 <= _0357_;
  always @(posedge nvdla_core_clk)
      dl_out_data88 <= _0356_;
  always @(posedge nvdla_core_clk)
      dl_out_data87 <= _0355_;
  always @(posedge nvdla_core_clk)
      dl_out_data86 <= _0354_;
  always @(posedge nvdla_core_clk)
      dl_out_data85 <= _0353_;
  always @(posedge nvdla_core_clk)
      dl_out_data84 <= _0352_;
  always @(posedge nvdla_core_clk)
      dl_out_data83 <= _0351_;
  always @(posedge nvdla_core_clk)
      dl_out_data82 <= _0350_;
  always @(posedge nvdla_core_clk)
      dl_out_data81 <= _0349_;
  always @(posedge nvdla_core_clk)
      dl_out_data80 <= _0348_;
  always @(posedge nvdla_core_clk)
      dl_out_data79 <= _0346_;
  always @(posedge nvdla_core_clk)
      dl_out_data78 <= _0345_;
  always @(posedge nvdla_core_clk)
      dl_out_data77 <= _0344_;
  always @(posedge nvdla_core_clk)
      dl_out_data76 <= _0343_;
  always @(posedge nvdla_core_clk)
      dl_out_data75 <= _0342_;
  always @(posedge nvdla_core_clk)
      dl_out_data74 <= _0341_;
  always @(posedge nvdla_core_clk)
      dl_out_data73 <= _0340_;
  always @(posedge nvdla_core_clk)
      dl_out_data72 <= _0339_;
  always @(posedge nvdla_core_clk)
      dl_out_data71 <= _0338_;
  always @(posedge nvdla_core_clk)
      dl_out_data70 <= _0337_;
  always @(posedge nvdla_core_clk)
      dl_out_data69 <= _0335_;
  always @(posedge nvdla_core_clk)
      dl_out_data68 <= _0334_;
  always @(posedge nvdla_core_clk)
      dl_out_data67 <= _0333_;
  always @(posedge nvdla_core_clk)
      dl_out_data66 <= _0332_;
  always @(posedge nvdla_core_clk)
      dl_out_data65 <= _0331_;
  always @(posedge nvdla_core_clk)
      dl_out_data64 <= _0330_;
  always @(posedge nvdla_core_clk)
      dl_out_data63 <= _0329_;
  always @(posedge nvdla_core_clk)
      dl_out_data62 <= _0328_;
  always @(posedge nvdla_core_clk)
      dl_out_data61 <= _0327_;
  always @(posedge nvdla_core_clk)
      dl_out_data60 <= _0326_;
  always @(posedge nvdla_core_clk)
      dl_out_data59 <= _0324_;
  always @(posedge nvdla_core_clk)
      dl_out_data58 <= _0323_;
  always @(posedge nvdla_core_clk)
      dl_out_data57 <= _0322_;
  always @(posedge nvdla_core_clk)
      dl_out_data56 <= _0321_;
  always @(posedge nvdla_core_clk)
      dl_out_data55 <= _0320_;
  always @(posedge nvdla_core_clk)
      dl_out_data54 <= _0319_;
  always @(posedge nvdla_core_clk)
      dl_out_data53 <= _0318_;
  always @(posedge nvdla_core_clk)
      dl_out_data52 <= _0317_;
  always @(posedge nvdla_core_clk)
      dl_out_data51 <= _0316_;
  always @(posedge nvdla_core_clk)
      dl_out_data50 <= _0315_;
  always @(posedge nvdla_core_clk)
      dl_out_data49 <= _0313_;
  always @(posedge nvdla_core_clk)
      dl_out_data48 <= _0312_;
  always @(posedge nvdla_core_clk)
      dl_out_data47 <= _0311_;
  always @(posedge nvdla_core_clk)
      dl_out_data46 <= _0310_;
  always @(posedge nvdla_core_clk)
      dl_out_data45 <= _0309_;
  always @(posedge nvdla_core_clk)
      dl_out_data44 <= _0308_;
  always @(posedge nvdla_core_clk)
      dl_out_data43 <= _0307_;
  always @(posedge nvdla_core_clk)
      dl_out_data42 <= _0306_;
  always @(posedge nvdla_core_clk)
      dl_out_data41 <= _0305_;
  always @(posedge nvdla_core_clk)
      dl_out_data40 <= _0304_;
  always @(posedge nvdla_core_clk)
      dl_out_data39 <= _0302_;
  always @(posedge nvdla_core_clk)
      dl_out_data38 <= _0301_;
  always @(posedge nvdla_core_clk)
      dl_out_data37 <= _0300_;
  always @(posedge nvdla_core_clk)
      dl_out_data36 <= _0299_;
  always @(posedge nvdla_core_clk)
      dl_out_data35 <= _0298_;
  always @(posedge nvdla_core_clk)
      dl_out_data34 <= _0297_;
  always @(posedge nvdla_core_clk)
      dl_out_data33 <= _0296_;
  always @(posedge nvdla_core_clk)
      dl_out_data32 <= _0295_;
  always @(posedge nvdla_core_clk)
      dl_out_data31 <= _0294_;
  always @(posedge nvdla_core_clk)
      dl_out_data30 <= _0293_;
  always @(posedge nvdla_core_clk)
      dl_out_data29 <= _0291_;
  always @(posedge nvdla_core_clk)
      dl_out_data28 <= _0290_;
  always @(posedge nvdla_core_clk)
      dl_out_data27 <= _0289_;
  always @(posedge nvdla_core_clk)
      dl_out_data26 <= _0288_;
  always @(posedge nvdla_core_clk)
      dl_out_data25 <= _0287_;
  always @(posedge nvdla_core_clk)
      dl_out_data24 <= _0286_;
  always @(posedge nvdla_core_clk)
      dl_out_data23 <= _0285_;
  always @(posedge nvdla_core_clk)
      dl_out_data22 <= _0284_;
  always @(posedge nvdla_core_clk)
      dl_out_data21 <= _0283_;
  always @(posedge nvdla_core_clk)
      dl_out_data20 <= _0282_;
  always @(posedge nvdla_core_clk)
      dl_out_data19 <= _0280_;
  always @(posedge nvdla_core_clk)
      dl_out_data18 <= _0279_;
  always @(posedge nvdla_core_clk)
      dl_out_data17 <= _0278_;
  always @(posedge nvdla_core_clk)
      dl_out_data16 <= _0277_;
  always @(posedge nvdla_core_clk)
      dl_out_data15 <= _0276_;
  always @(posedge nvdla_core_clk)
      dl_out_data14 <= _0275_;
  always @(posedge nvdla_core_clk)
      dl_out_data13 <= _0274_;
  always @(posedge nvdla_core_clk)
      dl_out_data12 <= _0273_;
  always @(posedge nvdla_core_clk)
      dl_out_data11 <= _0264_;
  always @(posedge nvdla_core_clk)
      dl_out_data10 <= _0253_;
  always @(posedge nvdla_core_clk)
      dl_out_data9 <= _0369_;
  always @(posedge nvdla_core_clk)
      dl_out_data8 <= _0358_;
  always @(posedge nvdla_core_clk)
      dl_out_data7 <= _0347_;
  always @(posedge nvdla_core_clk)
      dl_out_data6 <= _0336_;
  always @(posedge nvdla_core_clk)
      dl_out_data5 <= _0325_;
  always @(posedge nvdla_core_clk)
      dl_out_data4 <= _0314_;
  always @(posedge nvdla_core_clk)
      dl_out_data3 <= _0303_;
  always @(posedge nvdla_core_clk)
      dl_out_data2 <= _0292_;
  always @(posedge nvdla_core_clk)
      dl_out_data1 <= _0281_;
  always @(posedge nvdla_core_clk)
      dl_out_data0 <= _0242_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      dl_out_flag <= 9'b000000000;
    else
      dl_out_flag <= _0370_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      dl_out_mask <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    else
      dl_out_mask <= _0371_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      dl_out_pvld <= 1'b0;
    else
      dl_out_pvld <= dat_out_pvld;
  always @(posedge nvdla_core_clk)
      dat_rsp_wg_ch3_d1 <= _0222_;
  always @(posedge nvdla_core_clk)
      dat_rsp_wg_ch2_d1 <= _0221_;
  always @(posedge nvdla_core_clk)
      dat_rsp_wg_ch1_d1 <= _0220_;
  always @(posedge nvdla_core_clk)
      dat_rsp_wg_ch0_d1 <= _0219_;
  reg [0:0] \dat_rsp_pra_en_d1_reg[0] ;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      \dat_rsp_pra_en_d1_reg[0]  <= 1'b0;
    else
      \dat_rsp_pra_en_d1_reg[0]  <= dat_rsp_pra_en;
  assign dat_rsp_pra_en_d1[0] = \dat_rsp_pra_en_d1_reg[0] ;
  always @(posedge nvdla_core_clk)
      dat_out_bypass_data[1023:1016] <= _0025_;
  always @(posedge nvdla_core_clk)
      dat_out_bypass_data[1015:1008] <= _0024_;
  always @(posedge nvdla_core_clk)
      dat_out_bypass_data[1007:1000] <= _0023_;
  always @(posedge nvdla_core_clk)
      dat_out_bypass_data[999:992] <= _0150_;
  always @(posedge nvdla_core_clk)
      dat_out_bypass_data[991:984] <= _0149_;
  always @(posedge nvdla_core_clk)
      dat_out_bypass_data[983:976] <= _0148_;
  always @(posedge nvdla_core_clk)
      dat_out_bypass_data[975:968] <= _0147_;
  always @(posedge nvdla_core_clk)
      dat_out_bypass_data[967:960] <= _0146_;
  always @(posedge nvdla_core_clk)
      dat_out_bypass_data[959:952] <= _0144_;
  always @(posedge nvdla_core_clk)
      dat_out_bypass_data[951:944] <= _0143_;
  always @(posedge nvdla_core_clk)
      dat_out_bypass_data[943:936] <= _0142_;
  always @(posedge nvdla_core_clk)
      dat_out_bypass_data[935:928] <= _0141_;
  always @(posedge nvdla_core_clk)
      dat_out_bypass_data[927:920] <= _0140_;
  always @(posedge nvdla_core_clk)
      dat_out_bypass_data[919:912] <= _0139_;
  always @(posedge nvdla_core_clk)
      dat_out_bypass_data[911:904] <= _0138_;
  always @(posedge nvdla_core_clk)
      dat_out_bypass_data[903:896] <= _0137_;
  always @(posedge nvdla_core_clk)
      dat_out_bypass_data[895:888] <= _0136_;
  always @(posedge nvdla_core_clk)
      dat_out_bypass_data[887:880] <= _0135_;
  always @(posedge nvdla_core_clk)
      dat_out_bypass_data[879:872] <= _0133_;
  always @(posedge nvdla_core_clk)
      dat_out_bypass_data[871:864] <= _0132_;
  always @(posedge nvdla_core_clk)
      dat_out_bypass_data[863:856] <= _0131_;
  always @(posedge nvdla_core_clk)
      dat_out_bypass_data[855:848] <= _0130_;
  always @(posedge nvdla_core_clk)
      dat_out_bypass_data[847:840] <= _0129_;
  always @(posedge nvdla_core_clk)
      dat_out_bypass_data[839:832] <= _0128_;
  always @(posedge nvdla_core_clk)
      dat_out_bypass_data[831:824] <= _0127_;
  always @(posedge nvdla_core_clk)
      dat_out_bypass_data[823:816] <= _0126_;
  always @(posedge nvdla_core_clk)
      dat_out_bypass_data[815:808] <= _0125_;
  always @(posedge nvdla_core_clk)
      dat_out_bypass_data[807:800] <= _0124_;
  always @(posedge nvdla_core_clk)
      dat_out_bypass_data[799:792] <= _0121_;
  always @(posedge nvdla_core_clk)
      dat_out_bypass_data[791:784] <= _0120_;
  always @(posedge nvdla_core_clk)
      dat_out_bypass_data[783:776] <= _0119_;
  always @(posedge nvdla_core_clk)
      dat_out_bypass_data[775:768] <= _0118_;
  always @(posedge nvdla_core_clk)
      dat_out_bypass_data[767:760] <= _0117_;
  always @(posedge nvdla_core_clk)
      dat_out_bypass_data[759:752] <= _0116_;
  always @(posedge nvdla_core_clk)
      dat_out_bypass_data[751:744] <= _0115_;
  always @(posedge nvdla_core_clk)
      dat_out_bypass_data[743:736] <= _0114_;
  always @(posedge nvdla_core_clk)
      dat_out_bypass_data[735:728] <= _0113_;
  always @(posedge nvdla_core_clk)
      dat_out_bypass_data[727:720] <= _0112_;
  always @(posedge nvdla_core_clk)
      dat_out_bypass_data[719:712] <= _0110_;
  always @(posedge nvdla_core_clk)
      dat_out_bypass_data[711:704] <= _0109_;
  always @(posedge nvdla_core_clk)
      dat_out_bypass_data[703:696] <= _0108_;
  always @(posedge nvdla_core_clk)
      dat_out_bypass_data[695:688] <= _0107_;
  always @(posedge nvdla_core_clk)
      dat_out_bypass_data[687:680] <= _0106_;
  always @(posedge nvdla_core_clk)
      dat_out_bypass_data[679:672] <= _0105_;
  always @(posedge nvdla_core_clk)
      dat_out_bypass_data[671:664] <= _0104_;
  always @(posedge nvdla_core_clk)
      dat_out_bypass_data[663:656] <= _0103_;
  always @(posedge nvdla_core_clk)
      dat_out_bypass_data[655:648] <= _0102_;
  always @(posedge nvdla_core_clk)
      dat_out_bypass_data[647:640] <= _0101_;
  always @(posedge nvdla_core_clk)
      dat_out_bypass_data[639:632] <= _0099_;
  always @(posedge nvdla_core_clk)
      dat_out_bypass_data[631:624] <= _0098_;
  always @(posedge nvdla_core_clk)
      dat_out_bypass_data[623:616] <= _0097_;
  always @(posedge nvdla_core_clk)
      dat_out_bypass_data[615:608] <= _0096_;
  always @(posedge nvdla_core_clk)
      dat_out_bypass_data[607:600] <= _0095_;
  always @(posedge nvdla_core_clk)
      dat_out_bypass_data[599:592] <= _0094_;
  always @(posedge nvdla_core_clk)
      dat_out_bypass_data[591:584] <= _0093_;
  always @(posedge nvdla_core_clk)
      dat_out_bypass_data[583:576] <= _0092_;
  always @(posedge nvdla_core_clk)
      dat_out_bypass_data[575:568] <= _0091_;
  always @(posedge nvdla_core_clk)
      dat_out_bypass_data[567:560] <= _0090_;
  always @(posedge nvdla_core_clk)
      dat_out_bypass_data[559:552] <= _0088_;
  always @(posedge nvdla_core_clk)
      dat_out_bypass_data[551:544] <= _0087_;
  always @(posedge nvdla_core_clk)
      dat_out_bypass_data[543:536] <= _0086_;
  always @(posedge nvdla_core_clk)
      dat_out_bypass_data[535:528] <= _0085_;
  always @(posedge nvdla_core_clk)
      dat_out_bypass_data[527:520] <= _0084_;
  always @(posedge nvdla_core_clk)
      dat_out_bypass_data[519:512] <= _0083_;
  always @(posedge nvdla_core_clk)
      dat_out_bypass_data[511:504] <= _0082_;
  always @(posedge nvdla_core_clk)
      dat_out_bypass_data[503:496] <= _0081_;
  always @(posedge nvdla_core_clk)
      dat_out_bypass_data[495:488] <= _0080_;
  always @(posedge nvdla_core_clk)
      dat_out_bypass_data[487:480] <= _0079_;
  always @(posedge nvdla_core_clk)
      dat_out_bypass_data[479:472] <= _0077_;
  always @(posedge nvdla_core_clk)
      dat_out_bypass_data[471:464] <= _0076_;
  always @(posedge nvdla_core_clk)
      dat_out_bypass_data[463:456] <= _0075_;
  always @(posedge nvdla_core_clk)
      dat_out_bypass_data[455:448] <= _0074_;
  always @(posedge nvdla_core_clk)
      dat_out_bypass_data[447:440] <= _0073_;
  always @(posedge nvdla_core_clk)
      dat_out_bypass_data[439:432] <= _0072_;
  always @(posedge nvdla_core_clk)
      dat_out_bypass_data[431:424] <= _0071_;
  always @(posedge nvdla_core_clk)
      dat_out_bypass_data[423:416] <= _0070_;
  always @(posedge nvdla_core_clk)
      dat_out_bypass_data[415:408] <= _0069_;
  always @(posedge nvdla_core_clk)
      dat_out_bypass_data[407:400] <= _0068_;
  always @(posedge nvdla_core_clk)
      dat_out_bypass_data[399:392] <= _0066_;
  always @(posedge nvdla_core_clk)
      dat_out_bypass_data[391:384] <= _0065_;
  always @(posedge nvdla_core_clk)
      dat_out_bypass_data[383:376] <= _0064_;
  always @(posedge nvdla_core_clk)
      dat_out_bypass_data[375:368] <= _0063_;
  always @(posedge nvdla_core_clk)
      dat_out_bypass_data[367:360] <= _0062_;
  always @(posedge nvdla_core_clk)
      dat_out_bypass_data[359:352] <= _0061_;
  always @(posedge nvdla_core_clk)
      dat_out_bypass_data[351:344] <= _0060_;
  always @(posedge nvdla_core_clk)
      dat_out_bypass_data[343:336] <= _0059_;
  always @(posedge nvdla_core_clk)
      dat_out_bypass_data[335:328] <= _0058_;
  always @(posedge nvdla_core_clk)
      dat_out_bypass_data[327:320] <= _0057_;
  always @(posedge nvdla_core_clk)
      dat_out_bypass_data[319:312] <= _0055_;
  always @(posedge nvdla_core_clk)
      dat_out_bypass_data[311:304] <= _0054_;
  always @(posedge nvdla_core_clk)
      dat_out_bypass_data[303:296] <= _0053_;
  always @(posedge nvdla_core_clk)
      dat_out_bypass_data[295:288] <= _0052_;
  always @(posedge nvdla_core_clk)
      dat_out_bypass_data[287:280] <= _0051_;
  always @(posedge nvdla_core_clk)
      dat_out_bypass_data[279:272] <= _0050_;
  always @(posedge nvdla_core_clk)
      dat_out_bypass_data[271:264] <= _0049_;
  always @(posedge nvdla_core_clk)
      dat_out_bypass_data[263:256] <= _0048_;
  always @(posedge nvdla_core_clk)
      dat_out_bypass_data[255:248] <= _0047_;
  always @(posedge nvdla_core_clk)
      dat_out_bypass_data[247:240] <= _0046_;
  always @(posedge nvdla_core_clk)
      dat_out_bypass_data[239:232] <= _0044_;
  always @(posedge nvdla_core_clk)
      dat_out_bypass_data[231:224] <= _0043_;
  always @(posedge nvdla_core_clk)
      dat_out_bypass_data[223:216] <= _0042_;
  always @(posedge nvdla_core_clk)
      dat_out_bypass_data[215:208] <= _0041_;
  always @(posedge nvdla_core_clk)
      dat_out_bypass_data[207:200] <= _0040_;
  always @(posedge nvdla_core_clk)
      dat_out_bypass_data[199:192] <= _0039_;
  always @(posedge nvdla_core_clk)
      dat_out_bypass_data[191:184] <= _0038_;
  always @(posedge nvdla_core_clk)
      dat_out_bypass_data[183:176] <= _0037_;
  always @(posedge nvdla_core_clk)
      dat_out_bypass_data[175:168] <= _0036_;
  always @(posedge nvdla_core_clk)
      dat_out_bypass_data[167:160] <= _0035_;
  always @(posedge nvdla_core_clk)
      dat_out_bypass_data[159:152] <= _0033_;
  always @(posedge nvdla_core_clk)
      dat_out_bypass_data[151:144] <= _0032_;
  always @(posedge nvdla_core_clk)
      dat_out_bypass_data[143:136] <= _0031_;
  always @(posedge nvdla_core_clk)
      dat_out_bypass_data[135:128] <= _0030_;
  always @(posedge nvdla_core_clk)
      dat_out_bypass_data[127:120] <= _0029_;
  always @(posedge nvdla_core_clk)
      dat_out_bypass_data[119:112] <= _0028_;
  always @(posedge nvdla_core_clk)
      dat_out_bypass_data[111:104] <= _0027_;
  always @(posedge nvdla_core_clk)
      dat_out_bypass_data[103:96] <= _0026_;
  always @(posedge nvdla_core_clk)
      dat_out_bypass_data[95:88] <= _0145_;
  always @(posedge nvdla_core_clk)
      dat_out_bypass_data[87:80] <= _0134_;
  always @(posedge nvdla_core_clk)
      dat_out_bypass_data[79:72] <= _0122_;
  always @(posedge nvdla_core_clk)
      dat_out_bypass_data[71:64] <= _0111_;
  always @(posedge nvdla_core_clk)
      dat_out_bypass_data[63:56] <= _0100_;
  always @(posedge nvdla_core_clk)
      dat_out_bypass_data[55:48] <= _0089_;
  always @(posedge nvdla_core_clk)
      dat_out_bypass_data[47:40] <= _0078_;
  always @(posedge nvdla_core_clk)
      dat_out_bypass_data[39:32] <= _0067_;
  always @(posedge nvdla_core_clk)
      dat_out_bypass_data[31:24] <= _0056_;
  always @(posedge nvdla_core_clk)
      dat_out_bypass_data[23:16] <= _0045_;
  always @(posedge nvdla_core_clk)
      dat_out_bypass_data[15:8] <= _0034_;
  always @(posedge nvdla_core_clk)
      dat_out_bypass_data[7:0] <= _0123_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      dat_out_bypass_mask[127:64] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    else
      dat_out_bypass_mask[127:64] <= _0151_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      dat_out_bypass_mask[63:0] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    else
      dat_out_bypass_mask[63:0] <= _0152_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      dat_out_flag <= 9'b000000000;
    else
      dat_out_flag <= _0153_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      dat_out_pvld <= 1'b0;
    else
      dat_out_pvld <= dat_out_pvld_w;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      dat_out_flag_l5 <= 9'b000000000;
    else
      dat_out_flag_l5 <= _0158_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      dat_out_pvld_l5 <= 1'b0;
    else
      dat_out_pvld_l5 <= dat_out_pvld_l4;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      dat_out_flag_l4 <= 9'b000000000;
    else
      dat_out_flag_l4 <= _0157_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      dat_out_pvld_l4 <= 1'b0;
    else
      dat_out_pvld_l4 <= dat_out_pvld_l3;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      dat_out_flag_l3 <= 9'b000000000;
    else
      dat_out_flag_l3 <= _0156_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      dat_out_pvld_l3 <= 1'b0;
    else
      dat_out_pvld_l3 <= dat_out_pvld_l2;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      dat_out_flag_l2 <= 9'b000000000;
    else
      dat_out_flag_l2 <= _0155_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      dat_out_pvld_l2 <= 1'b0;
    else
      dat_out_pvld_l2 <= dat_out_pvld_l1;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      dat_out_flag_l1 <= 9'b000000000;
    else
      dat_out_flag_l1 <= _0154_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      dat_out_pvld_l1 <= 1'b0;
    else
      dat_out_pvld_l1 <= dat_rsp_pvld;
  always @(posedge nvdla_core_clk)
      dat_rsp_l2_sft_d3[255:128] <= _0208_;
  always @(posedge nvdla_core_clk)
      dat_rsp_l2_sft_d3[127:0] <= _0207_;
  always @(posedge nvdla_core_clk)
      dat_rsp_l1_sft_d3[255:128] <= _0206_;
  always @(posedge nvdla_core_clk)
      dat_rsp_l1_sft_d3[127:0] <= _0205_;
  always @(posedge nvdla_core_clk)
      dat_rsp_l1_sft_d2[255:128] <= _0204_;
  always @(posedge nvdla_core_clk)
      dat_rsp_l1_sft_d2[127:0] <= _0203_;
  always @(posedge nvdla_core_clk)
      dat_rsp_l0_sft_d3[255:128] <= _0202_;
  always @(posedge nvdla_core_clk)
      dat_rsp_l0_sft_d3[127:0] <= _0201_;
  always @(posedge nvdla_core_clk)
      dat_rsp_l0_sft_d2[255:128] <= _0200_;
  always @(posedge nvdla_core_clk)
      dat_rsp_l0_sft_d2[127:0] <= _0199_;
  always @(posedge nvdla_core_clk)
      dat_rsp_l0_sft_d1[511:256] <= _0198_;
  always @(posedge nvdla_core_clk)
      dat_rsp_l0_sft_d1[255:0] <= _0197_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      rsp_sft_cnt_l3_ori <= 8'b00000000;
    else
      rsp_sft_cnt_l3_ori <= _0419_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      rsp_sft_cnt_l2_ori <= 8'b00000000;
    else
      rsp_sft_cnt_l2_ori <= _0417_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      rsp_sft_cnt_l1_ori <= 8'b00000000;
    else
      rsp_sft_cnt_l1_ori <= _0415_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      rsp_sft_cnt_l0_ori <= 8'b00000000;
    else
      rsp_sft_cnt_l0_ori <= _0413_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      rsp_sft_cnt_l3 <= 8'b00000000;
    else
      rsp_sft_cnt_l3 <= _0418_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      rsp_sft_cnt_l2 <= 8'b00000000;
    else
      rsp_sft_cnt_l2 <= _0416_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      rsp_sft_cnt_l1 <= 8'b00000000;
    else
      rsp_sft_cnt_l1 <= _0414_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      rsp_sft_cnt_l0 <= 8'b00000000;
    else
      rsp_sft_cnt_l0 <= _0412_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      dat_rsp_pd_d4 <= 27'b000000000000000000000000000;
    else
      dat_rsp_pd_d4 <= _0212_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      dat_rsp_pvld_d4 <= 1'b0;
    else
      dat_rsp_pvld_d4 <= dat_rsp_pvld_d3;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      dat_rsp_pd_d3 <= 27'b000000000000000000000000000;
    else
      dat_rsp_pd_d3 <= _0211_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      dat_rsp_pvld_d3 <= 1'b0;
    else
      dat_rsp_pvld_d3 <= dat_rsp_pvld_d2;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      dat_rsp_pd_d2 <= 27'b000000000000000000000000000;
    else
      dat_rsp_pd_d2 <= _0210_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      dat_rsp_pvld_d2 <= 1'b0;
    else
      dat_rsp_pvld_d2 <= dat_rsp_pvld_d1;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      dat_rsp_pd_d1 <= 27'b000000000000000000000000000;
    else
      dat_rsp_pd_d1 <= _0209_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      dat_rsp_pvld_d1 <= 1'b0;
    else
      dat_rsp_pvld_d1 <= dat_rsp_pipe_pvld_d6;
  always @(posedge nvdla_core_clk)
      dat_l3c1_hi <= _0021_;
  always @(posedge nvdla_core_clk)
      dat_l3c1_lo <= _0022_;
  always @(posedge nvdla_core_clk)
      dat_l2c1_hi <= _0017_;
  always @(posedge nvdla_core_clk)
      dat_l2c1_lo <= _0018_;
  always @(posedge nvdla_core_clk)
      dat_l1c1_hi <= _0013_;
  always @(posedge nvdla_core_clk)
      dat_l1c1_lo <= _0014_;
  always @(posedge nvdla_core_clk)
      dat_l0c1_hi <= _0009_;
  always @(posedge nvdla_core_clk)
      dat_l0c1_lo <= _0010_;
  always @(posedge nvdla_core_clk)
      dat_l3c0_hi <= _0019_;
  always @(posedge nvdla_core_clk)
      dat_l3c0_lo <= _0020_;
  always @(posedge nvdla_core_clk)
      dat_l2c0_hi <= _0015_;
  always @(posedge nvdla_core_clk)
      dat_l2c0_lo <= _0016_;
  always @(posedge nvdla_core_clk)
      dat_l1c0_hi <= _0011_;
  always @(posedge nvdla_core_clk)
      dat_l1c0_lo <= _0012_;
  always @(posedge nvdla_core_clk)
      dat_l0c0_hi <= _0007_;
  always @(posedge nvdla_core_clk)
      dat_l0c0_lo <= _0008_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      dat_l3c1_dummy <= 1'b1;
    else
      dat_l3c1_dummy <= dat_l3c1_dummy_w;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      dat_l2c1_dummy <= 1'b1;
    else
      dat_l2c1_dummy <= dat_l2c1_dummy_w;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      dat_l1c1_dummy <= 1'b1;
    else
      dat_l1c1_dummy <= dat_l1c1_dummy_w;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      dat_l0c1_dummy <= 1'b1;
    else
      dat_l0c1_dummy <= dat_l0c1_dummy_w;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      dat_l3c0_dummy <= 1'b1;
    else
      dat_l3c0_dummy <= dat_l3c0_dummy_w;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      dat_l2c0_dummy <= 1'b1;
    else
      dat_l2c0_dummy <= dat_l2c0_dummy_w;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      dat_l1c0_dummy <= 1'b1;
    else
      dat_l1c0_dummy <= dat_l1c0_dummy_w;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      dat_l0c0_dummy <= 1'b1;
    else
      dat_l0c0_dummy <= dat_l0c0_dummy_w;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      dat_rsp_exec_sub_h_d6 <= 2'b00;
    else
      dat_rsp_exec_sub_h_d6 <= _0196_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      dat_rsp_exec_dummy_d6 <= 1'b0;
    else
      dat_rsp_exec_dummy_d6 <= _0190_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      dat_rsp_exec_pvld_d6 <= 1'b0;
    else
      dat_rsp_exec_pvld_d6 <= dat_rsp_exec_pvld_d5;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      dat_rsp_pipe_pd_d6 <= 29'b00000000000000000000000000000;
    else
      dat_rsp_pipe_pd_d6 <= _0218_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      dat_rsp_pipe_pvld_d6 <= 1'b0;
    else
      dat_rsp_pipe_pvld_d6 <= dat_rsp_pipe_pvld_d5;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      dat_rsp_exec_sub_h_d5 <= 2'b00;
    else
      dat_rsp_exec_sub_h_d5 <= _0195_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      dat_rsp_exec_dummy_d5 <= 1'b0;
    else
      dat_rsp_exec_dummy_d5 <= _0189_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      dat_rsp_exec_pvld_d5 <= 1'b0;
    else
      dat_rsp_exec_pvld_d5 <= dat_rsp_exec_pvld_d4;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      dat_rsp_pipe_pd_d5 <= 29'b00000000000000000000000000000;
    else
      dat_rsp_pipe_pd_d5 <= _0217_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      dat_rsp_pipe_pvld_d5 <= 1'b0;
    else
      dat_rsp_pipe_pvld_d5 <= dat_rsp_pipe_pvld_d4;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      dat_rsp_exec_sub_h_d4 <= 2'b00;
    else
      dat_rsp_exec_sub_h_d4 <= _0194_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      dat_rsp_exec_dummy_d4 <= 1'b0;
    else
      dat_rsp_exec_dummy_d4 <= _0188_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      dat_rsp_exec_pvld_d4 <= 1'b0;
    else
      dat_rsp_exec_pvld_d4 <= dat_rsp_exec_pvld_d3;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      dat_rsp_pipe_pd_d4 <= 29'b00000000000000000000000000000;
    else
      dat_rsp_pipe_pd_d4 <= _0216_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      dat_rsp_pipe_pvld_d4 <= 1'b0;
    else
      dat_rsp_pipe_pvld_d4 <= dat_rsp_pipe_pvld_d3;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      dat_rsp_exec_sub_h_d3 <= 2'b00;
    else
      dat_rsp_exec_sub_h_d3 <= _0193_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      dat_rsp_exec_dummy_d3 <= 1'b0;
    else
      dat_rsp_exec_dummy_d3 <= _0187_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      dat_rsp_exec_pvld_d3 <= 1'b0;
    else
      dat_rsp_exec_pvld_d3 <= dat_rsp_exec_pvld_d2;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      dat_rsp_pipe_pd_d3 <= 29'b00000000000000000000000000000;
    else
      dat_rsp_pipe_pd_d3 <= _0215_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      dat_rsp_pipe_pvld_d3 <= 1'b0;
    else
      dat_rsp_pipe_pvld_d3 <= dat_rsp_pipe_pvld_d2;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      dat_rsp_exec_sub_h_d2 <= 2'b00;
    else
      dat_rsp_exec_sub_h_d2 <= _0192_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      dat_rsp_exec_dummy_d2 <= 1'b0;
    else
      dat_rsp_exec_dummy_d2 <= _0186_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      dat_rsp_exec_pvld_d2 <= 1'b0;
    else
      dat_rsp_exec_pvld_d2 <= dat_rsp_exec_pvld_d1;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      dat_rsp_pipe_pd_d2 <= 29'b00000000000000000000000000000;
    else
      dat_rsp_pipe_pd_d2 <= _0214_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      dat_rsp_pipe_pvld_d2 <= 1'b0;
    else
      dat_rsp_pipe_pvld_d2 <= dat_rsp_pipe_pvld_d1;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      dat_rsp_exec_sub_h_d1 <= 2'b00;
    else
      dat_rsp_exec_sub_h_d1 <= _0191_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      dat_rsp_exec_dummy_d1 <= 1'b0;
    else
      dat_rsp_exec_dummy_d1 <= _0185_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      dat_rsp_exec_pvld_d1 <= 1'b0;
    else
      dat_rsp_exec_pvld_d1 <= dat_exec_valid_d2;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      dat_rsp_pipe_pd_d1 <= 29'b00000000000000000000000000000;
    else
      dat_rsp_pipe_pd_d1 <= _0213_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      dat_rsp_pipe_pvld_d1 <= 1'b0;
    else
      dat_rsp_pipe_pvld_d1 <= dat_pipe_valid_d2;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      dat_req_flag_d2 <= 9'b000000000;
    else
      dat_req_flag_d2 <= _0170_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      dat_req_rls_d2 <= 1'b0;
    else
      dat_req_rls_d2 <= _0172_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      dat_req_sub_w_st_d2 <= 1'b0;
    else
      dat_req_sub_w_st_d2 <= _0184_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      dat_req_cur_sub_h_d2 <= 2'b00;
    else
      dat_req_cur_sub_h_d2 <= _0166_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      dat_req_dummy_d2 <= 1'b0;
    else
      dat_req_dummy_d2 <= _0168_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      dat_req_bytes_d2 <= 8'b00000000;
    else
      dat_req_bytes_d2 <= _0160_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      dat_req_ch_odd_d2 <= 1'b0;
    else
      dat_req_ch_odd_d2 <= _0164_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      dat_req_ch_end_d2 <= 1'b0;
    else
      dat_req_ch_end_d2 <= _0162_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      dat_req_sub_c_d2 <= 1'b0;
    else
      dat_req_sub_c_d2 <= _0174_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      dat_req_sub_h_d2 <= 2'b00;
    else
      dat_req_sub_h_d2 <= _0180_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      dat_req_sub_w_d2 <= 2'b00;
    else
      dat_req_sub_w_d2 <= _0182_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      dat_exec_valid_d2 <= 1'b0;
    else
      dat_exec_valid_d2 <= dat_exec_valid_d1;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      dat_pipe_valid_d2 <= 1'b0;
    else
      dat_pipe_valid_d2 <= dat_pipe_valid_d1;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      sc2buf_dat_rd_addr <= 12'b111111111111;
    else
      sc2buf_dat_rd_addr <= _0420_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      sc2buf_dat_rd_en <= 1'b0;
    else
      sc2buf_dat_rd_en <= sc2buf_dat_rd_en_w;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      dat_req_sub_h_3_addr <= 12'b111111111111;
    else
      dat_req_sub_h_3_addr <= _0178_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      dat_req_sub_h_2_addr <= 12'b111111111111;
    else
      dat_req_sub_h_2_addr <= _0177_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      dat_req_sub_h_1_addr <= 12'b111111111111;
    else
      dat_req_sub_h_1_addr <= _0176_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      dat_req_sub_h_0_addr <= 12'b111111111111;
    else
      dat_req_sub_h_0_addr <= _0175_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      w_bias_d1 <= 12'b000000000000;
    else
      w_bias_d1 <= _0700_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      h_bias_3_d1 <= 12'b000000000000;
    else
      h_bias_3_d1 <= _0385_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      h_bias_2_d1 <= 12'b000000000000;
    else
      h_bias_2_d1 <= _0383_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      h_bias_1_d1 <= 12'b000000000000;
    else
      h_bias_1_d1 <= _0381_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      h_bias_0_d1 <= 12'b000000000000;
    else
      h_bias_0_d1 <= _0379_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      c_bias_d1 <= 12'b000000000000;
    else
      c_bias_d1 <= _0003_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      c_bias <= 12'b000000000000;
    else
      c_bias <= _0002_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      pixel_force_clr_d1 <= 1'b0;
    else
      pixel_force_clr_d1 <= _0396_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      pixel_force_fetch_d1 <= 1'b0;
    else
      pixel_force_fetch_d1 <= _0397_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      dat_req_rls_d1 <= 1'b0;
    else
      dat_req_rls_d1 <= _0171_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      dat_req_flag_d1 <= 9'b000000000;
    else
      dat_req_flag_d1 <= _0169_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      dat_req_sub_w_st_d1 <= 1'b0;
    else
      dat_req_sub_w_st_d1 <= _0183_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      dat_req_cur_sub_h_d1 <= 2'b00;
    else
      dat_req_cur_sub_h_d1 <= _0165_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      dat_req_dummy_d1 <= 1'b0;
    else
      dat_req_dummy_d1 <= _0167_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      dat_req_ch_odd_d1 <= 1'b0;
    else
      dat_req_ch_odd_d1 <= _0163_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      dat_req_ch_end_d1 <= 1'b0;
    else
      dat_req_ch_end_d1 <= _0161_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      dat_req_sub_c_d1 <= 1'b0;
    else
      dat_req_sub_c_d1 <= _0173_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      dat_req_sub_h_d1 <= 2'b00;
    else
      dat_req_sub_h_d1 <= _0179_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      dat_req_sub_w_d1 <= 2'b00;
    else
      dat_req_sub_w_d1 <= _0181_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      dat_req_valid_d1 <= 1'b0;
    else
      dat_req_valid_d1 <= dat_req_valid;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      datain_h_ori <= 14'b00000000000000;
    else
      datain_h_ori <= _0228_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      datain_h_cnt <= 14'b00000000000000;
    else
      datain_h_cnt <= _0227_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      pixel_req_ch_odd_ori <= 1'b0;
    else
      pixel_req_ch_odd_ori <= _0399_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      pixel_req_ch_odd <= 1'b0;
    else
      pixel_req_ch_odd <= _0398_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      pixel_w_ch_ori <= 16'b0000000000000000;
    else
      pixel_w_ch_ori <= _0400_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      pixel_w_ori <= 16'b0000000000000000;
    else
      pixel_w_ori <= _0402_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      pixel_w_cnt <= 16'b0000000000000000;
    else
      pixel_w_cnt <= _0401_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      datain_w_ori <= 14'b00000000000000;
    else
      datain_w_ori <= _0231_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      datain_w_cnt <= 14'b00000000000000;
    else
      datain_w_cnt <= _0230_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      datain_c_cnt <= 11'b00000000000;
    else
      datain_c_cnt <= _0225_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      dataout_w_ori <= 13'b0000000000000;
    else
      dataout_w_ori <= _0235_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      dataout_w_cnt <= 13'b0000000000000;
    else
      dataout_w_cnt <= _0234_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      dat_req_bytes_d1 <= 8'b00000000;
    else
      dat_req_bytes_d1 <= _0159_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      dat_exec_valid_d1 <= 1'b0;
    else
      dat_exec_valid_d1 <= dat_exec_valid;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      dat_pipe_valid_d1 <= 1'b0;
    else
      dat_pipe_valid_d1 <= dat_pipe_valid;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      dat_pipe_local_valid <= 1'b0;
    else
      dat_pipe_local_valid <= dat_pipe_local_valid_w;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      stripe_cnt <= 7'b0000000;
    else
      stripe_cnt <= _0684_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      sub_h_cnt <= 2'b00;
    else
      sub_h_cnt <= _0687_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      batch_cnt <= 5'b00000;
    else
      batch_cnt <= _0001_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      dl_pd_d4 <= 31'b0000000000000000000000000000000;
    else
      dl_pd_d4 <= _0375_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      dl_pvld_d4 <= 1'b0;
    else
      dl_pvld_d4 <= dl_pvld_d3;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      dl_pd_d3 <= 31'b0000000000000000000000000000000;
    else
      dl_pd_d3 <= _0374_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      dl_pvld_d3 <= 1'b0;
    else
      dl_pvld_d3 <= dl_pvld_d2;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      dl_pd_d2 <= 31'b0000000000000000000000000000000;
    else
      dl_pd_d2 <= _0373_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      dl_pvld_d2 <= 1'b0;
    else
      dl_pvld_d2 <= dl_pvld_d1;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      dl_pd_d1 <= 31'b0000000000000000000000000000000;
    else
      dl_pd_d1 <= _0372_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      dl_pvld_d1 <= 1'b0;
    else
      dl_pvld_d1 <= dl_in_pvld;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      dl_in_pd_d5 <= 31'b0000000000000000000000000000000;
    else
      dl_in_pd_d5 <= _0241_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      dl_in_pvld_d5 <= 1'b0;
    else
      dl_in_pvld_d5 <= dl_in_pvld_d4;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      dl_in_pd_d4 <= 31'b0000000000000000000000000000000;
    else
      dl_in_pd_d4 <= _0240_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      dl_in_pvld_d4 <= 1'b0;
    else
      dl_in_pvld_d4 <= dl_in_pvld_d3;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      dl_in_pd_d3 <= 31'b0000000000000000000000000000000;
    else
      dl_in_pd_d3 <= _0239_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      dl_in_pvld_d3 <= 1'b0;
    else
      dl_in_pvld_d3 <= dl_in_pvld_d2;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      dl_in_pd_d2 <= 31'b0000000000000000000000000000000;
    else
      dl_in_pd_d2 <= _0238_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      dl_in_pvld_d2 <= 1'b0;
    else
      dl_in_pvld_d2 <= dl_in_pvld_d1;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      dl_in_pd_d1 <= 31'b0000000000000000000000000000000;
    else
      dl_in_pd_d1 <= _0237_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      dl_in_pvld_d1 <= 1'b0;
    else
      dl_in_pvld_d1 <= sg2dl_pvld;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      sc2cdma_dat_entries <= 12'b000000000000;
    else
      sc2cdma_dat_entries <= _0421_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      sc2cdma_dat_slices <= 12'b000000000000;
    else
      sc2cdma_dat_slices <= _0422_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      sc2cdma_dat_updt <= 1'b0;
    else
      sc2cdma_dat_updt <= dat_rls;
  always @(posedge nvdla_core_ng_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      dat_entry_st <= 12'b000000000000;
    else
      dat_entry_st <= _0006_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      slcg_wg_en_d3 <= 1'b0;
    else
      slcg_wg_en_d3 <= slcg_wg_en_d2;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      slcg_wg_en_d2 <= 1'b0;
    else
      slcg_wg_en_d2 <= slcg_wg_en_d1;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      slcg_wg_en_d1 <= 1'b0;
    else
      slcg_wg_en_d1 <= slcg_wg_en_w;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      pra_precision <= 8'b00000000;
    else
      pra_precision <= _0408_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      pra_truncate <= 8'b00000000;
    else
      pra_truncate <= _0409_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      dataout_width_cmp <= 13'b0000000000000;
    else
      dataout_width_cmp <= _0236_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      last_entries <= 12'b000000000000;
    else
      last_entries <= _0392_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      last_slices <= 12'b000000000000;
    else
      last_slices <= _0393_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      slice_left <= 12'b000000000000;
    else
      slice_left <= _0683_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      rls_entries <= 12'b000000000000;
    else
      rls_entries <= _0410_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      rls_slices <= 12'b000000000000;
    else
      rls_slices <= _0411_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      h_bias_3_stride <= 12'b000000000000;
    else
      h_bias_3_stride <= _0386_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      h_bias_2_stride <= 12'b000000000000;
    else
      h_bias_2_stride <= _0384_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      h_bias_1_stride <= 12'b000000000000;
    else
      h_bias_1_stride <= _0382_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      h_bias_0_stride <= 12'b000000000000;
    else
      h_bias_0_stride <= _0380_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      h_offset_slice <= 12'b000000000000;
    else
      h_offset_slice <= _0387_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      entries_cmp <= 12'b000000000000;
    else
      entries_cmp <= _0378_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      entries_batch <= 12'b000000000000;
    else
      entries_batch <= _0377_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      entries <= 12'b000000000000;
    else
      entries <= _0376_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      pad_value <= 16'b0000000000000000;
    else
      pad_value <= _0394_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      y_dilate <= 6'b000000;
    else
      y_dilate <= _0702_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      x_dilate <= 6'b000000;
    else
      x_dilate <= _0701_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      pixel_ch_stride <= 12'b000000000000;
    else
      pixel_ch_stride <= _0395_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      pixel_x_byte_stride <= 7'b0000000;
    else
      pixel_x_byte_stride <= _0404_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      pixel_x_add <= 7'b0000000;
    else
      pixel_x_add <= _0403_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      pixel_x_init_offset <= 7'b0000000;
    else
      pixel_x_init_offset <= _0406_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      pixel_x_init <= 6'b000000;
    else
      pixel_x_init <= _0405_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      batch_cmp <= 5'b00000;
    else
      batch_cmp <= _0000_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      data_batch <= 6'b000000;
    else
      data_batch <= _0224_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      pixel_x_stride_odd <= 1'b0;
    else
      pixel_x_stride_odd <= _0407_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      conv_y_stride <= 4'b0000;
    else
      conv_y_stride <= _0005_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      conv_x_stride <= 4'b0000;
    else
      conv_x_stride <= _0004_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      sub_h_cmp_g1 <= 3'b001;
    else
      sub_h_cmp_g1 <= _0686_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      sub_h_cmp_g0 <= 3'b001;
    else
      sub_h_cmp_g0 <= _0685_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      sub_h_total_g11 <= 3'b001;
    else
      sub_h_total_g11 <= _0690_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      sub_h_total_g10 <= 3'b001;
    else
      sub_h_total_g10 <= _0689_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      sub_h_total_g9 <= 3'b001;
    else
      sub_h_total_g9 <= _0699_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      sub_h_total_g8 <= 3'b001;
    else
      sub_h_total_g8 <= _0698_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      sub_h_total_g7 <= 3'b001;
    else
      sub_h_total_g7 <= _0697_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      sub_h_total_g6 <= 3'b001;
    else
      sub_h_total_g6 <= _0696_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      sub_h_total_g5 <= 3'b001;
    else
      sub_h_total_g5 <= _0695_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      sub_h_total_g4 <= 3'b001;
    else
      sub_h_total_g4 <= _0694_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      sub_h_total_g3 <= 3'b001;
    else
      sub_h_total_g3 <= _0693_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      sub_h_total_g2 <= 2'b01;
    else
      sub_h_total_g2 <= _0692_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      sub_h_total_g1 <= 3'b001;
    else
      sub_h_total_g1 <= _0691_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      sub_h_total_g0 <= 3'b001;
    else
      sub_h_total_g0 <= _0688_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      datain_channel_cmp <= 11'b00000000000;
    else
      datain_channel_cmp <= _0226_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      datain_height_cmp <= 13'b0000000000000;
    else
      datain_height_cmp <= _0229_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      datain_width_cmp <= 13'b0000000000000;
    else
      datain_width_cmp <= _0233_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      datain_width <= 14'b00000000000000;
    else
      datain_width <= _0232_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      data_bank <= 4'b0000;
    else
      data_bank <= _0223_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      is_fp16_d1 <= 2'b00;
    else
      is_fp16_d1 <= _0388_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      is_int8_d1 <= 23'b00000000000000000000000;
    else
      is_int8_d1 <= _0390_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      is_img_d1 <= 34'b0000000000000000000000000000000000;
    else
      is_img_d1 <= _0389_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      is_winograd_d1 <= 22'b0000000000000000000000;
    else
      is_winograd_d1 <= _0391_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      layer_st_d1 <= 1'b0;
    else
      layer_st_d1 <= layer_st;
  assign _0583_ = dl_out_mask[127] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:22732" *) dl_out_data127 : sc2mac_dat_b_data127;
  assign _0582_ = dl_out_mask[126] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:22722" *) dl_out_data126 : sc2mac_dat_b_data126;
  assign _0581_ = dl_out_mask[125] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:22712" *) dl_out_data125 : sc2mac_dat_b_data125;
  assign _0580_ = dl_out_mask[124] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:22702" *) dl_out_data124 : sc2mac_dat_b_data124;
  assign _0579_ = dl_out_mask[123] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:22692" *) dl_out_data123 : sc2mac_dat_b_data123;
  assign _0578_ = dl_out_mask[122] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:22682" *) dl_out_data122 : sc2mac_dat_b_data122;
  assign _0577_ = dl_out_mask[121] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:22672" *) dl_out_data121 : sc2mac_dat_b_data121;
  assign _0576_ = dl_out_mask[120] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:22662" *) dl_out_data120 : sc2mac_dat_b_data120;
  assign _0574_ = dl_out_mask[119] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:22652" *) dl_out_data119 : sc2mac_dat_b_data119;
  assign _0573_ = dl_out_mask[118] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:22642" *) dl_out_data118 : sc2mac_dat_b_data118;
  assign _0572_ = dl_out_mask[117] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:22632" *) dl_out_data117 : sc2mac_dat_b_data117;
  assign _0571_ = dl_out_mask[116] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:22622" *) dl_out_data116 : sc2mac_dat_b_data116;
  assign _0570_ = dl_out_mask[115] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:22612" *) dl_out_data115 : sc2mac_dat_b_data115;
  assign _0569_ = dl_out_mask[114] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:22602" *) dl_out_data114 : sc2mac_dat_b_data114;
  assign _0568_ = dl_out_mask[113] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:22592" *) dl_out_data113 : sc2mac_dat_b_data113;
  assign _0567_ = dl_out_mask[112] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:22582" *) dl_out_data112 : sc2mac_dat_b_data112;
  assign _0566_ = dl_out_mask[111] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:22572" *) dl_out_data111 : sc2mac_dat_b_data111;
  assign _0565_ = dl_out_mask[110] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:22562" *) dl_out_data110 : sc2mac_dat_b_data110;
  assign _0563_ = dl_out_mask[109] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:22552" *) dl_out_data109 : sc2mac_dat_b_data109;
  assign _0562_ = dl_out_mask[108] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:22542" *) dl_out_data108 : sc2mac_dat_b_data108;
  assign _0561_ = dl_out_mask[107] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:22532" *) dl_out_data107 : sc2mac_dat_b_data107;
  assign _0560_ = dl_out_mask[106] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:22522" *) dl_out_data106 : sc2mac_dat_b_data106;
  assign _0559_ = dl_out_mask[105] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:22512" *) dl_out_data105 : sc2mac_dat_b_data105;
  assign _0558_ = dl_out_mask[104] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:22502" *) dl_out_data104 : sc2mac_dat_b_data104;
  assign _0557_ = dl_out_mask[103] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:22492" *) dl_out_data103 : sc2mac_dat_b_data103;
  assign _0556_ = dl_out_mask[102] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:22482" *) dl_out_data102 : sc2mac_dat_b_data102;
  assign _0555_ = dl_out_mask[101] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:22472" *) dl_out_data101 : sc2mac_dat_b_data101;
  assign _0554_ = dl_out_mask[100] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:22462" *) dl_out_data100 : sc2mac_dat_b_data100;
  assign _0679_ = dl_out_mask[99] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:22452" *) dl_out_data99 : sc2mac_dat_b_data99;
  assign _0678_ = dl_out_mask[98] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:22442" *) dl_out_data98 : sc2mac_dat_b_data98;
  assign _0677_ = dl_out_mask[97] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:22432" *) dl_out_data97 : sc2mac_dat_b_data97;
  assign _0676_ = dl_out_mask[96] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:22422" *) dl_out_data96 : sc2mac_dat_b_data96;
  assign _0675_ = dl_out_mask[95] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:22412" *) dl_out_data95 : sc2mac_dat_b_data95;
  assign _0674_ = dl_out_mask[94] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:22402" *) dl_out_data94 : sc2mac_dat_b_data94;
  assign _0673_ = dl_out_mask[93] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:22392" *) dl_out_data93 : sc2mac_dat_b_data93;
  assign _0672_ = dl_out_mask[92] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:22382" *) dl_out_data92 : sc2mac_dat_b_data92;
  assign _0671_ = dl_out_mask[91] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:22372" *) dl_out_data91 : sc2mac_dat_b_data91;
  assign _0670_ = dl_out_mask[90] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:22362" *) dl_out_data90 : sc2mac_dat_b_data90;
  assign _0668_ = dl_out_mask[89] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:22352" *) dl_out_data89 : sc2mac_dat_b_data89;
  assign _0667_ = dl_out_mask[88] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:22342" *) dl_out_data88 : sc2mac_dat_b_data88;
  assign _0666_ = dl_out_mask[87] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:22332" *) dl_out_data87 : sc2mac_dat_b_data87;
  assign _0665_ = dl_out_mask[86] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:22322" *) dl_out_data86 : sc2mac_dat_b_data86;
  assign _0664_ = dl_out_mask[85] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:22312" *) dl_out_data85 : sc2mac_dat_b_data85;
  assign _0663_ = dl_out_mask[84] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:22302" *) dl_out_data84 : sc2mac_dat_b_data84;
  assign _0662_ = dl_out_mask[83] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:22292" *) dl_out_data83 : sc2mac_dat_b_data83;
  assign _0661_ = dl_out_mask[82] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:22282" *) dl_out_data82 : sc2mac_dat_b_data82;
  assign _0660_ = dl_out_mask[81] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:22272" *) dl_out_data81 : sc2mac_dat_b_data81;
  assign _0659_ = dl_out_mask[80] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:22262" *) dl_out_data80 : sc2mac_dat_b_data80;
  assign _0657_ = dl_out_mask[79] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:22252" *) dl_out_data79 : sc2mac_dat_b_data79;
  assign _0656_ = dl_out_mask[78] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:22242" *) dl_out_data78 : sc2mac_dat_b_data78;
  assign _0655_ = dl_out_mask[77] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:22232" *) dl_out_data77 : sc2mac_dat_b_data77;
  assign _0654_ = dl_out_mask[76] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:22222" *) dl_out_data76 : sc2mac_dat_b_data76;
  assign _0653_ = dl_out_mask[75] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:22212" *) dl_out_data75 : sc2mac_dat_b_data75;
  assign _0652_ = dl_out_mask[74] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:22202" *) dl_out_data74 : sc2mac_dat_b_data74;
  assign _0651_ = dl_out_mask[73] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:22192" *) dl_out_data73 : sc2mac_dat_b_data73;
  assign _0650_ = dl_out_mask[72] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:22182" *) dl_out_data72 : sc2mac_dat_b_data72;
  assign _0649_ = dl_out_mask[71] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:22172" *) dl_out_data71 : sc2mac_dat_b_data71;
  assign _0648_ = dl_out_mask[70] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:22162" *) dl_out_data70 : sc2mac_dat_b_data70;
  assign _0646_ = dl_out_mask[69] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:22152" *) dl_out_data69 : sc2mac_dat_b_data69;
  assign _0645_ = dl_out_mask[68] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:22142" *) dl_out_data68 : sc2mac_dat_b_data68;
  assign _0644_ = dl_out_mask[67] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:22132" *) dl_out_data67 : sc2mac_dat_b_data67;
  assign _0643_ = dl_out_mask[66] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:22122" *) dl_out_data66 : sc2mac_dat_b_data66;
  assign _0642_ = dl_out_mask[65] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:22112" *) dl_out_data65 : sc2mac_dat_b_data65;
  assign _0641_ = dl_out_mask[64] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:22102" *) dl_out_data64 : sc2mac_dat_b_data64;
  assign _0640_ = dl_out_mask[63] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:22092" *) dl_out_data63 : sc2mac_dat_b_data63;
  assign _0639_ = dl_out_mask[62] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:22082" *) dl_out_data62 : sc2mac_dat_b_data62;
  assign _0638_ = dl_out_mask[61] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:22072" *) dl_out_data61 : sc2mac_dat_b_data61;
  assign _0637_ = dl_out_mask[60] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:22062" *) dl_out_data60 : sc2mac_dat_b_data60;
  assign _0635_ = dl_out_mask[59] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:22052" *) dl_out_data59 : sc2mac_dat_b_data59;
  assign _0634_ = dl_out_mask[58] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:22042" *) dl_out_data58 : sc2mac_dat_b_data58;
  assign _0633_ = dl_out_mask[57] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:22032" *) dl_out_data57 : sc2mac_dat_b_data57;
  assign _0632_ = dl_out_mask[56] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:22022" *) dl_out_data56 : sc2mac_dat_b_data56;
  assign _0631_ = dl_out_mask[55] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:22012" *) dl_out_data55 : sc2mac_dat_b_data55;
  assign _0630_ = dl_out_mask[54] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:22002" *) dl_out_data54 : sc2mac_dat_b_data54;
  assign _0629_ = dl_out_mask[53] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21992" *) dl_out_data53 : sc2mac_dat_b_data53;
  assign _0628_ = dl_out_mask[52] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21982" *) dl_out_data52 : sc2mac_dat_b_data52;
  assign _0627_ = dl_out_mask[51] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21972" *) dl_out_data51 : sc2mac_dat_b_data51;
  assign _0626_ = dl_out_mask[50] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21962" *) dl_out_data50 : sc2mac_dat_b_data50;
  assign _0624_ = dl_out_mask[49] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21952" *) dl_out_data49 : sc2mac_dat_b_data49;
  assign _0623_ = dl_out_mask[48] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21942" *) dl_out_data48 : sc2mac_dat_b_data48;
  assign _0622_ = dl_out_mask[47] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21932" *) dl_out_data47 : sc2mac_dat_b_data47;
  assign _0621_ = dl_out_mask[46] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21922" *) dl_out_data46 : sc2mac_dat_b_data46;
  assign _0620_ = dl_out_mask[45] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21912" *) dl_out_data45 : sc2mac_dat_b_data45;
  assign _0619_ = dl_out_mask[44] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21902" *) dl_out_data44 : sc2mac_dat_b_data44;
  assign _0618_ = dl_out_mask[43] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21892" *) dl_out_data43 : sc2mac_dat_b_data43;
  assign _0617_ = dl_out_mask[42] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21882" *) dl_out_data42 : sc2mac_dat_b_data42;
  assign _0616_ = dl_out_mask[41] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21872" *) dl_out_data41 : sc2mac_dat_b_data41;
  assign _0615_ = dl_out_mask[40] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21862" *) dl_out_data40 : sc2mac_dat_b_data40;
  assign _0613_ = dl_out_mask[39] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21852" *) dl_out_data39 : sc2mac_dat_b_data39;
  assign _0612_ = dl_out_mask[38] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21842" *) dl_out_data38 : sc2mac_dat_b_data38;
  assign _0611_ = dl_out_mask[37] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21832" *) dl_out_data37 : sc2mac_dat_b_data37;
  assign _0610_ = dl_out_mask[36] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21822" *) dl_out_data36 : sc2mac_dat_b_data36;
  assign _0609_ = dl_out_mask[35] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21812" *) dl_out_data35 : sc2mac_dat_b_data35;
  assign _0608_ = dl_out_mask[34] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21802" *) dl_out_data34 : sc2mac_dat_b_data34;
  assign _0607_ = dl_out_mask[33] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21792" *) dl_out_data33 : sc2mac_dat_b_data33;
  assign _0606_ = dl_out_mask[32] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21782" *) dl_out_data32 : sc2mac_dat_b_data32;
  assign _0605_ = dl_out_mask[31] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21772" *) dl_out_data31 : sc2mac_dat_b_data31;
  assign _0604_ = dl_out_mask[30] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21762" *) dl_out_data30 : sc2mac_dat_b_data30;
  assign _0602_ = dl_out_mask[29] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21752" *) dl_out_data29 : sc2mac_dat_b_data29;
  assign _0601_ = dl_out_mask[28] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21742" *) dl_out_data28 : sc2mac_dat_b_data28;
  assign _0600_ = dl_out_mask[27] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21732" *) dl_out_data27 : sc2mac_dat_b_data27;
  assign _0599_ = dl_out_mask[26] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21722" *) dl_out_data26 : sc2mac_dat_b_data26;
  assign _0598_ = dl_out_mask[25] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21712" *) dl_out_data25 : sc2mac_dat_b_data25;
  assign _0597_ = dl_out_mask[24] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21702" *) dl_out_data24 : sc2mac_dat_b_data24;
  assign _0596_ = dl_out_mask[23] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21692" *) dl_out_data23 : sc2mac_dat_b_data23;
  assign _0595_ = dl_out_mask[22] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21682" *) dl_out_data22 : sc2mac_dat_b_data22;
  assign _0594_ = dl_out_mask[21] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21672" *) dl_out_data21 : sc2mac_dat_b_data21;
  assign _0593_ = dl_out_mask[20] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21662" *) dl_out_data20 : sc2mac_dat_b_data20;
  assign _0591_ = dl_out_mask[19] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21652" *) dl_out_data19 : sc2mac_dat_b_data19;
  assign _0590_ = dl_out_mask[18] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21642" *) dl_out_data18 : sc2mac_dat_b_data18;
  assign _0589_ = dl_out_mask[17] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21632" *) dl_out_data17 : sc2mac_dat_b_data17;
  assign _0588_ = dl_out_mask[16] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21622" *) dl_out_data16 : sc2mac_dat_b_data16;
  assign _0587_ = dl_out_mask[15] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21612" *) dl_out_data15 : sc2mac_dat_b_data15;
  assign _0586_ = dl_out_mask[14] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21602" *) dl_out_data14 : sc2mac_dat_b_data14;
  assign _0585_ = dl_out_mask[13] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21592" *) dl_out_data13 : sc2mac_dat_b_data13;
  assign _0584_ = dl_out_mask[12] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21582" *) dl_out_data12 : sc2mac_dat_b_data12;
  assign _0575_ = dl_out_mask[11] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21572" *) dl_out_data11 : sc2mac_dat_b_data11;
  assign _0564_ = dl_out_mask[10] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21562" *) dl_out_data10 : sc2mac_dat_b_data10;
  assign _0680_ = dl_out_mask[9] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21552" *) dl_out_data9 : sc2mac_dat_b_data9;
  assign _0669_ = dl_out_mask[8] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21542" *) dl_out_data8 : sc2mac_dat_b_data8;
  assign _0658_ = dl_out_mask[7] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21532" *) dl_out_data7 : sc2mac_dat_b_data7;
  assign _0647_ = dl_out_mask[6] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21522" *) dl_out_data6 : sc2mac_dat_b_data6;
  assign _0636_ = dl_out_mask[5] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21512" *) dl_out_data5 : sc2mac_dat_b_data5;
  assign _0625_ = dl_out_mask[4] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21502" *) dl_out_data4 : sc2mac_dat_b_data4;
  assign _0614_ = dl_out_mask[3] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21492" *) dl_out_data3 : sc2mac_dat_b_data3;
  assign _0603_ = dl_out_mask[2] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21482" *) dl_out_data2 : sc2mac_dat_b_data2;
  assign _0592_ = dl_out_mask[1] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21472" *) dl_out_data1 : sc2mac_dat_b_data1;
  assign _0553_ = dl_out_mask[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21462" *) dl_out_data0 : sc2mac_dat_b_data0;
  assign _0453_ = dl_out_mask[127] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21452" *) dl_out_data127 : sc2mac_dat_a_data127;
  assign _0452_ = dl_out_mask[126] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21442" *) dl_out_data126 : sc2mac_dat_a_data126;
  assign _0451_ = dl_out_mask[125] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21432" *) dl_out_data125 : sc2mac_dat_a_data125;
  assign _0450_ = dl_out_mask[124] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21422" *) dl_out_data124 : sc2mac_dat_a_data124;
  assign _0449_ = dl_out_mask[123] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21412" *) dl_out_data123 : sc2mac_dat_a_data123;
  assign _0448_ = dl_out_mask[122] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21402" *) dl_out_data122 : sc2mac_dat_a_data122;
  assign _0447_ = dl_out_mask[121] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21392" *) dl_out_data121 : sc2mac_dat_a_data121;
  assign _0446_ = dl_out_mask[120] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21382" *) dl_out_data120 : sc2mac_dat_a_data120;
  assign _0444_ = dl_out_mask[119] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21372" *) dl_out_data119 : sc2mac_dat_a_data119;
  assign _0443_ = dl_out_mask[118] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21362" *) dl_out_data118 : sc2mac_dat_a_data118;
  assign _0442_ = dl_out_mask[117] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21352" *) dl_out_data117 : sc2mac_dat_a_data117;
  assign _0441_ = dl_out_mask[116] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21342" *) dl_out_data116 : sc2mac_dat_a_data116;
  assign _0440_ = dl_out_mask[115] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21332" *) dl_out_data115 : sc2mac_dat_a_data115;
  assign _0439_ = dl_out_mask[114] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21322" *) dl_out_data114 : sc2mac_dat_a_data114;
  assign _0438_ = dl_out_mask[113] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21312" *) dl_out_data113 : sc2mac_dat_a_data113;
  assign _0437_ = dl_out_mask[112] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21302" *) dl_out_data112 : sc2mac_dat_a_data112;
  assign _0436_ = dl_out_mask[111] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21292" *) dl_out_data111 : sc2mac_dat_a_data111;
  assign _0435_ = dl_out_mask[110] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21282" *) dl_out_data110 : sc2mac_dat_a_data110;
  assign _0433_ = dl_out_mask[109] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21272" *) dl_out_data109 : sc2mac_dat_a_data109;
  assign _0432_ = dl_out_mask[108] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21262" *) dl_out_data108 : sc2mac_dat_a_data108;
  assign _0431_ = dl_out_mask[107] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21252" *) dl_out_data107 : sc2mac_dat_a_data107;
  assign _0430_ = dl_out_mask[106] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21242" *) dl_out_data106 : sc2mac_dat_a_data106;
  assign _0429_ = dl_out_mask[105] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21232" *) dl_out_data105 : sc2mac_dat_a_data105;
  assign _0428_ = dl_out_mask[104] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21222" *) dl_out_data104 : sc2mac_dat_a_data104;
  assign _0427_ = dl_out_mask[103] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21212" *) dl_out_data103 : sc2mac_dat_a_data103;
  assign _0426_ = dl_out_mask[102] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21202" *) dl_out_data102 : sc2mac_dat_a_data102;
  assign _0425_ = dl_out_mask[101] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21192" *) dl_out_data101 : sc2mac_dat_a_data101;
  assign _0424_ = dl_out_mask[100] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21182" *) dl_out_data100 : sc2mac_dat_a_data100;
  assign _0549_ = dl_out_mask[99] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21172" *) dl_out_data99 : sc2mac_dat_a_data99;
  assign _0548_ = dl_out_mask[98] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21162" *) dl_out_data98 : sc2mac_dat_a_data98;
  assign _0547_ = dl_out_mask[97] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21152" *) dl_out_data97 : sc2mac_dat_a_data97;
  assign _0546_ = dl_out_mask[96] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21142" *) dl_out_data96 : sc2mac_dat_a_data96;
  assign _0545_ = dl_out_mask[95] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21132" *) dl_out_data95 : sc2mac_dat_a_data95;
  assign _0544_ = dl_out_mask[94] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21122" *) dl_out_data94 : sc2mac_dat_a_data94;
  assign _0543_ = dl_out_mask[93] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21112" *) dl_out_data93 : sc2mac_dat_a_data93;
  assign _0542_ = dl_out_mask[92] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21102" *) dl_out_data92 : sc2mac_dat_a_data92;
  assign _0541_ = dl_out_mask[91] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21092" *) dl_out_data91 : sc2mac_dat_a_data91;
  assign _0540_ = dl_out_mask[90] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21082" *) dl_out_data90 : sc2mac_dat_a_data90;
  assign _0538_ = dl_out_mask[89] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21072" *) dl_out_data89 : sc2mac_dat_a_data89;
  assign _0537_ = dl_out_mask[88] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21062" *) dl_out_data88 : sc2mac_dat_a_data88;
  assign _0536_ = dl_out_mask[87] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21052" *) dl_out_data87 : sc2mac_dat_a_data87;
  assign _0535_ = dl_out_mask[86] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21042" *) dl_out_data86 : sc2mac_dat_a_data86;
  assign _0534_ = dl_out_mask[85] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21032" *) dl_out_data85 : sc2mac_dat_a_data85;
  assign _0533_ = dl_out_mask[84] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21022" *) dl_out_data84 : sc2mac_dat_a_data84;
  assign _0532_ = dl_out_mask[83] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21012" *) dl_out_data83 : sc2mac_dat_a_data83;
  assign _0531_ = dl_out_mask[82] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:21002" *) dl_out_data82 : sc2mac_dat_a_data82;
  assign _0530_ = dl_out_mask[81] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:20992" *) dl_out_data81 : sc2mac_dat_a_data81;
  assign _0529_ = dl_out_mask[80] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:20982" *) dl_out_data80 : sc2mac_dat_a_data80;
  assign _0527_ = dl_out_mask[79] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:20972" *) dl_out_data79 : sc2mac_dat_a_data79;
  assign _0526_ = dl_out_mask[78] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:20962" *) dl_out_data78 : sc2mac_dat_a_data78;
  assign _0525_ = dl_out_mask[77] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:20952" *) dl_out_data77 : sc2mac_dat_a_data77;
  assign _0524_ = dl_out_mask[76] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:20942" *) dl_out_data76 : sc2mac_dat_a_data76;
  assign _0523_ = dl_out_mask[75] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:20932" *) dl_out_data75 : sc2mac_dat_a_data75;
  assign _0522_ = dl_out_mask[74] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:20922" *) dl_out_data74 : sc2mac_dat_a_data74;
  assign _0521_ = dl_out_mask[73] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:20912" *) dl_out_data73 : sc2mac_dat_a_data73;
  assign _0520_ = dl_out_mask[72] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:20902" *) dl_out_data72 : sc2mac_dat_a_data72;
  assign _0519_ = dl_out_mask[71] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:20892" *) dl_out_data71 : sc2mac_dat_a_data71;
  assign _0518_ = dl_out_mask[70] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:20882" *) dl_out_data70 : sc2mac_dat_a_data70;
  assign _0516_ = dl_out_mask[69] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:20872" *) dl_out_data69 : sc2mac_dat_a_data69;
  assign _0515_ = dl_out_mask[68] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:20862" *) dl_out_data68 : sc2mac_dat_a_data68;
  assign _0514_ = dl_out_mask[67] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:20852" *) dl_out_data67 : sc2mac_dat_a_data67;
  assign _0513_ = dl_out_mask[66] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:20842" *) dl_out_data66 : sc2mac_dat_a_data66;
  assign _0512_ = dl_out_mask[65] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:20832" *) dl_out_data65 : sc2mac_dat_a_data65;
  assign _0511_ = dl_out_mask[64] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:20822" *) dl_out_data64 : sc2mac_dat_a_data64;
  assign _0510_ = dl_out_mask[63] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:20812" *) dl_out_data63 : sc2mac_dat_a_data63;
  assign _0509_ = dl_out_mask[62] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:20802" *) dl_out_data62 : sc2mac_dat_a_data62;
  assign _0508_ = dl_out_mask[61] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:20792" *) dl_out_data61 : sc2mac_dat_a_data61;
  assign _0507_ = dl_out_mask[60] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:20782" *) dl_out_data60 : sc2mac_dat_a_data60;
  assign _0505_ = dl_out_mask[59] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:20772" *) dl_out_data59 : sc2mac_dat_a_data59;
  assign _0504_ = dl_out_mask[58] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:20762" *) dl_out_data58 : sc2mac_dat_a_data58;
  assign _0503_ = dl_out_mask[57] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:20752" *) dl_out_data57 : sc2mac_dat_a_data57;
  assign _0502_ = dl_out_mask[56] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:20742" *) dl_out_data56 : sc2mac_dat_a_data56;
  assign _0501_ = dl_out_mask[55] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:20732" *) dl_out_data55 : sc2mac_dat_a_data55;
  assign _0500_ = dl_out_mask[54] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:20722" *) dl_out_data54 : sc2mac_dat_a_data54;
  assign _0499_ = dl_out_mask[53] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:20712" *) dl_out_data53 : sc2mac_dat_a_data53;
  assign _0498_ = dl_out_mask[52] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:20702" *) dl_out_data52 : sc2mac_dat_a_data52;
  assign _0497_ = dl_out_mask[51] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:20692" *) dl_out_data51 : sc2mac_dat_a_data51;
  assign _0496_ = dl_out_mask[50] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:20682" *) dl_out_data50 : sc2mac_dat_a_data50;
  assign _0494_ = dl_out_mask[49] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:20672" *) dl_out_data49 : sc2mac_dat_a_data49;
  assign _0493_ = dl_out_mask[48] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:20662" *) dl_out_data48 : sc2mac_dat_a_data48;
  assign _0492_ = dl_out_mask[47] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:20652" *) dl_out_data47 : sc2mac_dat_a_data47;
  assign _0491_ = dl_out_mask[46] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:20642" *) dl_out_data46 : sc2mac_dat_a_data46;
  assign _0490_ = dl_out_mask[45] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:20632" *) dl_out_data45 : sc2mac_dat_a_data45;
  assign _0489_ = dl_out_mask[44] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:20622" *) dl_out_data44 : sc2mac_dat_a_data44;
  assign _0488_ = dl_out_mask[43] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:20612" *) dl_out_data43 : sc2mac_dat_a_data43;
  assign _0487_ = dl_out_mask[42] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:20602" *) dl_out_data42 : sc2mac_dat_a_data42;
  assign _0486_ = dl_out_mask[41] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:20592" *) dl_out_data41 : sc2mac_dat_a_data41;
  assign _0485_ = dl_out_mask[40] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:20582" *) dl_out_data40 : sc2mac_dat_a_data40;
  assign _0483_ = dl_out_mask[39] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:20572" *) dl_out_data39 : sc2mac_dat_a_data39;
  assign _0482_ = dl_out_mask[38] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:20562" *) dl_out_data38 : sc2mac_dat_a_data38;
  assign _0481_ = dl_out_mask[37] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:20552" *) dl_out_data37 : sc2mac_dat_a_data37;
  assign _0480_ = dl_out_mask[36] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:20542" *) dl_out_data36 : sc2mac_dat_a_data36;
  assign _0479_ = dl_out_mask[35] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:20532" *) dl_out_data35 : sc2mac_dat_a_data35;
  assign _0478_ = dl_out_mask[34] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:20522" *) dl_out_data34 : sc2mac_dat_a_data34;
  assign _0477_ = dl_out_mask[33] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:20512" *) dl_out_data33 : sc2mac_dat_a_data33;
  assign _0476_ = dl_out_mask[32] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:20502" *) dl_out_data32 : sc2mac_dat_a_data32;
  assign _0475_ = dl_out_mask[31] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:20492" *) dl_out_data31 : sc2mac_dat_a_data31;
  assign _0474_ = dl_out_mask[30] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:20482" *) dl_out_data30 : sc2mac_dat_a_data30;
  assign _0472_ = dl_out_mask[29] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:20472" *) dl_out_data29 : sc2mac_dat_a_data29;
  assign _0471_ = dl_out_mask[28] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:20462" *) dl_out_data28 : sc2mac_dat_a_data28;
  assign _0470_ = dl_out_mask[27] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:20452" *) dl_out_data27 : sc2mac_dat_a_data27;
  assign _0469_ = dl_out_mask[26] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:20442" *) dl_out_data26 : sc2mac_dat_a_data26;
  assign _0468_ = dl_out_mask[25] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:20432" *) dl_out_data25 : sc2mac_dat_a_data25;
  assign _0467_ = dl_out_mask[24] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:20422" *) dl_out_data24 : sc2mac_dat_a_data24;
  assign _0466_ = dl_out_mask[23] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:20412" *) dl_out_data23 : sc2mac_dat_a_data23;
  assign _0465_ = dl_out_mask[22] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:20402" *) dl_out_data22 : sc2mac_dat_a_data22;
  assign _0464_ = dl_out_mask[21] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:20392" *) dl_out_data21 : sc2mac_dat_a_data21;
  assign _0463_ = dl_out_mask[20] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:20382" *) dl_out_data20 : sc2mac_dat_a_data20;
  assign _0461_ = dl_out_mask[19] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:20372" *) dl_out_data19 : sc2mac_dat_a_data19;
  assign _0460_ = dl_out_mask[18] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:20362" *) dl_out_data18 : sc2mac_dat_a_data18;
  assign _0459_ = dl_out_mask[17] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:20352" *) dl_out_data17 : sc2mac_dat_a_data17;
  assign _0458_ = dl_out_mask[16] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:20342" *) dl_out_data16 : sc2mac_dat_a_data16;
  assign _0457_ = dl_out_mask[15] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:20332" *) dl_out_data15 : sc2mac_dat_a_data15;
  assign _0456_ = dl_out_mask[14] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:20322" *) dl_out_data14 : sc2mac_dat_a_data14;
  assign _0455_ = dl_out_mask[13] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:20312" *) dl_out_data13 : sc2mac_dat_a_data13;
  assign _0454_ = dl_out_mask[12] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:20302" *) dl_out_data12 : sc2mac_dat_a_data12;
  assign _0445_ = dl_out_mask[11] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:20292" *) dl_out_data11 : sc2mac_dat_a_data11;
  assign _0434_ = dl_out_mask[10] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:20282" *) dl_out_data10 : sc2mac_dat_a_data10;
  assign _0550_ = dl_out_mask[9] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:20272" *) dl_out_data9 : sc2mac_dat_a_data9;
  assign _0539_ = dl_out_mask[8] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:20262" *) dl_out_data8 : sc2mac_dat_a_data8;
  assign _0528_ = dl_out_mask[7] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:20252" *) dl_out_data7 : sc2mac_dat_a_data7;
  assign _0517_ = dl_out_mask[6] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:20242" *) dl_out_data6 : sc2mac_dat_a_data6;
  assign _0506_ = dl_out_mask[5] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:20232" *) dl_out_data5 : sc2mac_dat_a_data5;
  assign _0495_ = dl_out_mask[4] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:20222" *) dl_out_data4 : sc2mac_dat_a_data4;
  assign _0484_ = dl_out_mask[3] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:20212" *) dl_out_data3 : sc2mac_dat_a_data3;
  assign _0473_ = dl_out_mask[2] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:20202" *) dl_out_data2 : sc2mac_dat_a_data2;
  assign _0462_ = dl_out_mask[1] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:20192" *) dl_out_data1 : sc2mac_dat_a_data1;
  assign _0423_ = dl_out_mask[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:20182" *) dl_out_data0 : sc2mac_dat_a_data0;
  assign _0681_ = _1054_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:20124" *) dl_out_mask : sc2mac_dat_b_mask;
  assign _0551_ = _1054_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:20063" *) dl_out_mask : sc2mac_dat_a_mask;
  assign _0682_ = _1054_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:20002" *) sc2mac_dat_pd_w : sc2mac_dat_b_pd;
  assign _0552_ = _1054_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:19941" *) sc2mac_dat_pd_w : sc2mac_dat_a_pd;
  assign _0272_ = dat_out_mask[127] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:19898" *) dat_out_data[1023:1016] : dl_out_data127;
  assign _0271_ = dat_out_mask[126] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:19888" *) dat_out_data[1015:1008] : dl_out_data126;
  assign _0270_ = dat_out_mask[125] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:19878" *) dat_out_data[1007:1000] : dl_out_data125;
  assign _0269_ = dat_out_mask[124] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:19868" *) dat_out_data[999:992] : dl_out_data124;
  assign _0268_ = dat_out_mask[123] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:19858" *) dat_out_data[991:984] : dl_out_data123;
  assign _0267_ = dat_out_mask[122] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:19848" *) dat_out_data[983:976] : dl_out_data122;
  assign _0266_ = dat_out_mask[121] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:19838" *) dat_out_data[975:968] : dl_out_data121;
  assign _0265_ = dat_out_mask[120] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:19828" *) dat_out_data[967:960] : dl_out_data120;
  assign _0263_ = dat_out_mask[119] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:19818" *) dat_out_data[959:952] : dl_out_data119;
  assign _0262_ = dat_out_mask[118] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:19808" *) dat_out_data[951:944] : dl_out_data118;
  assign _0261_ = dat_out_mask[117] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:19798" *) dat_out_data[943:936] : dl_out_data117;
  assign _0260_ = dat_out_mask[116] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:19788" *) dat_out_data[935:928] : dl_out_data116;
  assign _0259_ = dat_out_mask[115] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:19778" *) dat_out_data[927:920] : dl_out_data115;
  assign _0258_ = dat_out_mask[114] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:19768" *) dat_out_data[919:912] : dl_out_data114;
  assign _0257_ = dat_out_mask[113] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:19758" *) dat_out_data[911:904] : dl_out_data113;
  assign _0256_ = dat_out_mask[112] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:19748" *) dat_out_data[903:896] : dl_out_data112;
  assign _0255_ = dat_out_mask[111] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:19738" *) dat_out_data[895:888] : dl_out_data111;
  assign _0254_ = dat_out_mask[110] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:19728" *) dat_out_data[887:880] : dl_out_data110;
  assign _0252_ = dat_out_mask[109] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:19718" *) dat_out_data[879:872] : dl_out_data109;
  assign _0251_ = dat_out_mask[108] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:19708" *) dat_out_data[871:864] : dl_out_data108;
  assign _0250_ = dat_out_mask[107] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:19698" *) dat_out_data[863:856] : dl_out_data107;
  assign _0249_ = dat_out_mask[106] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:19688" *) dat_out_data[855:848] : dl_out_data106;
  assign _0248_ = dat_out_mask[105] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:19678" *) dat_out_data[847:840] : dl_out_data105;
  assign _0247_ = dat_out_mask[104] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:19668" *) dat_out_data[839:832] : dl_out_data104;
  assign _0246_ = dat_out_mask[103] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:19658" *) dat_out_data[831:824] : dl_out_data103;
  assign _0245_ = dat_out_mask[102] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:19648" *) dat_out_data[823:816] : dl_out_data102;
  assign _0244_ = dat_out_mask[101] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:19638" *) dat_out_data[815:808] : dl_out_data101;
  assign _0243_ = dat_out_mask[100] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:19628" *) dat_out_data[807:800] : dl_out_data100;
  assign _0368_ = dat_out_mask[99] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:19618" *) dat_out_data[799:792] : dl_out_data99;
  assign _0367_ = dat_out_mask[98] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:19608" *) dat_out_data[791:784] : dl_out_data98;
  assign _0366_ = dat_out_mask[97] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:19598" *) dat_out_data[783:776] : dl_out_data97;
  assign _0365_ = dat_out_mask[96] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:19588" *) dat_out_data[775:768] : dl_out_data96;
  assign _0364_ = dat_out_mask[95] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:19578" *) dat_out_data[767:760] : dl_out_data95;
  assign _0363_ = dat_out_mask[94] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:19568" *) dat_out_data[759:752] : dl_out_data94;
  assign _0362_ = dat_out_mask[93] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:19558" *) dat_out_data[751:744] : dl_out_data93;
  assign _0361_ = dat_out_mask[92] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:19548" *) dat_out_data[743:736] : dl_out_data92;
  assign _0360_ = dat_out_mask[91] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:19538" *) dat_out_data[735:728] : dl_out_data91;
  assign _0359_ = dat_out_mask[90] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:19528" *) dat_out_data[727:720] : dl_out_data90;
  assign _0357_ = dat_out_mask[89] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:19518" *) dat_out_data[719:712] : dl_out_data89;
  assign _0356_ = dat_out_mask[88] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:19508" *) dat_out_data[711:704] : dl_out_data88;
  assign _0355_ = dat_out_mask[87] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:19498" *) dat_out_data[703:696] : dl_out_data87;
  assign _0354_ = dat_out_mask[86] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:19488" *) dat_out_data[695:688] : dl_out_data86;
  assign _0353_ = dat_out_mask[85] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:19478" *) dat_out_data[687:680] : dl_out_data85;
  assign _0352_ = dat_out_mask[84] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:19468" *) dat_out_data[679:672] : dl_out_data84;
  assign _0351_ = dat_out_mask[83] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:19458" *) dat_out_data[671:664] : dl_out_data83;
  assign _0350_ = dat_out_mask[82] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:19448" *) dat_out_data[663:656] : dl_out_data82;
  assign _0349_ = dat_out_mask[81] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:19438" *) dat_out_data[655:648] : dl_out_data81;
  assign _0348_ = dat_out_mask[80] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:19428" *) dat_out_data[647:640] : dl_out_data80;
  assign _0346_ = dat_out_mask[79] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:19418" *) dat_out_data[639:632] : dl_out_data79;
  assign _0345_ = dat_out_mask[78] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:19408" *) dat_out_data[631:624] : dl_out_data78;
  assign _0344_ = dat_out_mask[77] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:19398" *) dat_out_data[623:616] : dl_out_data77;
  assign _0343_ = dat_out_mask[76] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:19388" *) dat_out_data[615:608] : dl_out_data76;
  assign _0342_ = dat_out_mask[75] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:19378" *) dat_out_data[607:600] : dl_out_data75;
  assign _0341_ = dat_out_mask[74] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:19368" *) dat_out_data[599:592] : dl_out_data74;
  assign _0340_ = dat_out_mask[73] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:19358" *) dat_out_data[591:584] : dl_out_data73;
  assign _0339_ = dat_out_mask[72] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:19348" *) dat_out_data[583:576] : dl_out_data72;
  assign _0338_ = dat_out_mask[71] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:19338" *) dat_out_data[575:568] : dl_out_data71;
  assign _0337_ = dat_out_mask[70] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:19328" *) dat_out_data[567:560] : dl_out_data70;
  assign _0335_ = dat_out_mask[69] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:19318" *) dat_out_data[559:552] : dl_out_data69;
  assign _0334_ = dat_out_mask[68] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:19308" *) dat_out_data[551:544] : dl_out_data68;
  assign _0333_ = dat_out_mask[67] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:19298" *) dat_out_data[543:536] : dl_out_data67;
  assign _0332_ = dat_out_mask[66] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:19288" *) dat_out_data[535:528] : dl_out_data66;
  assign _0331_ = dat_out_mask[65] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:19278" *) dat_out_data[527:520] : dl_out_data65;
  assign _0330_ = dat_out_mask[64] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:19268" *) dat_out_data[519:512] : dl_out_data64;
  assign _0329_ = dat_out_mask[63] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:19258" *) dat_out_data[511:504] : dl_out_data63;
  assign _0328_ = dat_out_mask[62] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:19248" *) dat_out_data[503:496] : dl_out_data62;
  assign _0327_ = dat_out_mask[61] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:19238" *) dat_out_data[495:488] : dl_out_data61;
  assign _0326_ = dat_out_mask[60] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:19228" *) dat_out_data[487:480] : dl_out_data60;
  assign _0324_ = dat_out_mask[59] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:19218" *) dat_out_data[479:472] : dl_out_data59;
  assign _0323_ = dat_out_mask[58] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:19208" *) dat_out_data[471:464] : dl_out_data58;
  assign _0322_ = dat_out_mask[57] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:19198" *) dat_out_data[463:456] : dl_out_data57;
  assign _0321_ = dat_out_mask[56] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:19188" *) dat_out_data[455:448] : dl_out_data56;
  assign _0320_ = dat_out_mask[55] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:19178" *) dat_out_data[447:440] : dl_out_data55;
  assign _0319_ = dat_out_mask[54] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:19168" *) dat_out_data[439:432] : dl_out_data54;
  assign _0318_ = dat_out_mask[53] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:19158" *) dat_out_data[431:424] : dl_out_data53;
  assign _0317_ = dat_out_mask[52] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:19148" *) dat_out_data[423:416] : dl_out_data52;
  assign _0316_ = dat_out_mask[51] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:19138" *) dat_out_data[415:408] : dl_out_data51;
  assign _0315_ = dat_out_mask[50] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:19128" *) dat_out_data[407:400] : dl_out_data50;
  assign _0313_ = dat_out_mask[49] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:19118" *) dat_out_data[399:392] : dl_out_data49;
  assign _0312_ = dat_out_mask[48] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:19108" *) dat_out_data[391:384] : dl_out_data48;
  assign _0311_ = dat_out_mask[47] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:19098" *) dat_out_data[383:376] : dl_out_data47;
  assign _0310_ = dat_out_mask[46] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:19088" *) dat_out_data[375:368] : dl_out_data46;
  assign _0309_ = dat_out_mask[45] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:19078" *) dat_out_data[367:360] : dl_out_data45;
  assign _0308_ = dat_out_mask[44] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:19068" *) dat_out_data[359:352] : dl_out_data44;
  assign _0307_ = dat_out_mask[43] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:19058" *) dat_out_data[351:344] : dl_out_data43;
  assign _0306_ = dat_out_mask[42] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:19048" *) dat_out_data[343:336] : dl_out_data42;
  assign _0305_ = dat_out_mask[41] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:19038" *) dat_out_data[335:328] : dl_out_data41;
  assign _0304_ = dat_out_mask[40] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:19028" *) dat_out_data[327:320] : dl_out_data40;
  assign _0302_ = dat_out_mask[39] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:19018" *) dat_out_data[319:312] : dl_out_data39;
  assign _0301_ = dat_out_mask[38] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:19008" *) dat_out_data[311:304] : dl_out_data38;
  assign _0300_ = dat_out_mask[37] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18998" *) dat_out_data[303:296] : dl_out_data37;
  assign _0299_ = dat_out_mask[36] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18988" *) dat_out_data[295:288] : dl_out_data36;
  assign _0298_ = dat_out_mask[35] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18978" *) dat_out_data[287:280] : dl_out_data35;
  assign _0297_ = dat_out_mask[34] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18968" *) dat_out_data[279:272] : dl_out_data34;
  assign _0296_ = dat_out_mask[33] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18958" *) dat_out_data[271:264] : dl_out_data33;
  assign _0295_ = dat_out_mask[32] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18948" *) dat_out_data[263:256] : dl_out_data32;
  assign _0294_ = dat_out_mask[31] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18938" *) dat_out_data[255:248] : dl_out_data31;
  assign _0293_ = dat_out_mask[30] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18928" *) dat_out_data[247:240] : dl_out_data30;
  assign _0291_ = dat_out_mask[29] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18918" *) dat_out_data[239:232] : dl_out_data29;
  assign _0290_ = dat_out_mask[28] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18908" *) dat_out_data[231:224] : dl_out_data28;
  assign _0289_ = dat_out_mask[27] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18898" *) dat_out_data[223:216] : dl_out_data27;
  assign _0288_ = dat_out_mask[26] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18888" *) dat_out_data[215:208] : dl_out_data26;
  assign _0287_ = dat_out_mask[25] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18878" *) dat_out_data[207:200] : dl_out_data25;
  assign _0286_ = dat_out_mask[24] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18868" *) dat_out_data[199:192] : dl_out_data24;
  assign _0285_ = dat_out_mask[23] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18858" *) dat_out_data[191:184] : dl_out_data23;
  assign _0284_ = dat_out_mask[22] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18848" *) dat_out_data[183:176] : dl_out_data22;
  assign _0283_ = dat_out_mask[21] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18838" *) dat_out_data[175:168] : dl_out_data21;
  assign _0282_ = dat_out_mask[20] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18828" *) dat_out_data[167:160] : dl_out_data20;
  assign _0280_ = dat_out_mask[19] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18818" *) dat_out_data[159:152] : dl_out_data19;
  assign _0279_ = dat_out_mask[18] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18808" *) dat_out_data[151:144] : dl_out_data18;
  assign _0278_ = dat_out_mask[17] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18798" *) dat_out_data[143:136] : dl_out_data17;
  assign _0277_ = dat_out_mask[16] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18788" *) dat_out_data[135:128] : dl_out_data16;
  assign _0276_ = dat_out_mask[15] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18778" *) dat_out_data[127:120] : dl_out_data15;
  assign _0275_ = dat_out_mask[14] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18768" *) dat_out_data[119:112] : dl_out_data14;
  assign _0274_ = dat_out_mask[13] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18758" *) dat_out_data[111:104] : dl_out_data13;
  assign _0273_ = dat_out_mask[12] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18748" *) dat_out_data[103:96] : dl_out_data12;
  assign _0264_ = dat_out_mask[11] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18738" *) dat_out_data[95:88] : dl_out_data11;
  assign _0253_ = dat_out_mask[10] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18728" *) dat_out_data[87:80] : dl_out_data10;
  assign _0369_ = dat_out_mask[9] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18718" *) dat_out_data[79:72] : dl_out_data9;
  assign _0358_ = dat_out_mask[8] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18708" *) dat_out_data[71:64] : dl_out_data8;
  assign _0347_ = dat_out_mask[7] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18698" *) dat_out_data[63:56] : dl_out_data7;
  assign _0336_ = dat_out_mask[6] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18688" *) dat_out_data[55:48] : dl_out_data6;
  assign _0325_ = dat_out_mask[5] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18678" *) dat_out_data[47:40] : dl_out_data5;
  assign _0314_ = dat_out_mask[4] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18668" *) dat_out_data[39:32] : dl_out_data4;
  assign _0303_ = dat_out_mask[3] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18658" *) dat_out_data[31:24] : dl_out_data3;
  assign _0292_ = dat_out_mask[2] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18648" *) dat_out_data[23:16] : dl_out_data2;
  assign _0281_ = dat_out_mask[1] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18638" *) dat_out_data[15:8] : dl_out_data1;
  assign _0242_ = dat_out_mask[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18628" *) dat_out_data[7:0] : dl_out_data0;
  assign _0370_ = dat_out_pvld ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18570" *) dat_out_flag : dl_out_flag;
  assign _0371_ = _1053_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18509" *) dat_out_mask : dl_out_mask;
  assign _0222_ = dat_rsp_pra_en ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18251" *) dat_rsp_wg_ch3 : dat_rsp_wg_ch3_d1;
  assign _0221_ = dat_rsp_pra_en ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18241" *) dat_rsp_wg_ch2 : dat_rsp_wg_ch2_d1;
  assign _0220_ = dat_rsp_pra_en ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18231" *) dat_rsp_wg_ch1 : dat_rsp_wg_ch1_d1;
  assign _0219_ = dat_rsp_pra_en ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18221" *) dat_rsp_wg_ch0 : dat_rsp_wg_ch0_d1;
  assign _0025_ = _0974_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18193" *) dat_out_bypass_data_w[1023:1016] : dat_out_bypass_data[1023:1016];
  assign _0024_ = _0973_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18183" *) dat_out_bypass_data_w[1015:1008] : dat_out_bypass_data[1015:1008];
  assign _0023_ = _0972_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18173" *) dat_out_bypass_data_w[1007:1000] : dat_out_bypass_data[1007:1000];
  assign _0150_ = _0971_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18163" *) dat_out_bypass_data_w[999:992] : dat_out_bypass_data[999:992];
  assign _0149_ = _0970_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18153" *) dat_out_bypass_data_w[991:984] : dat_out_bypass_data[991:984];
  assign _0148_ = _0969_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18143" *) dat_out_bypass_data_w[983:976] : dat_out_bypass_data[983:976];
  assign _0147_ = _0968_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18133" *) dat_out_bypass_data_w[975:968] : dat_out_bypass_data[975:968];
  assign _0146_ = _0967_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18123" *) dat_out_bypass_data_w[967:960] : dat_out_bypass_data[967:960];
  assign _0144_ = _0966_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18113" *) dat_out_bypass_data_w[959:952] : dat_out_bypass_data[959:952];
  assign _0143_ = _0965_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18103" *) dat_out_bypass_data_w[951:944] : dat_out_bypass_data[951:944];
  assign _0142_ = _0964_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18093" *) dat_out_bypass_data_w[943:936] : dat_out_bypass_data[943:936];
  assign _0141_ = _0963_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18083" *) dat_out_bypass_data_w[935:928] : dat_out_bypass_data[935:928];
  assign _0140_ = _0962_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18073" *) dat_out_bypass_data_w[927:920] : dat_out_bypass_data[927:920];
  assign _0139_ = _0961_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18063" *) dat_out_bypass_data_w[919:912] : dat_out_bypass_data[919:912];
  assign _0138_ = _0960_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18053" *) dat_out_bypass_data_w[911:904] : dat_out_bypass_data[911:904];
  assign _0137_ = _0959_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18043" *) dat_out_bypass_data_w[903:896] : dat_out_bypass_data[903:896];
  assign _0136_ = _0958_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18033" *) dat_out_bypass_data_w[895:888] : dat_out_bypass_data[895:888];
  assign _0135_ = _0957_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18023" *) dat_out_bypass_data_w[887:880] : dat_out_bypass_data[887:880];
  assign _0133_ = _0956_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18013" *) dat_out_bypass_data_w[879:872] : dat_out_bypass_data[879:872];
  assign _0132_ = _0955_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18003" *) dat_out_bypass_data_w[871:864] : dat_out_bypass_data[871:864];
  assign _0131_ = _0954_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17993" *) dat_out_bypass_data_w[863:856] : dat_out_bypass_data[863:856];
  assign _0130_ = _0953_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17983" *) dat_out_bypass_data_w[855:848] : dat_out_bypass_data[855:848];
  assign _0129_ = _0952_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17973" *) dat_out_bypass_data_w[847:840] : dat_out_bypass_data[847:840];
  assign _0128_ = _0951_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17963" *) dat_out_bypass_data_w[839:832] : dat_out_bypass_data[839:832];
  assign _0127_ = _0950_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17953" *) dat_out_bypass_data_w[831:824] : dat_out_bypass_data[831:824];
  assign _0126_ = _0949_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17943" *) dat_out_bypass_data_w[823:816] : dat_out_bypass_data[823:816];
  assign _0125_ = _0948_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17933" *) dat_out_bypass_data_w[815:808] : dat_out_bypass_data[815:808];
  assign _0124_ = _0947_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17923" *) dat_out_bypass_data_w[807:800] : dat_out_bypass_data[807:800];
  assign _0121_ = _0946_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17913" *) dat_out_bypass_data_w[799:792] : dat_out_bypass_data[799:792];
  assign _0120_ = _0945_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17903" *) dat_out_bypass_data_w[791:784] : dat_out_bypass_data[791:784];
  assign _0119_ = _0944_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17893" *) dat_out_bypass_data_w[783:776] : dat_out_bypass_data[783:776];
  assign _0118_ = _0943_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17883" *) dat_out_bypass_data_w[775:768] : dat_out_bypass_data[775:768];
  assign _0117_ = _0942_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17873" *) dat_out_bypass_data_w[767:760] : dat_out_bypass_data[767:760];
  assign _0116_ = _0941_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17863" *) dat_out_bypass_data_w[759:752] : dat_out_bypass_data[759:752];
  assign _0115_ = _0940_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17853" *) dat_out_bypass_data_w[751:744] : dat_out_bypass_data[751:744];
  assign _0114_ = _0939_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17843" *) dat_out_bypass_data_w[743:736] : dat_out_bypass_data[743:736];
  assign _0113_ = _0938_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17833" *) dat_out_bypass_data_w[735:728] : dat_out_bypass_data[735:728];
  assign _0112_ = _0937_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17823" *) dat_out_bypass_data_w[727:720] : dat_out_bypass_data[727:720];
  assign _0110_ = _0936_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17813" *) dat_out_bypass_data_w[719:712] : dat_out_bypass_data[719:712];
  assign _0109_ = _0935_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17803" *) dat_out_bypass_data_w[711:704] : dat_out_bypass_data[711:704];
  assign _0108_ = _0934_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17793" *) dat_out_bypass_data_w[703:696] : dat_out_bypass_data[703:696];
  assign _0107_ = _0933_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17783" *) dat_out_bypass_data_w[695:688] : dat_out_bypass_data[695:688];
  assign _0106_ = _0932_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17773" *) dat_out_bypass_data_w[687:680] : dat_out_bypass_data[687:680];
  assign _0105_ = _0931_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17763" *) dat_out_bypass_data_w[679:672] : dat_out_bypass_data[679:672];
  assign _0104_ = _0930_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17753" *) dat_out_bypass_data_w[671:664] : dat_out_bypass_data[671:664];
  assign _0103_ = _0929_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17743" *) dat_out_bypass_data_w[663:656] : dat_out_bypass_data[663:656];
  assign _0102_ = _0928_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17733" *) dat_out_bypass_data_w[655:648] : dat_out_bypass_data[655:648];
  assign _0101_ = _0927_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17723" *) dat_out_bypass_data_w[647:640] : dat_out_bypass_data[647:640];
  assign _0099_ = _0926_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17713" *) dat_out_bypass_data_w[639:632] : dat_out_bypass_data[639:632];
  assign _0098_ = _0925_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17703" *) dat_out_bypass_data_w[631:624] : dat_out_bypass_data[631:624];
  assign _0097_ = _0924_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17693" *) dat_out_bypass_data_w[623:616] : dat_out_bypass_data[623:616];
  assign _0096_ = _0923_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17683" *) dat_out_bypass_data_w[615:608] : dat_out_bypass_data[615:608];
  assign _0095_ = _0922_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17673" *) dat_out_bypass_data_w[607:600] : dat_out_bypass_data[607:600];
  assign _0094_ = _0921_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17663" *) dat_out_bypass_data_w[599:592] : dat_out_bypass_data[599:592];
  assign _0093_ = _0920_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17653" *) dat_out_bypass_data_w[591:584] : dat_out_bypass_data[591:584];
  assign _0092_ = _0919_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17643" *) dat_out_bypass_data_w[583:576] : dat_out_bypass_data[583:576];
  assign _0091_ = _0918_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17633" *) dat_out_bypass_data_w[575:568] : dat_out_bypass_data[575:568];
  assign _0090_ = _0917_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17623" *) dat_out_bypass_data_w[567:560] : dat_out_bypass_data[567:560];
  assign _0088_ = _0916_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17613" *) dat_out_bypass_data_w[559:552] : dat_out_bypass_data[559:552];
  assign _0087_ = _0915_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17603" *) dat_out_bypass_data_w[551:544] : dat_out_bypass_data[551:544];
  assign _0086_ = _0914_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17593" *) dat_out_bypass_data_w[543:536] : dat_out_bypass_data[543:536];
  assign _0085_ = _0913_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17583" *) dat_out_bypass_data_w[535:528] : dat_out_bypass_data[535:528];
  assign _0084_ = _0912_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17573" *) dat_out_bypass_data_w[527:520] : dat_out_bypass_data[527:520];
  assign _0083_ = _0911_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17563" *) dat_out_bypass_data_w[519:512] : dat_out_bypass_data[519:512];
  assign _0082_ = _0910_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17553" *) dat_out_bypass_data_w[511:504] : dat_out_bypass_data[511:504];
  assign _0081_ = _0909_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17543" *) dat_out_bypass_data_w[503:496] : dat_out_bypass_data[503:496];
  assign _0080_ = _0908_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17533" *) dat_out_bypass_data_w[495:488] : dat_out_bypass_data[495:488];
  assign _0079_ = _0907_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17523" *) dat_out_bypass_data_w[487:480] : dat_out_bypass_data[487:480];
  assign _0077_ = _0906_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17513" *) dat_out_bypass_data_w[479:472] : dat_out_bypass_data[479:472];
  assign _0076_ = _0905_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17503" *) dat_out_bypass_data_w[471:464] : dat_out_bypass_data[471:464];
  assign _0075_ = _0904_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17493" *) dat_out_bypass_data_w[463:456] : dat_out_bypass_data[463:456];
  assign _0074_ = _0903_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17483" *) dat_out_bypass_data_w[455:448] : dat_out_bypass_data[455:448];
  assign _0073_ = _0902_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17473" *) dat_out_bypass_data_w[447:440] : dat_out_bypass_data[447:440];
  assign _0072_ = _0901_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17463" *) dat_out_bypass_data_w[439:432] : dat_out_bypass_data[439:432];
  assign _0071_ = _0900_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17453" *) dat_out_bypass_data_w[431:424] : dat_out_bypass_data[431:424];
  assign _0070_ = _0899_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17443" *) dat_out_bypass_data_w[423:416] : dat_out_bypass_data[423:416];
  assign _0069_ = _0898_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17433" *) dat_out_bypass_data_w[415:408] : dat_out_bypass_data[415:408];
  assign _0068_ = _0897_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17423" *) dat_out_bypass_data_w[407:400] : dat_out_bypass_data[407:400];
  assign _0066_ = _0896_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17413" *) dat_out_bypass_data_w[399:392] : dat_out_bypass_data[399:392];
  assign _0065_ = _0895_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17403" *) dat_out_bypass_data_w[391:384] : dat_out_bypass_data[391:384];
  assign _0064_ = _0894_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17393" *) dat_out_bypass_data_w[383:376] : dat_out_bypass_data[383:376];
  assign _0063_ = _0893_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17383" *) dat_out_bypass_data_w[375:368] : dat_out_bypass_data[375:368];
  assign _0062_ = _0892_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17373" *) dat_out_bypass_data_w[367:360] : dat_out_bypass_data[367:360];
  assign _0061_ = _0891_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17363" *) dat_out_bypass_data_w[359:352] : dat_out_bypass_data[359:352];
  assign _0060_ = _0890_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17353" *) dat_out_bypass_data_w[351:344] : dat_out_bypass_data[351:344];
  assign _0059_ = _0889_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17343" *) dat_out_bypass_data_w[343:336] : dat_out_bypass_data[343:336];
  assign _0058_ = _0888_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17333" *) dat_out_bypass_data_w[335:328] : dat_out_bypass_data[335:328];
  assign _0057_ = _0887_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17323" *) dat_out_bypass_data_w[327:320] : dat_out_bypass_data[327:320];
  assign _0055_ = _0886_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17313" *) dat_out_bypass_data_w[319:312] : dat_out_bypass_data[319:312];
  assign _0054_ = _0885_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17303" *) dat_out_bypass_data_w[311:304] : dat_out_bypass_data[311:304];
  assign _0053_ = _0884_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17293" *) dat_out_bypass_data_w[303:296] : dat_out_bypass_data[303:296];
  assign _0052_ = _0883_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17283" *) dat_out_bypass_data_w[295:288] : dat_out_bypass_data[295:288];
  assign _0051_ = _0882_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17273" *) dat_out_bypass_data_w[287:280] : dat_out_bypass_data[287:280];
  assign _0050_ = _0881_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17263" *) dat_out_bypass_data_w[279:272] : dat_out_bypass_data[279:272];
  assign _0049_ = _0880_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17253" *) dat_out_bypass_data_w[271:264] : dat_out_bypass_data[271:264];
  assign _0048_ = _0879_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17243" *) dat_out_bypass_data_w[263:256] : dat_out_bypass_data[263:256];
  assign _0047_ = _0878_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17233" *) dat_out_bypass_data_w[255:248] : dat_out_bypass_data[255:248];
  assign _0046_ = _0877_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17223" *) dat_out_bypass_data_w[247:240] : dat_out_bypass_data[247:240];
  assign _0044_ = _0876_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17213" *) dat_out_bypass_data_w[239:232] : dat_out_bypass_data[239:232];
  assign _0043_ = _0875_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17203" *) dat_out_bypass_data_w[231:224] : dat_out_bypass_data[231:224];
  assign _0042_ = _0874_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17193" *) dat_out_bypass_data_w[223:216] : dat_out_bypass_data[223:216];
  assign _0041_ = _0873_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17183" *) dat_out_bypass_data_w[215:208] : dat_out_bypass_data[215:208];
  assign _0040_ = _0872_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17173" *) dat_out_bypass_data_w[207:200] : dat_out_bypass_data[207:200];
  assign _0039_ = _0871_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17163" *) dat_out_bypass_data_w[199:192] : dat_out_bypass_data[199:192];
  assign _0038_ = _0870_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17153" *) dat_out_bypass_data_w[191:184] : dat_out_bypass_data[191:184];
  assign _0037_ = _0869_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17143" *) dat_out_bypass_data_w[183:176] : dat_out_bypass_data[183:176];
  assign _0036_ = _0868_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17133" *) dat_out_bypass_data_w[175:168] : dat_out_bypass_data[175:168];
  assign _0035_ = _0867_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17123" *) dat_out_bypass_data_w[167:160] : dat_out_bypass_data[167:160];
  assign _0033_ = _0866_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17113" *) dat_out_bypass_data_w[159:152] : dat_out_bypass_data[159:152];
  assign _0032_ = _0865_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17103" *) dat_out_bypass_data_w[151:144] : dat_out_bypass_data[151:144];
  assign _0031_ = _0864_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17093" *) dat_out_bypass_data_w[143:136] : dat_out_bypass_data[143:136];
  assign _0030_ = _0863_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17083" *) dat_out_bypass_data_w[135:128] : dat_out_bypass_data[135:128];
  assign _0029_ = _0862_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17073" *) dat_out_bypass_data_w[127:120] : dat_out_bypass_data[127:120];
  assign _0028_ = _0861_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17063" *) dat_out_bypass_data_w[119:112] : dat_out_bypass_data[119:112];
  assign _0027_ = _0860_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17053" *) dat_out_bypass_data_w[111:104] : dat_out_bypass_data[111:104];
  assign _0026_ = _0859_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17043" *) dat_out_bypass_data_w[103:96] : dat_out_bypass_data[103:96];
  assign _0145_ = _0858_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17033" *) dat_out_bypass_data_w[95:88] : dat_out_bypass_data[95:88];
  assign _0134_ = _0857_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17023" *) dat_out_bypass_data_w[87:80] : dat_out_bypass_data[87:80];
  assign _0122_ = _0856_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17013" *) dat_out_bypass_data_w[79:72] : dat_out_bypass_data[79:72];
  assign _0111_ = _0855_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:17003" *) dat_out_bypass_data_w[71:64] : dat_out_bypass_data[71:64];
  assign _0100_ = _0854_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16993" *) dat_out_bypass_data_w[63:56] : dat_out_bypass_data[63:56];
  assign _0089_ = _0853_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16983" *) dat_out_bypass_data_w[55:48] : dat_out_bypass_data[55:48];
  assign _0078_ = _0852_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16973" *) dat_out_bypass_data_w[47:40] : dat_out_bypass_data[47:40];
  assign _0067_ = _0851_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16963" *) dat_out_bypass_data_w[39:32] : dat_out_bypass_data[39:32];
  assign _0056_ = _0850_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16953" *) dat_out_bypass_data_w[31:24] : dat_out_bypass_data[31:24];
  assign _0045_ = _0849_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16943" *) dat_out_bypass_data_w[23:16] : dat_out_bypass_data[23:16];
  assign _0034_ = _0848_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16933" *) dat_out_bypass_data_w[15:8] : dat_out_bypass_data[15:8];
  assign _0123_ = _0847_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16923" *) dat_out_bypass_data_w[7:0] : dat_out_bypass_data[7:0];
  assign _0151_ = dat_out_bypass_p1_vld_w ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16865" *) dat_out_bypass_mask_w[127:64] : dat_out_bypass_mask[127:64];
  assign _0152_ = dat_out_bypass_p0_vld_w ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16804" *) dat_out_bypass_mask_w[63:0] : dat_out_bypass_mask[63:0];
  assign _0153_ = dat_out_pvld_w ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16743" *) dat_out_flag_w : dat_out_flag;
  assign _0158_ = dat_out_pvld_l4 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16669" *) dat_out_flag_l4 : dat_out_flag_l5;
  assign _0157_ = dat_out_pvld_l3 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16601" *) dat_out_flag_l3 : dat_out_flag_l4;
  assign _0156_ = dat_out_pvld_l2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16533" *) dat_out_flag_l2 : dat_out_flag_l3;
  assign _0155_ = dat_out_pvld_l1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16465" *) dat_out_flag_l1 : dat_out_flag_l2;
  assign _0154_ = dat_rsp_pvld ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16397" *) dat_rsp_pd[26:18] : dat_out_flag_l1;
  assign _0208_ = dat_rsp_sft_hi_d3_en ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16258" *) dat_rsp_l2_sft[255:128] : dat_rsp_l2_sft_d3[255:128];
  assign _0207_ = dat_rsp_sft_lo_d3_en ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16248" *) dat_rsp_l2_sft[127:0] : dat_rsp_l2_sft_d3[127:0];
  assign _0206_ = dat_rsp_sft_hi_d3_en ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16238" *) dat_rsp_l1_sft_d2[255:128] : dat_rsp_l1_sft_d3[255:128];
  assign _0205_ = dat_rsp_sft_lo_d3_en ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16228" *) dat_rsp_l1_sft_d2[127:0] : dat_rsp_l1_sft_d3[127:0];
  assign _0204_ = dat_rsp_sft_hi_d2_en ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16218" *) dat_rsp_l1_sft[255:128] : dat_rsp_l1_sft_d2[255:128];
  assign _0203_ = dat_rsp_sft_lo_d2_en ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16208" *) dat_rsp_l1_sft[127:0] : dat_rsp_l1_sft_d2[127:0];
  assign _0202_ = dat_rsp_sft_hi_d3_en ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16198" *) dat_rsp_l0_sft_d2[255:128] : dat_rsp_l0_sft_d3[255:128];
  assign _0201_ = dat_rsp_sft_lo_d3_en ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16188" *) dat_rsp_l0_sft_d2[127:0] : dat_rsp_l0_sft_d3[127:0];
  assign _0200_ = dat_rsp_sft_hi_d2_en ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16178" *) dat_rsp_l0_sft_d1[255:128] : dat_rsp_l0_sft_d2[255:128];
  assign _0199_ = dat_rsp_sft_lo_d2_en ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16168" *) dat_rsp_l0_sft_d1[127:0] : dat_rsp_l0_sft_d2[127:0];
  assign _0198_ = dat_rsp_sft_hi_d1_en ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16158" *) dat_rsp_l0_sft[511:256] : dat_rsp_l0_sft_d1[511:256];
  assign _0197_ = dat_rsp_sft_lo_d1_en ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16148" *) dat_rsp_l0_sft[255:0] : dat_rsp_l0_sft_d1[255:0];
  assign _0419_ = rsp_sft_cnt_l3_ori_en ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15697" *) rsp_sft_cnt_l3_w : rsp_sft_cnt_l3_ori;
  assign _0417_ = rsp_sft_cnt_l2_ori_en ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15636" *) rsp_sft_cnt_l2_w : rsp_sft_cnt_l2_ori;
  assign _0415_ = rsp_sft_cnt_l1_ori_en ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15575" *) rsp_sft_cnt_l1_w : rsp_sft_cnt_l1_ori;
  assign _0413_ = rsp_sft_cnt_l0_ori_en ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15514" *) rsp_sft_cnt_l0_w : rsp_sft_cnt_l0_ori;
  assign _0418_ = rsp_sft_cnt_l3_en ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15453" *) rsp_sft_cnt_l3_w : rsp_sft_cnt_l3;
  assign _0416_ = rsp_sft_cnt_l2_en ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15392" *) rsp_sft_cnt_l2_w : rsp_sft_cnt_l2;
  assign _0414_ = rsp_sft_cnt_l1_en ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15331" *) rsp_sft_cnt_l1_w : rsp_sft_cnt_l1;
  assign _0412_ = rsp_sft_cnt_l0_en ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15270" *) rsp_sft_cnt_l0_w : rsp_sft_cnt_l0;
  assign _0212_ = dat_rsp_pvld_d3 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:14978" *) dat_rsp_pd_d3 : dat_rsp_pd_d4;
  assign _0211_ = dat_rsp_pvld_d2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:14910" *) dat_rsp_pd_d2 : dat_rsp_pd_d3;
  assign _0210_ = dat_rsp_pvld_d1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:14842" *) dat_rsp_pd_d1 : dat_rsp_pd_d2;
  assign _0209_ = dat_rsp_pipe_pvld_d6 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:14774" *) { dat_rsp_pipe_pd_d6[28:19], dat_rsp_pipe_pd_d6[16:0] } : dat_rsp_pd_d1;
  assign _0021_ = dat_l3c1_en ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:14740" *) dat_l3c0_hi : dat_l3c1_hi;
  assign _0022_ = dat_l3c1_en ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:14740" *) dat_l3c0_lo : dat_l3c1_lo;
  assign _0017_ = dat_l2c1_en ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:14730" *) dat_l2c0_hi : dat_l2c1_hi;
  assign _0018_ = dat_l2c1_en ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:14730" *) dat_l2c0_lo : dat_l2c1_lo;
  assign _0013_ = dat_l1c1_hi_en ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:14720" *) dat_l1c0_hi : dat_l1c1_hi;
  assign _0014_ = dat_l1c1_en ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:14710" *) dat_l1c0_lo : dat_l1c1_lo;
  assign _0009_ = dat_l0c1_en ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:14700" *) dat_l0c0_hi : dat_l0c1_hi;
  assign _0010_ = dat_l0c1_en ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:14700" *) dat_l0c0_lo : dat_l0c1_lo;
  assign _0019_ = dat_l3c0_en ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:14690" *) sc2buf_dat_rd_data[1023:512] : dat_l3c0_hi;
  assign _0020_ = dat_l3c0_en ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:14690" *) sc2buf_dat_rd_data[511:0] : dat_l3c0_lo;
  assign _0015_ = dat_l2c0_en ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:14680" *) sc2buf_dat_rd_data[1023:512] : dat_l2c0_hi;
  assign _0016_ = dat_l2c0_en ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:14680" *) sc2buf_dat_rd_data[511:0] : dat_l2c0_lo;
  assign _0011_ = dat_l1c0_hi_en ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:14670" *) sc2buf_dat_rd_data[1023:512] : dat_l1c0_hi;
  assign _0012_ = dat_l1c0_en ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:14660" *) sc2buf_dat_rd_data[511:0] : dat_l1c0_lo;
  assign _0007_ = dat_l0c0_en ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:14650" *) sc2buf_dat_rd_data[1023:512] : dat_l0c0_hi;
  assign _0008_ = dat_l0c0_en ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:14650" *) sc2buf_dat_rd_data[511:0] : dat_l0c0_lo;
  assign _0196_ = dat_rsp_exec_pvld_d5 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:14402" *) dat_rsp_exec_sub_h_d5 : dat_rsp_exec_sub_h_d6;
  assign _0190_ = dat_rsp_exec_pvld_d5 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:14341" *) dat_rsp_exec_dummy_d5 : dat_rsp_exec_dummy_d6;
  assign _0218_ = dat_rsp_pipe_pvld_d5 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:14273" *) dat_rsp_pipe_pd_d5 : dat_rsp_pipe_pd_d6;
  assign _0195_ = dat_rsp_exec_pvld_d4 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:14205" *) dat_rsp_exec_sub_h_d4 : dat_rsp_exec_sub_h_d5;
  assign _0189_ = dat_rsp_exec_pvld_d4 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:14144" *) dat_rsp_exec_dummy_d4 : dat_rsp_exec_dummy_d5;
  assign _0217_ = dat_rsp_pipe_pvld_d4 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:14076" *) dat_rsp_pipe_pd_d4 : dat_rsp_pipe_pd_d5;
  assign _0194_ = dat_rsp_exec_pvld_d3 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:14008" *) dat_rsp_exec_sub_h_d3 : dat_rsp_exec_sub_h_d4;
  assign _0188_ = dat_rsp_exec_pvld_d3 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:13947" *) dat_rsp_exec_dummy_d3 : dat_rsp_exec_dummy_d4;
  assign _0216_ = dat_rsp_pipe_pvld_d3 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:13879" *) dat_rsp_pipe_pd_d3 : dat_rsp_pipe_pd_d4;
  assign _0193_ = dat_rsp_exec_pvld_d2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:13811" *) dat_rsp_exec_sub_h_d2 : dat_rsp_exec_sub_h_d3;
  assign _0187_ = dat_rsp_exec_pvld_d2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:13750" *) dat_rsp_exec_dummy_d2 : dat_rsp_exec_dummy_d3;
  assign _0215_ = dat_rsp_pipe_pvld_d2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:13682" *) dat_rsp_pipe_pd_d2 : dat_rsp_pipe_pd_d3;
  assign _0192_ = dat_rsp_exec_pvld_d1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:13614" *) dat_rsp_exec_sub_h_d1 : dat_rsp_exec_sub_h_d2;
  assign _0186_ = dat_rsp_exec_pvld_d1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:13553" *) dat_rsp_exec_dummy_d1 : dat_rsp_exec_dummy_d2;
  assign _0214_ = dat_rsp_pipe_pvld_d1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:13485" *) dat_rsp_pipe_pd_d1 : dat_rsp_pipe_pd_d2;
  assign _0191_ = dat_exec_valid_d2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:13417" *) dat_req_sub_h_d2 : dat_rsp_exec_sub_h_d1;
  assign _0185_ = dat_exec_valid_d2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:13356" *) dat_req_dummy_d2 : dat_rsp_exec_dummy_d1;
  assign _0213_ = dat_pipe_valid_d2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:13288" *) { dat_req_flag_d2, dat_req_rls_d2, dat_req_sub_w_st_d2, dat_req_dummy_d2, dat_req_cur_sub_h_d2, dat_req_bytes_d2, dat_req_ch_odd_d2, dat_req_ch_end_d2, dat_req_sub_c_d2, dat_req_sub_h_d2, dat_req_sub_w_d2 } : dat_rsp_pipe_pd_d1;
  assign _0170_ = dat_exec_valid_d1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:13138" *) dat_req_flag_d1 : dat_req_flag_d2;
  assign _0172_ = dat_exec_valid_d1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:13077" *) dat_req_rls_d1 : dat_req_rls_d2;
  assign _0184_ = dat_exec_valid_d1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:13016" *) dat_req_sub_w_st_d1 : dat_req_sub_w_st_d2;
  assign _0166_ = dat_exec_valid_d1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:12955" *) dat_req_cur_sub_h_d1 : dat_req_cur_sub_h_d2;
  assign _0168_ = dat_exec_valid_d1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:12894" *) dat_req_dummy_d1 : dat_req_dummy_d2;
  assign _0160_ = dat_exec_valid_d1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:12833" *) dat_req_bytes_d1 : dat_req_bytes_d2;
  assign _0164_ = dat_exec_valid_d1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:12772" *) dat_req_ch_odd_d1 : dat_req_ch_odd_d2;
  assign _0162_ = dat_exec_valid_d1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:12711" *) dat_req_ch_end_d1 : dat_req_ch_end_d2;
  assign _0174_ = dat_exec_valid_d1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:12650" *) dat_req_sub_c_d1 : dat_req_sub_c_d2;
  assign _0180_ = dat_exec_valid_d1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:12589" *) dat_req_sub_h_d1 : dat_req_sub_h_d2;
  assign _0182_ = dat_exec_valid_d1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:12528" *) dat_req_sub_w_d1 : dat_req_sub_w_d2;
  assign _0420_ = _1031_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:12453" *) dat_req_addr_w : sc2buf_dat_rd_addr;
  assign _0178_ = dat_req_sub_h_3_addr_en ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:12385" *) dat_req_addr_w : dat_req_sub_h_3_addr;
  assign _0177_ = dat_req_sub_h_2_addr_en ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:12324" *) dat_req_addr_w : dat_req_sub_h_2_addr;
  assign _0176_ = dat_req_sub_h_1_addr_en ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:12263" *) dat_req_addr_w : dat_req_sub_h_1_addr;
  assign _0175_ = dat_req_sub_h_0_addr_en ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:12202" *) dat_req_addr_w : dat_req_sub_h_0_addr;
  assign _0700_ = dat_exec_valid ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:11802" *) w_bias_w[13:2] : w_bias_d1;
  assign _0385_ = h_bias_reg_en[1] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:11741" *) h_bias_3_w : h_bias_3_d1;
  assign _0383_ = dat_exec_valid ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:11680" *) h_bias_2_w : h_bias_2_d1;
  assign _0381_ = dat_exec_valid ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:11619" *) h_bias_1_w : h_bias_1_d1;
  assign _0379_ = dat_exec_valid ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:11558" *) h_bias_0_w : h_bias_0_d1;
  assign _0003_ = c_bias_d1_reg_en ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:11497" *) c_bias : c_bias_d1;
  assign _0002_ = c_bias_reg_en ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:11436" *) c_bias_w : c_bias;
  assign _0396_ = dat_exec_valid ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:11168" *) pixel_force_clr : pixel_force_clr_d1;
  assign _0397_ = dat_exec_valid ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:11107" *) pixel_force_fetch : pixel_force_fetch_d1;
  assign _0171_ = dat_exec_valid ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:11046" *) _0743_ : dat_req_rls_d1;
  assign _0169_ = dat_exec_valid ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:10985" *) { dl_pd[29], dl_pd[27], dat_req_stripe_end, dat_req_stripe_st, batch_cnt } : dat_req_flag_d1;
  assign _0183_ = dat_req_sub_w_st_en ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:10924" *) dat_req_stripe_st : dat_req_sub_w_st_d1;
  assign _0165_ = dat_exec_valid ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:10863" *) dl_pd[25:24] : dat_req_cur_sub_h_d1;
  assign _0167_ = dat_exec_valid ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:10802" *) dat_req_dummy : dat_req_dummy_d1;
  assign _0163_ = dat_exec_valid ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:10741" *) pixel_req_ch_odd_w : dat_req_ch_odd_d1;
  assign _0161_ = dat_exec_valid ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:10680" *) is_last_channel : dat_req_ch_end_d1;
  assign _0173_ = dat_exec_valid ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:10619" *) dat_req_sub_c_w : dat_req_sub_c_d1;
  assign _0179_ = dat_exec_valid ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:10558" *) sub_h_cnt : dat_req_sub_h_d1;
  assign _0181_ = dat_exec_valid ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:10497" *) dat_req_sub_w_w : dat_req_sub_w_d1;
  assign _0228_ = datain_h_ori_reg_en ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:10345" *) datain_h_cnt_w : datain_h_ori;
  assign _0227_ = datain_h_cnt_reg_en ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:10284" *) datain_h_cnt_w : datain_h_cnt;
  assign _0399_ = pixel_ch_ori_reg_en ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:10114" *) pixel_req_ch_odd_w : pixel_req_ch_odd_ori;
  assign _0398_ = pixel_req_ch_odd_en ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:10053" *) pixel_req_ch_odd_w : pixel_req_ch_odd;
  assign _0400_ = pixel_ch_ori_reg_en ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:9992" *) pixel_w_cnt_w : pixel_w_ch_ori;
  assign _0402_ = pixel_req_ch_odd_en ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:9931" *) pixel_w_cnt_w : pixel_w_ori;
  assign _0401_ = pixel_w_cnt_reg_en ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:9870" *) pixel_w_cnt_w : pixel_w_cnt;
  assign _0231_ = datain_w_ori_reg_en ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:9809" *) datain_w_cnt_w : datain_w_ori;
  assign _0230_ = datain_w_cnt_reg_en ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:9748" *) datain_w_cnt_w : datain_w_cnt;
  assign _0225_ = c_bias_reg_en ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:9543" *) datain_c_cnt_w : datain_c_cnt;
  assign _0235_ = datain_h_ori_reg_en ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:9452" *) dataout_w_cnt_w : dataout_w_ori;
  assign _0234_ = dataout_w_cnt_reg_en ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:9391" *) dataout_w_cnt_w : dataout_w_cnt;
  assign _0159_ = dat_exec_valid ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:9182" *) dat_req_bytes : dat_req_bytes_d1;
  assign _0684_ = stripe_cnt_reg_en ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:8835" *) stripe_cnt_w : stripe_cnt;
  assign _0687_ = sub_h_cnt_reg_en ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:8734" *) sub_h_cnt_w : sub_h_cnt;
  assign _0001_ = _1061_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:8551" *) batch_cnt_w : batch_cnt;
  assign _0375_ = dl_pvld_d3 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:8442" *) dl_pd_d3 : dl_pd_d4;
  assign _0374_ = dl_pvld_d2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:8374" *) dl_pd_d2 : dl_pd_d3;
  assign _0373_ = dl_pvld_d1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:8306" *) dl_pd_d1 : dl_pd_d2;
  assign _0372_ = dl_in_pvld ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:8238" *) dl_pd_d0 : dl_pd_d1;
  assign _0241_ = dl_in_pvld_d4 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:8166" *) dl_in_pd_d4 : dl_in_pd_d5;
  assign _0240_ = dl_in_pvld_d3 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:8098" *) dl_in_pd_d3 : dl_in_pd_d4;
  assign _0239_ = dl_in_pvld_d2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:8030" *) dl_in_pd_d2 : dl_in_pd_d3;
  assign _0238_ = dl_in_pvld_d1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:7962" *) dl_in_pd_d1 : dl_in_pd_d2;
  assign _0237_ = sg2dl_pvld ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:7894" *) sg2dl_pd : dl_in_pd_d1;
  assign _0421_ = dat_rls ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:7536" *) sc2cdma_dat_entries_w : sc2cdma_dat_entries;
  assign _0422_ = dat_rls ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:7475" *) sc2cdma_dat_slices_w : sc2cdma_dat_slices;
  assign _0006_ = _1060_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:6884" *) dat_entry_st_w : dat_entry_st;
  assign _0408_ = layer_st ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:5284" *) { reg2dp_proc_precision, reg2dp_proc_precision, reg2dp_proc_precision, reg2dp_proc_precision } : pra_precision;
  assign _0409_ = layer_st ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:5223" *) { pra_truncate_w, pra_truncate_w, pra_truncate_w, pra_truncate_w } : pra_truncate;
  assign _0236_ = layer_st ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:5162" *) reg2dp_dataout_width : dataout_width_cmp;
  assign _0392_ = is_sg_done ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:5101" *) slice_entries_w : last_entries;
  assign _0393_ = is_sg_done ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:5040" *) slice_left : last_slices;
  assign _0683_ = layer_st ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:4979" *) slice_left_w : slice_left;
  assign _0410_ = layer_st_d1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:4918" *) slice_entries_w : rls_entries;
  assign _0411_ = layer_st ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:4857" *) rls_slices_w : rls_slices;
  assign _0386_ = layer_st_d1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:4796" *) entries : h_bias_3_stride;
  assign _0384_ = layer_st_d1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:4735" *) entries : h_bias_2_stride;
  assign _0382_ = layer_st_d1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:4674" *) h_bias_1_stride_w : h_bias_1_stride;
  assign _0380_ = layer_st_d1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:4613" *) h_bias_0_stride_w : h_bias_0_stride;
  assign _0387_ = layer_st ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:4552" *) h_offset_slice_w : h_offset_slice;
  assign _0378_ = layer_st ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:4491" *) reg2dp_entries : entries_cmp;
  assign _0377_ = layer_st ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:4430" *) entries_batch_w : entries_batch;
  assign _0376_ = layer_st ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:4369" *) entries_w : entries;
  assign _0394_ = layer_st ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:4308" *) reg2dp_pad_value : pad_value;
  assign _0702_ = layer_st ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:4247" *) y_dilate_w : y_dilate;
  assign _0701_ = layer_st ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:4186" *) x_dilate_w : x_dilate;
  assign _0395_ = layer_st ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:4125" *) { pixel_x_stride_w, 6'b000000 } : pixel_ch_stride;
  assign _0404_ = layer_st ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:4064" *) pixel_x_byte_stride_w : pixel_x_byte_stride;
  assign _0403_ = layer_st ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:4003" *) pixel_x_add_w : pixel_x_add;
  assign _0406_ = layer_st ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:3942" *) pixel_x_init_offset_w : pixel_x_init_offset;
  assign _0405_ = layer_st ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:3881" *) pixel_x_init_w : pixel_x_init;
  assign _0000_ = layer_st ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:3820" *) batch_cmp_w : batch_cmp;
  assign _0224_ = layer_st ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:3759" *) data_batch_w : data_batch;
  assign _0407_ = layer_st ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:3698" *) pixel_x_stride_w[0] : pixel_x_stride_odd;
  assign _0005_ = layer_st ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:3637" *) conv_y_stride_w : conv_y_stride;
  assign _0004_ = layer_st ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:3576" *) conv_x_stride_w : conv_x_stride;
  assign _0686_ = layer_st ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:3515" *) sub_h_cmp_w : sub_h_cmp_g1;
  assign _0685_ = layer_st ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:3454" *) sub_h_cmp_w : sub_h_cmp_g0;
  assign _0690_ = layer_st ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:3393" *) sub_h_total_w : sub_h_total_g11;
  assign _0689_ = layer_st ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:3332" *) sub_h_total_w : sub_h_total_g10;
  assign _0699_ = layer_st ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:3271" *) sub_h_total_w : sub_h_total_g9;
  assign _0698_ = layer_st ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:3210" *) sub_h_total_w : sub_h_total_g8;
  assign _0697_ = layer_st ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:3149" *) sub_h_total_w : sub_h_total_g7;
  assign _0696_ = layer_st ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:3088" *) sub_h_total_w : sub_h_total_g6;
  assign _0695_ = layer_st ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:3027" *) sub_h_total_w : sub_h_total_g5;
  assign _0694_ = layer_st ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:2966" *) sub_h_total_w : sub_h_total_g4;
  assign _0693_ = layer_st ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:2905" *) sub_h_total_w : sub_h_total_g3;
  assign _0692_ = layer_st ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:2844" *) sub_h_total_w[2:1] : sub_h_total_g2;
  assign _0691_ = layer_st ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:2783" *) sub_h_total_w : sub_h_total_g1;
  assign _0688_ = layer_st ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:2722" *) sub_h_total_w : sub_h_total_g0;
  assign _0226_ = layer_st ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:2661" *) datain_channel_cmp_w : datain_channel_cmp;
  assign _0229_ = layer_st ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:2600" *) reg2dp_datain_height_ext : datain_height_cmp;
  assign _0233_ = layer_st ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:2539" *) reg2dp_datain_width_ext : datain_width_cmp;
  assign _0232_ = layer_st ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:2478" *) datain_width_w : datain_width;
  assign _0223_ = layer_st ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:2417" *) data_bank_w : data_bank;
  assign _0388_ = layer_st ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:2356" *) { is_fp16, is_fp16 } : is_fp16_d1;
  assign _0390_ = layer_st ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:2295" *) { is_int8, is_int8, is_int8, is_int8, is_int8, is_int8, is_int8, is_int8, is_int8, is_int8, is_int8, is_int8, is_int8, is_int8, is_int8, is_int8, is_int8, is_int8, is_int8, is_int8, is_int8, is_int8, is_int8 } : is_int8_d1;
  assign _0389_ = layer_st ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:2234" *) { is_img, is_img, is_img, is_img, is_img, is_img, is_img, is_img, is_img, is_img, is_img, is_img, is_img, is_img, is_img, is_img, is_img, is_img, is_img, is_img, is_img, is_img, is_img, is_img, is_img, is_img, is_img, is_img, is_img, is_img, is_img, is_img, is_img, is_img } : is_img_d1;
  assign _0391_ = layer_st ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:2173" *) { reg2dp_conv_mode, reg2dp_conv_mode, reg2dp_conv_mode, reg2dp_conv_mode, reg2dp_conv_mode, reg2dp_conv_mode, reg2dp_conv_mode, reg2dp_conv_mode, reg2dp_conv_mode, reg2dp_conv_mode, reg2dp_conv_mode, reg2dp_conv_mode, reg2dp_conv_mode, reg2dp_conv_mode, reg2dp_conv_mode, reg2dp_conv_mode, reg2dp_conv_mode, reg2dp_conv_mode, reg2dp_conv_mode, reg2dp_conv_mode, reg2dp_conv_mode, reg2dp_conv_mode } : is_winograd_d1;
  assign _1157_ = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:10417" *) { datain_w_cur[2], datain_w_cur[3], datain_w_cur[4], datain_w_cur[5], datain_w_cur[6], datain_w_cur[7], datain_w_cur[8], datain_w_cur[9], datain_w_cur[10], datain_w_cur[11], datain_w_cur[12], datain_w_cur[13] };
  assign _1158_ = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:10417" *) { stripe_cnt[1], stripe_cnt[2], stripe_cnt[3], stripe_cnt[4], stripe_cnt[5], stripe_cnt[6] };
  assign _1159_ = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:14581" *) { sub_h_total_g2[0], sub_h_total_g2[1] };
  assign dat_rsp_mask_val_int8[56] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16327" *) { dat_out_bypass_data_w[448], dat_out_bypass_data_w[449], dat_out_bypass_data_w[450], dat_out_bypass_data_w[451], dat_out_bypass_data_w[452], dat_out_bypass_data_w[453], dat_out_bypass_data_w[454], dat_out_bypass_data_w[455] };
  assign dat_rsp_mask_val_int8[57] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16327" *) { dat_out_bypass_data_w[456], dat_out_bypass_data_w[457], dat_out_bypass_data_w[458], dat_out_bypass_data_w[459], dat_out_bypass_data_w[460], dat_out_bypass_data_w[461], dat_out_bypass_data_w[462], dat_out_bypass_data_w[463] };
  assign dat_rsp_mask_val_int8[58] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16327" *) { dat_out_bypass_data_w[464], dat_out_bypass_data_w[465], dat_out_bypass_data_w[466], dat_out_bypass_data_w[467], dat_out_bypass_data_w[468], dat_out_bypass_data_w[469], dat_out_bypass_data_w[470], dat_out_bypass_data_w[471] };
  assign dat_rsp_mask_val_int8[59] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16327" *) { dat_out_bypass_data_w[472], dat_out_bypass_data_w[473], dat_out_bypass_data_w[474], dat_out_bypass_data_w[475], dat_out_bypass_data_w[476], dat_out_bypass_data_w[477], dat_out_bypass_data_w[478], dat_out_bypass_data_w[479] };
  assign dat_rsp_mask_val_int8[60] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16327" *) { dat_out_bypass_data_w[480], dat_out_bypass_data_w[481], dat_out_bypass_data_w[482], dat_out_bypass_data_w[483], dat_out_bypass_data_w[484], dat_out_bypass_data_w[485], dat_out_bypass_data_w[486], dat_out_bypass_data_w[487] };
  assign dat_rsp_mask_val_int8[61] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16327" *) { dat_out_bypass_data_w[488], dat_out_bypass_data_w[489], dat_out_bypass_data_w[490], dat_out_bypass_data_w[491], dat_out_bypass_data_w[492], dat_out_bypass_data_w[493], dat_out_bypass_data_w[494], dat_out_bypass_data_w[495] };
  assign dat_rsp_mask_val_int8[62] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16327" *) { dat_out_bypass_data_w[496], dat_out_bypass_data_w[497], dat_out_bypass_data_w[498], dat_out_bypass_data_w[499], dat_out_bypass_data_w[500], dat_out_bypass_data_w[501], dat_out_bypass_data_w[502], dat_out_bypass_data_w[503] };
  assign dat_rsp_mask_val_int8[63] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16327" *) { dat_out_bypass_data_w[504], dat_out_bypass_data_w[505], dat_out_bypass_data_w[506], dat_out_bypass_data_w[507], dat_out_bypass_data_w[508], dat_out_bypass_data_w[509], dat_out_bypass_data_w[510], dat_out_bypass_data_w[511] };
  assign dat_rsp_mask_val_int8[48] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16328" *) { dat_out_bypass_data_w[384], dat_out_bypass_data_w[385], dat_out_bypass_data_w[386], dat_out_bypass_data_w[387], dat_out_bypass_data_w[388], dat_out_bypass_data_w[389], dat_out_bypass_data_w[390], dat_out_bypass_data_w[391] };
  assign dat_rsp_mask_val_int8[49] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16328" *) { dat_out_bypass_data_w[392], dat_out_bypass_data_w[393], dat_out_bypass_data_w[394], dat_out_bypass_data_w[395], dat_out_bypass_data_w[396], dat_out_bypass_data_w[397], dat_out_bypass_data_w[398], dat_out_bypass_data_w[399] };
  assign dat_rsp_mask_val_int8[50] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16328" *) { dat_out_bypass_data_w[400], dat_out_bypass_data_w[401], dat_out_bypass_data_w[402], dat_out_bypass_data_w[403], dat_out_bypass_data_w[404], dat_out_bypass_data_w[405], dat_out_bypass_data_w[406], dat_out_bypass_data_w[407] };
  assign dat_rsp_mask_val_int8[51] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16328" *) { dat_out_bypass_data_w[408], dat_out_bypass_data_w[409], dat_out_bypass_data_w[410], dat_out_bypass_data_w[411], dat_out_bypass_data_w[412], dat_out_bypass_data_w[413], dat_out_bypass_data_w[414], dat_out_bypass_data_w[415] };
  assign dat_rsp_mask_val_int8[52] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16328" *) { dat_out_bypass_data_w[416], dat_out_bypass_data_w[417], dat_out_bypass_data_w[418], dat_out_bypass_data_w[419], dat_out_bypass_data_w[420], dat_out_bypass_data_w[421], dat_out_bypass_data_w[422], dat_out_bypass_data_w[423] };
  assign dat_rsp_mask_val_int8[53] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16328" *) { dat_out_bypass_data_w[424], dat_out_bypass_data_w[425], dat_out_bypass_data_w[426], dat_out_bypass_data_w[427], dat_out_bypass_data_w[428], dat_out_bypass_data_w[429], dat_out_bypass_data_w[430], dat_out_bypass_data_w[431] };
  assign dat_rsp_mask_val_int8[54] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16328" *) { dat_out_bypass_data_w[432], dat_out_bypass_data_w[433], dat_out_bypass_data_w[434], dat_out_bypass_data_w[435], dat_out_bypass_data_w[436], dat_out_bypass_data_w[437], dat_out_bypass_data_w[438], dat_out_bypass_data_w[439] };
  assign dat_rsp_mask_val_int8[55] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16328" *) { dat_out_bypass_data_w[440], dat_out_bypass_data_w[441], dat_out_bypass_data_w[442], dat_out_bypass_data_w[443], dat_out_bypass_data_w[444], dat_out_bypass_data_w[445], dat_out_bypass_data_w[446], dat_out_bypass_data_w[447] };
  assign dat_rsp_mask_val_int8[40] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16329" *) { dat_out_bypass_data_w[320], dat_out_bypass_data_w[321], dat_out_bypass_data_w[322], dat_out_bypass_data_w[323], dat_out_bypass_data_w[324], dat_out_bypass_data_w[325], dat_out_bypass_data_w[326], dat_out_bypass_data_w[327] };
  assign dat_rsp_mask_val_int8[41] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16329" *) { dat_out_bypass_data_w[328], dat_out_bypass_data_w[329], dat_out_bypass_data_w[330], dat_out_bypass_data_w[331], dat_out_bypass_data_w[332], dat_out_bypass_data_w[333], dat_out_bypass_data_w[334], dat_out_bypass_data_w[335] };
  assign dat_rsp_mask_val_int8[42] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16329" *) { dat_out_bypass_data_w[336], dat_out_bypass_data_w[337], dat_out_bypass_data_w[338], dat_out_bypass_data_w[339], dat_out_bypass_data_w[340], dat_out_bypass_data_w[341], dat_out_bypass_data_w[342], dat_out_bypass_data_w[343] };
  assign dat_rsp_mask_val_int8[43] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16329" *) { dat_out_bypass_data_w[344], dat_out_bypass_data_w[345], dat_out_bypass_data_w[346], dat_out_bypass_data_w[347], dat_out_bypass_data_w[348], dat_out_bypass_data_w[349], dat_out_bypass_data_w[350], dat_out_bypass_data_w[351] };
  assign dat_rsp_mask_val_int8[44] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16329" *) { dat_out_bypass_data_w[352], dat_out_bypass_data_w[353], dat_out_bypass_data_w[354], dat_out_bypass_data_w[355], dat_out_bypass_data_w[356], dat_out_bypass_data_w[357], dat_out_bypass_data_w[358], dat_out_bypass_data_w[359] };
  assign dat_rsp_mask_val_int8[45] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16329" *) { dat_out_bypass_data_w[360], dat_out_bypass_data_w[361], dat_out_bypass_data_w[362], dat_out_bypass_data_w[363], dat_out_bypass_data_w[364], dat_out_bypass_data_w[365], dat_out_bypass_data_w[366], dat_out_bypass_data_w[367] };
  assign dat_rsp_mask_val_int8[46] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16329" *) { dat_out_bypass_data_w[368], dat_out_bypass_data_w[369], dat_out_bypass_data_w[370], dat_out_bypass_data_w[371], dat_out_bypass_data_w[372], dat_out_bypass_data_w[373], dat_out_bypass_data_w[374], dat_out_bypass_data_w[375] };
  assign dat_rsp_mask_val_int8[47] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16329" *) { dat_out_bypass_data_w[376], dat_out_bypass_data_w[377], dat_out_bypass_data_w[378], dat_out_bypass_data_w[379], dat_out_bypass_data_w[380], dat_out_bypass_data_w[381], dat_out_bypass_data_w[382], dat_out_bypass_data_w[383] };
  assign dat_rsp_mask_val_int8[32] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16330" *) { dat_out_bypass_data_w[256], dat_out_bypass_data_w[257], dat_out_bypass_data_w[258], dat_out_bypass_data_w[259], dat_out_bypass_data_w[260], dat_out_bypass_data_w[261], dat_out_bypass_data_w[262], dat_out_bypass_data_w[263] };
  assign dat_rsp_mask_val_int8[33] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16330" *) { dat_out_bypass_data_w[264], dat_out_bypass_data_w[265], dat_out_bypass_data_w[266], dat_out_bypass_data_w[267], dat_out_bypass_data_w[268], dat_out_bypass_data_w[269], dat_out_bypass_data_w[270], dat_out_bypass_data_w[271] };
  assign dat_rsp_mask_val_int8[34] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16330" *) { dat_out_bypass_data_w[272], dat_out_bypass_data_w[273], dat_out_bypass_data_w[274], dat_out_bypass_data_w[275], dat_out_bypass_data_w[276], dat_out_bypass_data_w[277], dat_out_bypass_data_w[278], dat_out_bypass_data_w[279] };
  assign dat_rsp_mask_val_int8[35] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16330" *) { dat_out_bypass_data_w[280], dat_out_bypass_data_w[281], dat_out_bypass_data_w[282], dat_out_bypass_data_w[283], dat_out_bypass_data_w[284], dat_out_bypass_data_w[285], dat_out_bypass_data_w[286], dat_out_bypass_data_w[287] };
  assign dat_rsp_mask_val_int8[36] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16330" *) { dat_out_bypass_data_w[288], dat_out_bypass_data_w[289], dat_out_bypass_data_w[290], dat_out_bypass_data_w[291], dat_out_bypass_data_w[292], dat_out_bypass_data_w[293], dat_out_bypass_data_w[294], dat_out_bypass_data_w[295] };
  assign dat_rsp_mask_val_int8[37] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16330" *) { dat_out_bypass_data_w[296], dat_out_bypass_data_w[297], dat_out_bypass_data_w[298], dat_out_bypass_data_w[299], dat_out_bypass_data_w[300], dat_out_bypass_data_w[301], dat_out_bypass_data_w[302], dat_out_bypass_data_w[303] };
  assign dat_rsp_mask_val_int8[38] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16330" *) { dat_out_bypass_data_w[304], dat_out_bypass_data_w[305], dat_out_bypass_data_w[306], dat_out_bypass_data_w[307], dat_out_bypass_data_w[308], dat_out_bypass_data_w[309], dat_out_bypass_data_w[310], dat_out_bypass_data_w[311] };
  assign dat_rsp_mask_val_int8[39] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16330" *) { dat_out_bypass_data_w[312], dat_out_bypass_data_w[313], dat_out_bypass_data_w[314], dat_out_bypass_data_w[315], dat_out_bypass_data_w[316], dat_out_bypass_data_w[317], dat_out_bypass_data_w[318], dat_out_bypass_data_w[319] };
  assign dat_rsp_mask_val_int8[24] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16331" *) { dat_out_bypass_data_w[192], dat_out_bypass_data_w[193], dat_out_bypass_data_w[194], dat_out_bypass_data_w[195], dat_out_bypass_data_w[196], dat_out_bypass_data_w[197], dat_out_bypass_data_w[198], dat_out_bypass_data_w[199] };
  assign dat_rsp_mask_val_int8[25] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16331" *) { dat_out_bypass_data_w[200], dat_out_bypass_data_w[201], dat_out_bypass_data_w[202], dat_out_bypass_data_w[203], dat_out_bypass_data_w[204], dat_out_bypass_data_w[205], dat_out_bypass_data_w[206], dat_out_bypass_data_w[207] };
  assign dat_rsp_mask_val_int8[26] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16331" *) { dat_out_bypass_data_w[208], dat_out_bypass_data_w[209], dat_out_bypass_data_w[210], dat_out_bypass_data_w[211], dat_out_bypass_data_w[212], dat_out_bypass_data_w[213], dat_out_bypass_data_w[214], dat_out_bypass_data_w[215] };
  assign dat_rsp_mask_val_int8[27] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16331" *) { dat_out_bypass_data_w[216], dat_out_bypass_data_w[217], dat_out_bypass_data_w[218], dat_out_bypass_data_w[219], dat_out_bypass_data_w[220], dat_out_bypass_data_w[221], dat_out_bypass_data_w[222], dat_out_bypass_data_w[223] };
  assign dat_rsp_mask_val_int8[28] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16331" *) { dat_out_bypass_data_w[224], dat_out_bypass_data_w[225], dat_out_bypass_data_w[226], dat_out_bypass_data_w[227], dat_out_bypass_data_w[228], dat_out_bypass_data_w[229], dat_out_bypass_data_w[230], dat_out_bypass_data_w[231] };
  assign dat_rsp_mask_val_int8[29] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16331" *) { dat_out_bypass_data_w[232], dat_out_bypass_data_w[233], dat_out_bypass_data_w[234], dat_out_bypass_data_w[235], dat_out_bypass_data_w[236], dat_out_bypass_data_w[237], dat_out_bypass_data_w[238], dat_out_bypass_data_w[239] };
  assign dat_rsp_mask_val_int8[30] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16331" *) { dat_out_bypass_data_w[240], dat_out_bypass_data_w[241], dat_out_bypass_data_w[242], dat_out_bypass_data_w[243], dat_out_bypass_data_w[244], dat_out_bypass_data_w[245], dat_out_bypass_data_w[246], dat_out_bypass_data_w[247] };
  assign dat_rsp_mask_val_int8[31] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16331" *) { dat_out_bypass_data_w[248], dat_out_bypass_data_w[249], dat_out_bypass_data_w[250], dat_out_bypass_data_w[251], dat_out_bypass_data_w[252], dat_out_bypass_data_w[253], dat_out_bypass_data_w[254], dat_out_bypass_data_w[255] };
  assign dat_rsp_mask_val_int8[16] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16332" *) { dat_out_bypass_data_w[128], dat_out_bypass_data_w[129], dat_out_bypass_data_w[130], dat_out_bypass_data_w[131], dat_out_bypass_data_w[132], dat_out_bypass_data_w[133], dat_out_bypass_data_w[134], dat_out_bypass_data_w[135] };
  assign dat_rsp_mask_val_int8[17] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16332" *) { dat_out_bypass_data_w[136], dat_out_bypass_data_w[137], dat_out_bypass_data_w[138], dat_out_bypass_data_w[139], dat_out_bypass_data_w[140], dat_out_bypass_data_w[141], dat_out_bypass_data_w[142], dat_out_bypass_data_w[143] };
  assign dat_rsp_mask_val_int8[18] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16332" *) { dat_out_bypass_data_w[144], dat_out_bypass_data_w[145], dat_out_bypass_data_w[146], dat_out_bypass_data_w[147], dat_out_bypass_data_w[148], dat_out_bypass_data_w[149], dat_out_bypass_data_w[150], dat_out_bypass_data_w[151] };
  assign dat_rsp_mask_val_int8[19] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16332" *) { dat_out_bypass_data_w[152], dat_out_bypass_data_w[153], dat_out_bypass_data_w[154], dat_out_bypass_data_w[155], dat_out_bypass_data_w[156], dat_out_bypass_data_w[157], dat_out_bypass_data_w[158], dat_out_bypass_data_w[159] };
  assign dat_rsp_mask_val_int8[20] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16332" *) { dat_out_bypass_data_w[160], dat_out_bypass_data_w[161], dat_out_bypass_data_w[162], dat_out_bypass_data_w[163], dat_out_bypass_data_w[164], dat_out_bypass_data_w[165], dat_out_bypass_data_w[166], dat_out_bypass_data_w[167] };
  assign dat_rsp_mask_val_int8[21] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16332" *) { dat_out_bypass_data_w[168], dat_out_bypass_data_w[169], dat_out_bypass_data_w[170], dat_out_bypass_data_w[171], dat_out_bypass_data_w[172], dat_out_bypass_data_w[173], dat_out_bypass_data_w[174], dat_out_bypass_data_w[175] };
  assign dat_rsp_mask_val_int8[22] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16332" *) { dat_out_bypass_data_w[176], dat_out_bypass_data_w[177], dat_out_bypass_data_w[178], dat_out_bypass_data_w[179], dat_out_bypass_data_w[180], dat_out_bypass_data_w[181], dat_out_bypass_data_w[182], dat_out_bypass_data_w[183] };
  assign dat_rsp_mask_val_int8[23] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16332" *) { dat_out_bypass_data_w[184], dat_out_bypass_data_w[185], dat_out_bypass_data_w[186], dat_out_bypass_data_w[187], dat_out_bypass_data_w[188], dat_out_bypass_data_w[189], dat_out_bypass_data_w[190], dat_out_bypass_data_w[191] };
  assign dat_rsp_mask_val_int8[8] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16333" *) { dat_out_bypass_data_w[64], dat_out_bypass_data_w[65], dat_out_bypass_data_w[66], dat_out_bypass_data_w[67], dat_out_bypass_data_w[68], dat_out_bypass_data_w[69], dat_out_bypass_data_w[70], dat_out_bypass_data_w[71] };
  assign dat_rsp_mask_val_int8[9] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16333" *) { dat_out_bypass_data_w[72], dat_out_bypass_data_w[73], dat_out_bypass_data_w[74], dat_out_bypass_data_w[75], dat_out_bypass_data_w[76], dat_out_bypass_data_w[77], dat_out_bypass_data_w[78], dat_out_bypass_data_w[79] };
  assign dat_rsp_mask_val_int8[10] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16333" *) { dat_out_bypass_data_w[80], dat_out_bypass_data_w[81], dat_out_bypass_data_w[82], dat_out_bypass_data_w[83], dat_out_bypass_data_w[84], dat_out_bypass_data_w[85], dat_out_bypass_data_w[86], dat_out_bypass_data_w[87] };
  assign dat_rsp_mask_val_int8[11] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16333" *) { dat_out_bypass_data_w[88], dat_out_bypass_data_w[89], dat_out_bypass_data_w[90], dat_out_bypass_data_w[91], dat_out_bypass_data_w[92], dat_out_bypass_data_w[93], dat_out_bypass_data_w[94], dat_out_bypass_data_w[95] };
  assign dat_rsp_mask_val_int8[12] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16333" *) { dat_out_bypass_data_w[96], dat_out_bypass_data_w[97], dat_out_bypass_data_w[98], dat_out_bypass_data_w[99], dat_out_bypass_data_w[100], dat_out_bypass_data_w[101], dat_out_bypass_data_w[102], dat_out_bypass_data_w[103] };
  assign dat_rsp_mask_val_int8[13] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16333" *) { dat_out_bypass_data_w[104], dat_out_bypass_data_w[105], dat_out_bypass_data_w[106], dat_out_bypass_data_w[107], dat_out_bypass_data_w[108], dat_out_bypass_data_w[109], dat_out_bypass_data_w[110], dat_out_bypass_data_w[111] };
  assign dat_rsp_mask_val_int8[14] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16333" *) { dat_out_bypass_data_w[112], dat_out_bypass_data_w[113], dat_out_bypass_data_w[114], dat_out_bypass_data_w[115], dat_out_bypass_data_w[116], dat_out_bypass_data_w[117], dat_out_bypass_data_w[118], dat_out_bypass_data_w[119] };
  assign dat_rsp_mask_val_int8[15] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16333" *) { dat_out_bypass_data_w[120], dat_out_bypass_data_w[121], dat_out_bypass_data_w[122], dat_out_bypass_data_w[123], dat_out_bypass_data_w[124], dat_out_bypass_data_w[125], dat_out_bypass_data_w[126], dat_out_bypass_data_w[127] };
  assign dat_rsp_mask_val_int8[0] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16334" *) { dat_out_bypass_data_w[0], dat_out_bypass_data_w[1], dat_out_bypass_data_w[2], dat_out_bypass_data_w[3], dat_out_bypass_data_w[4], dat_out_bypass_data_w[5], dat_out_bypass_data_w[6], dat_out_bypass_data_w[7] };
  assign dat_rsp_mask_val_int8[1] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16334" *) { dat_out_bypass_data_w[8], dat_out_bypass_data_w[9], dat_out_bypass_data_w[10], dat_out_bypass_data_w[11], dat_out_bypass_data_w[12], dat_out_bypass_data_w[13], dat_out_bypass_data_w[14], dat_out_bypass_data_w[15] };
  assign dat_rsp_mask_val_int8[2] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16334" *) { dat_out_bypass_data_w[16], dat_out_bypass_data_w[17], dat_out_bypass_data_w[18], dat_out_bypass_data_w[19], dat_out_bypass_data_w[20], dat_out_bypass_data_w[21], dat_out_bypass_data_w[22], dat_out_bypass_data_w[23] };
  assign dat_rsp_mask_val_int8[3] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16334" *) { dat_out_bypass_data_w[24], dat_out_bypass_data_w[25], dat_out_bypass_data_w[26], dat_out_bypass_data_w[27], dat_out_bypass_data_w[28], dat_out_bypass_data_w[29], dat_out_bypass_data_w[30], dat_out_bypass_data_w[31] };
  assign dat_rsp_mask_val_int8[4] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16334" *) { dat_out_bypass_data_w[32], dat_out_bypass_data_w[33], dat_out_bypass_data_w[34], dat_out_bypass_data_w[35], dat_out_bypass_data_w[36], dat_out_bypass_data_w[37], dat_out_bypass_data_w[38], dat_out_bypass_data_w[39] };
  assign dat_rsp_mask_val_int8[5] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16334" *) { dat_out_bypass_data_w[40], dat_out_bypass_data_w[41], dat_out_bypass_data_w[42], dat_out_bypass_data_w[43], dat_out_bypass_data_w[44], dat_out_bypass_data_w[45], dat_out_bypass_data_w[46], dat_out_bypass_data_w[47] };
  assign dat_rsp_mask_val_int8[6] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16334" *) { dat_out_bypass_data_w[48], dat_out_bypass_data_w[49], dat_out_bypass_data_w[50], dat_out_bypass_data_w[51], dat_out_bypass_data_w[52], dat_out_bypass_data_w[53], dat_out_bypass_data_w[54], dat_out_bypass_data_w[55] };
  assign dat_rsp_mask_val_int8[7] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16334" *) { dat_out_bypass_data_w[56], dat_out_bypass_data_w[57], dat_out_bypass_data_w[58], dat_out_bypass_data_w[59], dat_out_bypass_data_w[60], dat_out_bypass_data_w[61], dat_out_bypass_data_w[62], dat_out_bypass_data_w[63] };
  assign dat_rsp_mask_val_fp16[113] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16339" *) { dat_out_bypass_data_w[896], dat_out_bypass_data_w[897], dat_out_bypass_data_w[898], dat_out_bypass_data_w[899], dat_out_bypass_data_w[900], dat_out_bypass_data_w[901], dat_out_bypass_data_w[902], dat_out_bypass_data_w[903], dat_out_bypass_data_w[904], dat_out_bypass_data_w[905], dat_out_bypass_data_w[906], dat_out_bypass_data_w[907], dat_out_bypass_data_w[908], dat_out_bypass_data_w[909], dat_out_bypass_data_w[910] };
  assign dat_rsp_mask_val_fp16[115] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16339" *) { dat_out_bypass_data_w[912], dat_out_bypass_data_w[913], dat_out_bypass_data_w[914], dat_out_bypass_data_w[915], dat_out_bypass_data_w[916], dat_out_bypass_data_w[917], dat_out_bypass_data_w[918], dat_out_bypass_data_w[919], dat_out_bypass_data_w[920], dat_out_bypass_data_w[921], dat_out_bypass_data_w[922], dat_out_bypass_data_w[923], dat_out_bypass_data_w[924], dat_out_bypass_data_w[925], dat_out_bypass_data_w[926] };
  assign dat_rsp_mask_val_fp16[117] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16339" *) { dat_out_bypass_data_w[928], dat_out_bypass_data_w[929], dat_out_bypass_data_w[930], dat_out_bypass_data_w[931], dat_out_bypass_data_w[932], dat_out_bypass_data_w[933], dat_out_bypass_data_w[934], dat_out_bypass_data_w[935], dat_out_bypass_data_w[936], dat_out_bypass_data_w[937], dat_out_bypass_data_w[938], dat_out_bypass_data_w[939], dat_out_bypass_data_w[940], dat_out_bypass_data_w[941], dat_out_bypass_data_w[942] };
  assign dat_rsp_mask_val_fp16[119] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16339" *) { dat_out_bypass_data_w[944], dat_out_bypass_data_w[945], dat_out_bypass_data_w[946], dat_out_bypass_data_w[947], dat_out_bypass_data_w[948], dat_out_bypass_data_w[949], dat_out_bypass_data_w[950], dat_out_bypass_data_w[951], dat_out_bypass_data_w[952], dat_out_bypass_data_w[953], dat_out_bypass_data_w[954], dat_out_bypass_data_w[955], dat_out_bypass_data_w[956], dat_out_bypass_data_w[957], dat_out_bypass_data_w[958] };
  assign dat_rsp_mask_val_fp16[121] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16339" *) { dat_out_bypass_data_w[960], dat_out_bypass_data_w[961], dat_out_bypass_data_w[962], dat_out_bypass_data_w[963], dat_out_bypass_data_w[964], dat_out_bypass_data_w[965], dat_out_bypass_data_w[966], dat_out_bypass_data_w[967], dat_out_bypass_data_w[968], dat_out_bypass_data_w[969], dat_out_bypass_data_w[970], dat_out_bypass_data_w[971], dat_out_bypass_data_w[972], dat_out_bypass_data_w[973], dat_out_bypass_data_w[974] };
  assign dat_rsp_mask_val_fp16[123] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16339" *) { dat_out_bypass_data_w[976], dat_out_bypass_data_w[977], dat_out_bypass_data_w[978], dat_out_bypass_data_w[979], dat_out_bypass_data_w[980], dat_out_bypass_data_w[981], dat_out_bypass_data_w[982], dat_out_bypass_data_w[983], dat_out_bypass_data_w[984], dat_out_bypass_data_w[985], dat_out_bypass_data_w[986], dat_out_bypass_data_w[987], dat_out_bypass_data_w[988], dat_out_bypass_data_w[989], dat_out_bypass_data_w[990] };
  assign dat_rsp_mask_val_fp16[125] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16339" *) { dat_out_bypass_data_w[992], dat_out_bypass_data_w[993], dat_out_bypass_data_w[994], dat_out_bypass_data_w[995], dat_out_bypass_data_w[996], dat_out_bypass_data_w[997], dat_out_bypass_data_w[998], dat_out_bypass_data_w[999], dat_out_bypass_data_w[1000], dat_out_bypass_data_w[1001], dat_out_bypass_data_w[1002], dat_out_bypass_data_w[1003], dat_out_bypass_data_w[1004], dat_out_bypass_data_w[1005], dat_out_bypass_data_w[1006] };
  assign dat_rsp_mask_val_fp16[127] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16339" *) { dat_out_bypass_data_w[1008], dat_out_bypass_data_w[1009], dat_out_bypass_data_w[1010], dat_out_bypass_data_w[1011], dat_out_bypass_data_w[1012], dat_out_bypass_data_w[1013], dat_out_bypass_data_w[1014], dat_out_bypass_data_w[1015], dat_out_bypass_data_w[1016], dat_out_bypass_data_w[1017], dat_out_bypass_data_w[1018], dat_out_bypass_data_w[1019], dat_out_bypass_data_w[1020], dat_out_bypass_data_w[1021], dat_out_bypass_data_w[1022] };
  assign dat_rsp_mask_val_fp16[97] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16340" *) { dat_out_bypass_data_w[768], dat_out_bypass_data_w[769], dat_out_bypass_data_w[770], dat_out_bypass_data_w[771], dat_out_bypass_data_w[772], dat_out_bypass_data_w[773], dat_out_bypass_data_w[774], dat_out_bypass_data_w[775], dat_out_bypass_data_w[776], dat_out_bypass_data_w[777], dat_out_bypass_data_w[778], dat_out_bypass_data_w[779], dat_out_bypass_data_w[780], dat_out_bypass_data_w[781], dat_out_bypass_data_w[782] };
  assign dat_rsp_mask_val_fp16[99] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16340" *) { dat_out_bypass_data_w[784], dat_out_bypass_data_w[785], dat_out_bypass_data_w[786], dat_out_bypass_data_w[787], dat_out_bypass_data_w[788], dat_out_bypass_data_w[789], dat_out_bypass_data_w[790], dat_out_bypass_data_w[791], dat_out_bypass_data_w[792], dat_out_bypass_data_w[793], dat_out_bypass_data_w[794], dat_out_bypass_data_w[795], dat_out_bypass_data_w[796], dat_out_bypass_data_w[797], dat_out_bypass_data_w[798] };
  assign dat_rsp_mask_val_fp16[101] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16340" *) { dat_out_bypass_data_w[800], dat_out_bypass_data_w[801], dat_out_bypass_data_w[802], dat_out_bypass_data_w[803], dat_out_bypass_data_w[804], dat_out_bypass_data_w[805], dat_out_bypass_data_w[806], dat_out_bypass_data_w[807], dat_out_bypass_data_w[808], dat_out_bypass_data_w[809], dat_out_bypass_data_w[810], dat_out_bypass_data_w[811], dat_out_bypass_data_w[812], dat_out_bypass_data_w[813], dat_out_bypass_data_w[814] };
  assign dat_rsp_mask_val_fp16[103] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16340" *) { dat_out_bypass_data_w[816], dat_out_bypass_data_w[817], dat_out_bypass_data_w[818], dat_out_bypass_data_w[819], dat_out_bypass_data_w[820], dat_out_bypass_data_w[821], dat_out_bypass_data_w[822], dat_out_bypass_data_w[823], dat_out_bypass_data_w[824], dat_out_bypass_data_w[825], dat_out_bypass_data_w[826], dat_out_bypass_data_w[827], dat_out_bypass_data_w[828], dat_out_bypass_data_w[829], dat_out_bypass_data_w[830] };
  assign dat_rsp_mask_val_fp16[105] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16340" *) { dat_out_bypass_data_w[832], dat_out_bypass_data_w[833], dat_out_bypass_data_w[834], dat_out_bypass_data_w[835], dat_out_bypass_data_w[836], dat_out_bypass_data_w[837], dat_out_bypass_data_w[838], dat_out_bypass_data_w[839], dat_out_bypass_data_w[840], dat_out_bypass_data_w[841], dat_out_bypass_data_w[842], dat_out_bypass_data_w[843], dat_out_bypass_data_w[844], dat_out_bypass_data_w[845], dat_out_bypass_data_w[846] };
  assign dat_rsp_mask_val_fp16[107] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16340" *) { dat_out_bypass_data_w[848], dat_out_bypass_data_w[849], dat_out_bypass_data_w[850], dat_out_bypass_data_w[851], dat_out_bypass_data_w[852], dat_out_bypass_data_w[853], dat_out_bypass_data_w[854], dat_out_bypass_data_w[855], dat_out_bypass_data_w[856], dat_out_bypass_data_w[857], dat_out_bypass_data_w[858], dat_out_bypass_data_w[859], dat_out_bypass_data_w[860], dat_out_bypass_data_w[861], dat_out_bypass_data_w[862] };
  assign dat_rsp_mask_val_fp16[109] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16340" *) { dat_out_bypass_data_w[864], dat_out_bypass_data_w[865], dat_out_bypass_data_w[866], dat_out_bypass_data_w[867], dat_out_bypass_data_w[868], dat_out_bypass_data_w[869], dat_out_bypass_data_w[870], dat_out_bypass_data_w[871], dat_out_bypass_data_w[872], dat_out_bypass_data_w[873], dat_out_bypass_data_w[874], dat_out_bypass_data_w[875], dat_out_bypass_data_w[876], dat_out_bypass_data_w[877], dat_out_bypass_data_w[878] };
  assign dat_rsp_mask_val_fp16[111] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16340" *) { dat_out_bypass_data_w[880], dat_out_bypass_data_w[881], dat_out_bypass_data_w[882], dat_out_bypass_data_w[883], dat_out_bypass_data_w[884], dat_out_bypass_data_w[885], dat_out_bypass_data_w[886], dat_out_bypass_data_w[887], dat_out_bypass_data_w[888], dat_out_bypass_data_w[889], dat_out_bypass_data_w[890], dat_out_bypass_data_w[891], dat_out_bypass_data_w[892], dat_out_bypass_data_w[893], dat_out_bypass_data_w[894] };
  assign dat_rsp_mask_val_fp16[81] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16341" *) { dat_out_bypass_data_w[640], dat_out_bypass_data_w[641], dat_out_bypass_data_w[642], dat_out_bypass_data_w[643], dat_out_bypass_data_w[644], dat_out_bypass_data_w[645], dat_out_bypass_data_w[646], dat_out_bypass_data_w[647], dat_out_bypass_data_w[648], dat_out_bypass_data_w[649], dat_out_bypass_data_w[650], dat_out_bypass_data_w[651], dat_out_bypass_data_w[652], dat_out_bypass_data_w[653], dat_out_bypass_data_w[654] };
  assign dat_rsp_mask_val_fp16[83] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16341" *) { dat_out_bypass_data_w[656], dat_out_bypass_data_w[657], dat_out_bypass_data_w[658], dat_out_bypass_data_w[659], dat_out_bypass_data_w[660], dat_out_bypass_data_w[661], dat_out_bypass_data_w[662], dat_out_bypass_data_w[663], dat_out_bypass_data_w[664], dat_out_bypass_data_w[665], dat_out_bypass_data_w[666], dat_out_bypass_data_w[667], dat_out_bypass_data_w[668], dat_out_bypass_data_w[669], dat_out_bypass_data_w[670] };
  assign dat_rsp_mask_val_fp16[85] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16341" *) { dat_out_bypass_data_w[672], dat_out_bypass_data_w[673], dat_out_bypass_data_w[674], dat_out_bypass_data_w[675], dat_out_bypass_data_w[676], dat_out_bypass_data_w[677], dat_out_bypass_data_w[678], dat_out_bypass_data_w[679], dat_out_bypass_data_w[680], dat_out_bypass_data_w[681], dat_out_bypass_data_w[682], dat_out_bypass_data_w[683], dat_out_bypass_data_w[684], dat_out_bypass_data_w[685], dat_out_bypass_data_w[686] };
  assign dat_rsp_mask_val_fp16[87] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16341" *) { dat_out_bypass_data_w[688], dat_out_bypass_data_w[689], dat_out_bypass_data_w[690], dat_out_bypass_data_w[691], dat_out_bypass_data_w[692], dat_out_bypass_data_w[693], dat_out_bypass_data_w[694], dat_out_bypass_data_w[695], dat_out_bypass_data_w[696], dat_out_bypass_data_w[697], dat_out_bypass_data_w[698], dat_out_bypass_data_w[699], dat_out_bypass_data_w[700], dat_out_bypass_data_w[701], dat_out_bypass_data_w[702] };
  assign dat_rsp_mask_val_fp16[89] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16341" *) { dat_out_bypass_data_w[704], dat_out_bypass_data_w[705], dat_out_bypass_data_w[706], dat_out_bypass_data_w[707], dat_out_bypass_data_w[708], dat_out_bypass_data_w[709], dat_out_bypass_data_w[710], dat_out_bypass_data_w[711], dat_out_bypass_data_w[712], dat_out_bypass_data_w[713], dat_out_bypass_data_w[714], dat_out_bypass_data_w[715], dat_out_bypass_data_w[716], dat_out_bypass_data_w[717], dat_out_bypass_data_w[718] };
  assign dat_rsp_mask_val_fp16[91] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16341" *) { dat_out_bypass_data_w[720], dat_out_bypass_data_w[721], dat_out_bypass_data_w[722], dat_out_bypass_data_w[723], dat_out_bypass_data_w[724], dat_out_bypass_data_w[725], dat_out_bypass_data_w[726], dat_out_bypass_data_w[727], dat_out_bypass_data_w[728], dat_out_bypass_data_w[729], dat_out_bypass_data_w[730], dat_out_bypass_data_w[731], dat_out_bypass_data_w[732], dat_out_bypass_data_w[733], dat_out_bypass_data_w[734] };
  assign dat_rsp_mask_val_fp16[93] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16341" *) { dat_out_bypass_data_w[736], dat_out_bypass_data_w[737], dat_out_bypass_data_w[738], dat_out_bypass_data_w[739], dat_out_bypass_data_w[740], dat_out_bypass_data_w[741], dat_out_bypass_data_w[742], dat_out_bypass_data_w[743], dat_out_bypass_data_w[744], dat_out_bypass_data_w[745], dat_out_bypass_data_w[746], dat_out_bypass_data_w[747], dat_out_bypass_data_w[748], dat_out_bypass_data_w[749], dat_out_bypass_data_w[750] };
  assign dat_rsp_mask_val_fp16[95] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16341" *) { dat_out_bypass_data_w[752], dat_out_bypass_data_w[753], dat_out_bypass_data_w[754], dat_out_bypass_data_w[755], dat_out_bypass_data_w[756], dat_out_bypass_data_w[757], dat_out_bypass_data_w[758], dat_out_bypass_data_w[759], dat_out_bypass_data_w[760], dat_out_bypass_data_w[761], dat_out_bypass_data_w[762], dat_out_bypass_data_w[763], dat_out_bypass_data_w[764], dat_out_bypass_data_w[765], dat_out_bypass_data_w[766] };
  assign dat_rsp_mask_val_fp16[65] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16342" *) { dat_out_bypass_data_w[512], dat_out_bypass_data_w[513], dat_out_bypass_data_w[514], dat_out_bypass_data_w[515], dat_out_bypass_data_w[516], dat_out_bypass_data_w[517], dat_out_bypass_data_w[518], dat_out_bypass_data_w[519], dat_out_bypass_data_w[520], dat_out_bypass_data_w[521], dat_out_bypass_data_w[522], dat_out_bypass_data_w[523], dat_out_bypass_data_w[524], dat_out_bypass_data_w[525], dat_out_bypass_data_w[526] };
  assign dat_rsp_mask_val_fp16[67] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16342" *) { dat_out_bypass_data_w[528], dat_out_bypass_data_w[529], dat_out_bypass_data_w[530], dat_out_bypass_data_w[531], dat_out_bypass_data_w[532], dat_out_bypass_data_w[533], dat_out_bypass_data_w[534], dat_out_bypass_data_w[535], dat_out_bypass_data_w[536], dat_out_bypass_data_w[537], dat_out_bypass_data_w[538], dat_out_bypass_data_w[539], dat_out_bypass_data_w[540], dat_out_bypass_data_w[541], dat_out_bypass_data_w[542] };
  assign dat_rsp_mask_val_fp16[69] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16342" *) { dat_out_bypass_data_w[544], dat_out_bypass_data_w[545], dat_out_bypass_data_w[546], dat_out_bypass_data_w[547], dat_out_bypass_data_w[548], dat_out_bypass_data_w[549], dat_out_bypass_data_w[550], dat_out_bypass_data_w[551], dat_out_bypass_data_w[552], dat_out_bypass_data_w[553], dat_out_bypass_data_w[554], dat_out_bypass_data_w[555], dat_out_bypass_data_w[556], dat_out_bypass_data_w[557], dat_out_bypass_data_w[558] };
  assign dat_rsp_mask_val_fp16[71] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16342" *) { dat_out_bypass_data_w[560], dat_out_bypass_data_w[561], dat_out_bypass_data_w[562], dat_out_bypass_data_w[563], dat_out_bypass_data_w[564], dat_out_bypass_data_w[565], dat_out_bypass_data_w[566], dat_out_bypass_data_w[567], dat_out_bypass_data_w[568], dat_out_bypass_data_w[569], dat_out_bypass_data_w[570], dat_out_bypass_data_w[571], dat_out_bypass_data_w[572], dat_out_bypass_data_w[573], dat_out_bypass_data_w[574] };
  assign dat_rsp_mask_val_fp16[73] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16342" *) { dat_out_bypass_data_w[576], dat_out_bypass_data_w[577], dat_out_bypass_data_w[578], dat_out_bypass_data_w[579], dat_out_bypass_data_w[580], dat_out_bypass_data_w[581], dat_out_bypass_data_w[582], dat_out_bypass_data_w[583], dat_out_bypass_data_w[584], dat_out_bypass_data_w[585], dat_out_bypass_data_w[586], dat_out_bypass_data_w[587], dat_out_bypass_data_w[588], dat_out_bypass_data_w[589], dat_out_bypass_data_w[590] };
  assign dat_rsp_mask_val_fp16[75] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16342" *) { dat_out_bypass_data_w[592], dat_out_bypass_data_w[593], dat_out_bypass_data_w[594], dat_out_bypass_data_w[595], dat_out_bypass_data_w[596], dat_out_bypass_data_w[597], dat_out_bypass_data_w[598], dat_out_bypass_data_w[599], dat_out_bypass_data_w[600], dat_out_bypass_data_w[601], dat_out_bypass_data_w[602], dat_out_bypass_data_w[603], dat_out_bypass_data_w[604], dat_out_bypass_data_w[605], dat_out_bypass_data_w[606] };
  assign dat_rsp_mask_val_fp16[77] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16342" *) { dat_out_bypass_data_w[608], dat_out_bypass_data_w[609], dat_out_bypass_data_w[610], dat_out_bypass_data_w[611], dat_out_bypass_data_w[612], dat_out_bypass_data_w[613], dat_out_bypass_data_w[614], dat_out_bypass_data_w[615], dat_out_bypass_data_w[616], dat_out_bypass_data_w[617], dat_out_bypass_data_w[618], dat_out_bypass_data_w[619], dat_out_bypass_data_w[620], dat_out_bypass_data_w[621], dat_out_bypass_data_w[622] };
  assign dat_rsp_mask_val_fp16[79] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16342" *) { dat_out_bypass_data_w[624], dat_out_bypass_data_w[625], dat_out_bypass_data_w[626], dat_out_bypass_data_w[627], dat_out_bypass_data_w[628], dat_out_bypass_data_w[629], dat_out_bypass_data_w[630], dat_out_bypass_data_w[631], dat_out_bypass_data_w[632], dat_out_bypass_data_w[633], dat_out_bypass_data_w[634], dat_out_bypass_data_w[635], dat_out_bypass_data_w[636], dat_out_bypass_data_w[637], dat_out_bypass_data_w[638] };
  assign dat_rsp_mask_val_fp16[49] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16343" *) { dat_out_bypass_data_w[384], dat_out_bypass_data_w[385], dat_out_bypass_data_w[386], dat_out_bypass_data_w[387], dat_out_bypass_data_w[388], dat_out_bypass_data_w[389], dat_out_bypass_data_w[390], dat_out_bypass_data_w[391], dat_out_bypass_data_w[392], dat_out_bypass_data_w[393], dat_out_bypass_data_w[394], dat_out_bypass_data_w[395], dat_out_bypass_data_w[396], dat_out_bypass_data_w[397], dat_out_bypass_data_w[398] };
  assign dat_rsp_mask_val_fp16[51] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16343" *) { dat_out_bypass_data_w[400], dat_out_bypass_data_w[401], dat_out_bypass_data_w[402], dat_out_bypass_data_w[403], dat_out_bypass_data_w[404], dat_out_bypass_data_w[405], dat_out_bypass_data_w[406], dat_out_bypass_data_w[407], dat_out_bypass_data_w[408], dat_out_bypass_data_w[409], dat_out_bypass_data_w[410], dat_out_bypass_data_w[411], dat_out_bypass_data_w[412], dat_out_bypass_data_w[413], dat_out_bypass_data_w[414] };
  assign dat_rsp_mask_val_fp16[53] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16343" *) { dat_out_bypass_data_w[416], dat_out_bypass_data_w[417], dat_out_bypass_data_w[418], dat_out_bypass_data_w[419], dat_out_bypass_data_w[420], dat_out_bypass_data_w[421], dat_out_bypass_data_w[422], dat_out_bypass_data_w[423], dat_out_bypass_data_w[424], dat_out_bypass_data_w[425], dat_out_bypass_data_w[426], dat_out_bypass_data_w[427], dat_out_bypass_data_w[428], dat_out_bypass_data_w[429], dat_out_bypass_data_w[430] };
  assign dat_rsp_mask_val_fp16[55] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16343" *) { dat_out_bypass_data_w[432], dat_out_bypass_data_w[433], dat_out_bypass_data_w[434], dat_out_bypass_data_w[435], dat_out_bypass_data_w[436], dat_out_bypass_data_w[437], dat_out_bypass_data_w[438], dat_out_bypass_data_w[439], dat_out_bypass_data_w[440], dat_out_bypass_data_w[441], dat_out_bypass_data_w[442], dat_out_bypass_data_w[443], dat_out_bypass_data_w[444], dat_out_bypass_data_w[445], dat_out_bypass_data_w[446] };
  assign dat_rsp_mask_val_fp16[57] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16343" *) { dat_out_bypass_data_w[448], dat_out_bypass_data_w[449], dat_out_bypass_data_w[450], dat_out_bypass_data_w[451], dat_out_bypass_data_w[452], dat_out_bypass_data_w[453], dat_out_bypass_data_w[454], dat_out_bypass_data_w[455], dat_out_bypass_data_w[456], dat_out_bypass_data_w[457], dat_out_bypass_data_w[458], dat_out_bypass_data_w[459], dat_out_bypass_data_w[460], dat_out_bypass_data_w[461], dat_out_bypass_data_w[462] };
  assign dat_rsp_mask_val_fp16[59] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16343" *) { dat_out_bypass_data_w[464], dat_out_bypass_data_w[465], dat_out_bypass_data_w[466], dat_out_bypass_data_w[467], dat_out_bypass_data_w[468], dat_out_bypass_data_w[469], dat_out_bypass_data_w[470], dat_out_bypass_data_w[471], dat_out_bypass_data_w[472], dat_out_bypass_data_w[473], dat_out_bypass_data_w[474], dat_out_bypass_data_w[475], dat_out_bypass_data_w[476], dat_out_bypass_data_w[477], dat_out_bypass_data_w[478] };
  assign dat_rsp_mask_val_fp16[61] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16343" *) { dat_out_bypass_data_w[480], dat_out_bypass_data_w[481], dat_out_bypass_data_w[482], dat_out_bypass_data_w[483], dat_out_bypass_data_w[484], dat_out_bypass_data_w[485], dat_out_bypass_data_w[486], dat_out_bypass_data_w[487], dat_out_bypass_data_w[488], dat_out_bypass_data_w[489], dat_out_bypass_data_w[490], dat_out_bypass_data_w[491], dat_out_bypass_data_w[492], dat_out_bypass_data_w[493], dat_out_bypass_data_w[494] };
  assign dat_rsp_mask_val_fp16[63] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16343" *) { dat_out_bypass_data_w[496], dat_out_bypass_data_w[497], dat_out_bypass_data_w[498], dat_out_bypass_data_w[499], dat_out_bypass_data_w[500], dat_out_bypass_data_w[501], dat_out_bypass_data_w[502], dat_out_bypass_data_w[503], dat_out_bypass_data_w[504], dat_out_bypass_data_w[505], dat_out_bypass_data_w[506], dat_out_bypass_data_w[507], dat_out_bypass_data_w[508], dat_out_bypass_data_w[509], dat_out_bypass_data_w[510] };
  assign dat_rsp_mask_val_fp16[33] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16344" *) { dat_out_bypass_data_w[256], dat_out_bypass_data_w[257], dat_out_bypass_data_w[258], dat_out_bypass_data_w[259], dat_out_bypass_data_w[260], dat_out_bypass_data_w[261], dat_out_bypass_data_w[262], dat_out_bypass_data_w[263], dat_out_bypass_data_w[264], dat_out_bypass_data_w[265], dat_out_bypass_data_w[266], dat_out_bypass_data_w[267], dat_out_bypass_data_w[268], dat_out_bypass_data_w[269], dat_out_bypass_data_w[270] };
  assign dat_rsp_mask_val_fp16[35] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16344" *) { dat_out_bypass_data_w[272], dat_out_bypass_data_w[273], dat_out_bypass_data_w[274], dat_out_bypass_data_w[275], dat_out_bypass_data_w[276], dat_out_bypass_data_w[277], dat_out_bypass_data_w[278], dat_out_bypass_data_w[279], dat_out_bypass_data_w[280], dat_out_bypass_data_w[281], dat_out_bypass_data_w[282], dat_out_bypass_data_w[283], dat_out_bypass_data_w[284], dat_out_bypass_data_w[285], dat_out_bypass_data_w[286] };
  assign dat_rsp_mask_val_fp16[37] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16344" *) { dat_out_bypass_data_w[288], dat_out_bypass_data_w[289], dat_out_bypass_data_w[290], dat_out_bypass_data_w[291], dat_out_bypass_data_w[292], dat_out_bypass_data_w[293], dat_out_bypass_data_w[294], dat_out_bypass_data_w[295], dat_out_bypass_data_w[296], dat_out_bypass_data_w[297], dat_out_bypass_data_w[298], dat_out_bypass_data_w[299], dat_out_bypass_data_w[300], dat_out_bypass_data_w[301], dat_out_bypass_data_w[302] };
  assign dat_rsp_mask_val_fp16[39] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16344" *) { dat_out_bypass_data_w[304], dat_out_bypass_data_w[305], dat_out_bypass_data_w[306], dat_out_bypass_data_w[307], dat_out_bypass_data_w[308], dat_out_bypass_data_w[309], dat_out_bypass_data_w[310], dat_out_bypass_data_w[311], dat_out_bypass_data_w[312], dat_out_bypass_data_w[313], dat_out_bypass_data_w[314], dat_out_bypass_data_w[315], dat_out_bypass_data_w[316], dat_out_bypass_data_w[317], dat_out_bypass_data_w[318] };
  assign dat_rsp_mask_val_fp16[41] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16344" *) { dat_out_bypass_data_w[320], dat_out_bypass_data_w[321], dat_out_bypass_data_w[322], dat_out_bypass_data_w[323], dat_out_bypass_data_w[324], dat_out_bypass_data_w[325], dat_out_bypass_data_w[326], dat_out_bypass_data_w[327], dat_out_bypass_data_w[328], dat_out_bypass_data_w[329], dat_out_bypass_data_w[330], dat_out_bypass_data_w[331], dat_out_bypass_data_w[332], dat_out_bypass_data_w[333], dat_out_bypass_data_w[334] };
  assign dat_rsp_mask_val_fp16[43] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16344" *) { dat_out_bypass_data_w[336], dat_out_bypass_data_w[337], dat_out_bypass_data_w[338], dat_out_bypass_data_w[339], dat_out_bypass_data_w[340], dat_out_bypass_data_w[341], dat_out_bypass_data_w[342], dat_out_bypass_data_w[343], dat_out_bypass_data_w[344], dat_out_bypass_data_w[345], dat_out_bypass_data_w[346], dat_out_bypass_data_w[347], dat_out_bypass_data_w[348], dat_out_bypass_data_w[349], dat_out_bypass_data_w[350] };
  assign dat_rsp_mask_val_fp16[45] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16344" *) { dat_out_bypass_data_w[352], dat_out_bypass_data_w[353], dat_out_bypass_data_w[354], dat_out_bypass_data_w[355], dat_out_bypass_data_w[356], dat_out_bypass_data_w[357], dat_out_bypass_data_w[358], dat_out_bypass_data_w[359], dat_out_bypass_data_w[360], dat_out_bypass_data_w[361], dat_out_bypass_data_w[362], dat_out_bypass_data_w[363], dat_out_bypass_data_w[364], dat_out_bypass_data_w[365], dat_out_bypass_data_w[366] };
  assign dat_rsp_mask_val_fp16[47] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16344" *) { dat_out_bypass_data_w[368], dat_out_bypass_data_w[369], dat_out_bypass_data_w[370], dat_out_bypass_data_w[371], dat_out_bypass_data_w[372], dat_out_bypass_data_w[373], dat_out_bypass_data_w[374], dat_out_bypass_data_w[375], dat_out_bypass_data_w[376], dat_out_bypass_data_w[377], dat_out_bypass_data_w[378], dat_out_bypass_data_w[379], dat_out_bypass_data_w[380], dat_out_bypass_data_w[381], dat_out_bypass_data_w[382] };
  assign dat_rsp_mask_val_fp16[17] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16345" *) { dat_out_bypass_data_w[128], dat_out_bypass_data_w[129], dat_out_bypass_data_w[130], dat_out_bypass_data_w[131], dat_out_bypass_data_w[132], dat_out_bypass_data_w[133], dat_out_bypass_data_w[134], dat_out_bypass_data_w[135], dat_out_bypass_data_w[136], dat_out_bypass_data_w[137], dat_out_bypass_data_w[138], dat_out_bypass_data_w[139], dat_out_bypass_data_w[140], dat_out_bypass_data_w[141], dat_out_bypass_data_w[142] };
  assign dat_rsp_mask_val_fp16[19] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16345" *) { dat_out_bypass_data_w[144], dat_out_bypass_data_w[145], dat_out_bypass_data_w[146], dat_out_bypass_data_w[147], dat_out_bypass_data_w[148], dat_out_bypass_data_w[149], dat_out_bypass_data_w[150], dat_out_bypass_data_w[151], dat_out_bypass_data_w[152], dat_out_bypass_data_w[153], dat_out_bypass_data_w[154], dat_out_bypass_data_w[155], dat_out_bypass_data_w[156], dat_out_bypass_data_w[157], dat_out_bypass_data_w[158] };
  assign dat_rsp_mask_val_fp16[21] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16345" *) { dat_out_bypass_data_w[160], dat_out_bypass_data_w[161], dat_out_bypass_data_w[162], dat_out_bypass_data_w[163], dat_out_bypass_data_w[164], dat_out_bypass_data_w[165], dat_out_bypass_data_w[166], dat_out_bypass_data_w[167], dat_out_bypass_data_w[168], dat_out_bypass_data_w[169], dat_out_bypass_data_w[170], dat_out_bypass_data_w[171], dat_out_bypass_data_w[172], dat_out_bypass_data_w[173], dat_out_bypass_data_w[174] };
  assign dat_rsp_mask_val_fp16[23] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16345" *) { dat_out_bypass_data_w[176], dat_out_bypass_data_w[177], dat_out_bypass_data_w[178], dat_out_bypass_data_w[179], dat_out_bypass_data_w[180], dat_out_bypass_data_w[181], dat_out_bypass_data_w[182], dat_out_bypass_data_w[183], dat_out_bypass_data_w[184], dat_out_bypass_data_w[185], dat_out_bypass_data_w[186], dat_out_bypass_data_w[187], dat_out_bypass_data_w[188], dat_out_bypass_data_w[189], dat_out_bypass_data_w[190] };
  assign dat_rsp_mask_val_fp16[25] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16345" *) { dat_out_bypass_data_w[192], dat_out_bypass_data_w[193], dat_out_bypass_data_w[194], dat_out_bypass_data_w[195], dat_out_bypass_data_w[196], dat_out_bypass_data_w[197], dat_out_bypass_data_w[198], dat_out_bypass_data_w[199], dat_out_bypass_data_w[200], dat_out_bypass_data_w[201], dat_out_bypass_data_w[202], dat_out_bypass_data_w[203], dat_out_bypass_data_w[204], dat_out_bypass_data_w[205], dat_out_bypass_data_w[206] };
  assign dat_rsp_mask_val_fp16[27] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16345" *) { dat_out_bypass_data_w[208], dat_out_bypass_data_w[209], dat_out_bypass_data_w[210], dat_out_bypass_data_w[211], dat_out_bypass_data_w[212], dat_out_bypass_data_w[213], dat_out_bypass_data_w[214], dat_out_bypass_data_w[215], dat_out_bypass_data_w[216], dat_out_bypass_data_w[217], dat_out_bypass_data_w[218], dat_out_bypass_data_w[219], dat_out_bypass_data_w[220], dat_out_bypass_data_w[221], dat_out_bypass_data_w[222] };
  assign dat_rsp_mask_val_fp16[29] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16345" *) { dat_out_bypass_data_w[224], dat_out_bypass_data_w[225], dat_out_bypass_data_w[226], dat_out_bypass_data_w[227], dat_out_bypass_data_w[228], dat_out_bypass_data_w[229], dat_out_bypass_data_w[230], dat_out_bypass_data_w[231], dat_out_bypass_data_w[232], dat_out_bypass_data_w[233], dat_out_bypass_data_w[234], dat_out_bypass_data_w[235], dat_out_bypass_data_w[236], dat_out_bypass_data_w[237], dat_out_bypass_data_w[238] };
  assign dat_rsp_mask_val_fp16[31] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16345" *) { dat_out_bypass_data_w[240], dat_out_bypass_data_w[241], dat_out_bypass_data_w[242], dat_out_bypass_data_w[243], dat_out_bypass_data_w[244], dat_out_bypass_data_w[245], dat_out_bypass_data_w[246], dat_out_bypass_data_w[247], dat_out_bypass_data_w[248], dat_out_bypass_data_w[249], dat_out_bypass_data_w[250], dat_out_bypass_data_w[251], dat_out_bypass_data_w[252], dat_out_bypass_data_w[253], dat_out_bypass_data_w[254] };
  assign dat_rsp_mask_val_fp16[1] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16346" *) { dat_out_bypass_data_w[0], dat_out_bypass_data_w[1], dat_out_bypass_data_w[2], dat_out_bypass_data_w[3], dat_out_bypass_data_w[4], dat_out_bypass_data_w[5], dat_out_bypass_data_w[6], dat_out_bypass_data_w[7], dat_out_bypass_data_w[8], dat_out_bypass_data_w[9], dat_out_bypass_data_w[10], dat_out_bypass_data_w[11], dat_out_bypass_data_w[12], dat_out_bypass_data_w[13], dat_out_bypass_data_w[14] };
  assign dat_rsp_mask_val_fp16[3] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16346" *) { dat_out_bypass_data_w[16], dat_out_bypass_data_w[17], dat_out_bypass_data_w[18], dat_out_bypass_data_w[19], dat_out_bypass_data_w[20], dat_out_bypass_data_w[21], dat_out_bypass_data_w[22], dat_out_bypass_data_w[23], dat_out_bypass_data_w[24], dat_out_bypass_data_w[25], dat_out_bypass_data_w[26], dat_out_bypass_data_w[27], dat_out_bypass_data_w[28], dat_out_bypass_data_w[29], dat_out_bypass_data_w[30] };
  assign dat_rsp_mask_val_fp16[5] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16346" *) { dat_out_bypass_data_w[32], dat_out_bypass_data_w[33], dat_out_bypass_data_w[34], dat_out_bypass_data_w[35], dat_out_bypass_data_w[36], dat_out_bypass_data_w[37], dat_out_bypass_data_w[38], dat_out_bypass_data_w[39], dat_out_bypass_data_w[40], dat_out_bypass_data_w[41], dat_out_bypass_data_w[42], dat_out_bypass_data_w[43], dat_out_bypass_data_w[44], dat_out_bypass_data_w[45], dat_out_bypass_data_w[46] };
  assign dat_rsp_mask_val_fp16[7] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16346" *) { dat_out_bypass_data_w[48], dat_out_bypass_data_w[49], dat_out_bypass_data_w[50], dat_out_bypass_data_w[51], dat_out_bypass_data_w[52], dat_out_bypass_data_w[53], dat_out_bypass_data_w[54], dat_out_bypass_data_w[55], dat_out_bypass_data_w[56], dat_out_bypass_data_w[57], dat_out_bypass_data_w[58], dat_out_bypass_data_w[59], dat_out_bypass_data_w[60], dat_out_bypass_data_w[61], dat_out_bypass_data_w[62] };
  assign dat_rsp_mask_val_fp16[9] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16346" *) { dat_out_bypass_data_w[64], dat_out_bypass_data_w[65], dat_out_bypass_data_w[66], dat_out_bypass_data_w[67], dat_out_bypass_data_w[68], dat_out_bypass_data_w[69], dat_out_bypass_data_w[70], dat_out_bypass_data_w[71], dat_out_bypass_data_w[72], dat_out_bypass_data_w[73], dat_out_bypass_data_w[74], dat_out_bypass_data_w[75], dat_out_bypass_data_w[76], dat_out_bypass_data_w[77], dat_out_bypass_data_w[78] };
  assign dat_rsp_mask_val_fp16[11] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16346" *) { dat_out_bypass_data_w[80], dat_out_bypass_data_w[81], dat_out_bypass_data_w[82], dat_out_bypass_data_w[83], dat_out_bypass_data_w[84], dat_out_bypass_data_w[85], dat_out_bypass_data_w[86], dat_out_bypass_data_w[87], dat_out_bypass_data_w[88], dat_out_bypass_data_w[89], dat_out_bypass_data_w[90], dat_out_bypass_data_w[91], dat_out_bypass_data_w[92], dat_out_bypass_data_w[93], dat_out_bypass_data_w[94] };
  assign dat_rsp_mask_val_fp16[13] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16346" *) { dat_out_bypass_data_w[96], dat_out_bypass_data_w[97], dat_out_bypass_data_w[98], dat_out_bypass_data_w[99], dat_out_bypass_data_w[100], dat_out_bypass_data_w[101], dat_out_bypass_data_w[102], dat_out_bypass_data_w[103], dat_out_bypass_data_w[104], dat_out_bypass_data_w[105], dat_out_bypass_data_w[106], dat_out_bypass_data_w[107], dat_out_bypass_data_w[108], dat_out_bypass_data_w[109], dat_out_bypass_data_w[110] };
  assign dat_rsp_mask_val_fp16[15] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16346" *) { dat_out_bypass_data_w[112], dat_out_bypass_data_w[113], dat_out_bypass_data_w[114], dat_out_bypass_data_w[115], dat_out_bypass_data_w[116], dat_out_bypass_data_w[117], dat_out_bypass_data_w[118], dat_out_bypass_data_w[119], dat_out_bypass_data_w[120], dat_out_bypass_data_w[121], dat_out_bypass_data_w[122], dat_out_bypass_data_w[123], dat_out_bypass_data_w[124], dat_out_bypass_data_w[125], dat_out_bypass_data_w[126] };
  assign dat_rsp_mask_val_int16[113] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16351" *) { dat_out_bypass_data_w[896], dat_out_bypass_data_w[897], dat_out_bypass_data_w[898], dat_out_bypass_data_w[899], dat_out_bypass_data_w[900], dat_out_bypass_data_w[901], dat_out_bypass_data_w[902], dat_out_bypass_data_w[903], dat_out_bypass_data_w[904], dat_out_bypass_data_w[905], dat_out_bypass_data_w[906], dat_out_bypass_data_w[907], dat_out_bypass_data_w[908], dat_out_bypass_data_w[909], dat_out_bypass_data_w[910], dat_out_bypass_data_w[911] };
  assign dat_rsp_mask_val_int16[115] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16351" *) { dat_out_bypass_data_w[912], dat_out_bypass_data_w[913], dat_out_bypass_data_w[914], dat_out_bypass_data_w[915], dat_out_bypass_data_w[916], dat_out_bypass_data_w[917], dat_out_bypass_data_w[918], dat_out_bypass_data_w[919], dat_out_bypass_data_w[920], dat_out_bypass_data_w[921], dat_out_bypass_data_w[922], dat_out_bypass_data_w[923], dat_out_bypass_data_w[924], dat_out_bypass_data_w[925], dat_out_bypass_data_w[926], dat_out_bypass_data_w[927] };
  assign dat_rsp_mask_val_int16[117] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16351" *) { dat_out_bypass_data_w[928], dat_out_bypass_data_w[929], dat_out_bypass_data_w[930], dat_out_bypass_data_w[931], dat_out_bypass_data_w[932], dat_out_bypass_data_w[933], dat_out_bypass_data_w[934], dat_out_bypass_data_w[935], dat_out_bypass_data_w[936], dat_out_bypass_data_w[937], dat_out_bypass_data_w[938], dat_out_bypass_data_w[939], dat_out_bypass_data_w[940], dat_out_bypass_data_w[941], dat_out_bypass_data_w[942], dat_out_bypass_data_w[943] };
  assign dat_rsp_mask_val_int16[119] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16351" *) { dat_out_bypass_data_w[944], dat_out_bypass_data_w[945], dat_out_bypass_data_w[946], dat_out_bypass_data_w[947], dat_out_bypass_data_w[948], dat_out_bypass_data_w[949], dat_out_bypass_data_w[950], dat_out_bypass_data_w[951], dat_out_bypass_data_w[952], dat_out_bypass_data_w[953], dat_out_bypass_data_w[954], dat_out_bypass_data_w[955], dat_out_bypass_data_w[956], dat_out_bypass_data_w[957], dat_out_bypass_data_w[958], dat_out_bypass_data_w[959] };
  assign dat_rsp_mask_val_int16[121] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16351" *) { dat_out_bypass_data_w[960], dat_out_bypass_data_w[961], dat_out_bypass_data_w[962], dat_out_bypass_data_w[963], dat_out_bypass_data_w[964], dat_out_bypass_data_w[965], dat_out_bypass_data_w[966], dat_out_bypass_data_w[967], dat_out_bypass_data_w[968], dat_out_bypass_data_w[969], dat_out_bypass_data_w[970], dat_out_bypass_data_w[971], dat_out_bypass_data_w[972], dat_out_bypass_data_w[973], dat_out_bypass_data_w[974], dat_out_bypass_data_w[975] };
  assign dat_rsp_mask_val_int16[123] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16351" *) { dat_out_bypass_data_w[976], dat_out_bypass_data_w[977], dat_out_bypass_data_w[978], dat_out_bypass_data_w[979], dat_out_bypass_data_w[980], dat_out_bypass_data_w[981], dat_out_bypass_data_w[982], dat_out_bypass_data_w[983], dat_out_bypass_data_w[984], dat_out_bypass_data_w[985], dat_out_bypass_data_w[986], dat_out_bypass_data_w[987], dat_out_bypass_data_w[988], dat_out_bypass_data_w[989], dat_out_bypass_data_w[990], dat_out_bypass_data_w[991] };
  assign dat_rsp_mask_val_int16[125] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16351" *) { dat_out_bypass_data_w[992], dat_out_bypass_data_w[993], dat_out_bypass_data_w[994], dat_out_bypass_data_w[995], dat_out_bypass_data_w[996], dat_out_bypass_data_w[997], dat_out_bypass_data_w[998], dat_out_bypass_data_w[999], dat_out_bypass_data_w[1000], dat_out_bypass_data_w[1001], dat_out_bypass_data_w[1002], dat_out_bypass_data_w[1003], dat_out_bypass_data_w[1004], dat_out_bypass_data_w[1005], dat_out_bypass_data_w[1006], dat_out_bypass_data_w[1007] };
  assign dat_rsp_mask_val_int16[127] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16351" *) { dat_out_bypass_data_w[1008], dat_out_bypass_data_w[1009], dat_out_bypass_data_w[1010], dat_out_bypass_data_w[1011], dat_out_bypass_data_w[1012], dat_out_bypass_data_w[1013], dat_out_bypass_data_w[1014], dat_out_bypass_data_w[1015], dat_out_bypass_data_w[1016], dat_out_bypass_data_w[1017], dat_out_bypass_data_w[1018], dat_out_bypass_data_w[1019], dat_out_bypass_data_w[1020], dat_out_bypass_data_w[1021], dat_out_bypass_data_w[1022], dat_out_bypass_data_w[1023] };
  assign dat_rsp_mask_val_int16[97] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16352" *) { dat_out_bypass_data_w[768], dat_out_bypass_data_w[769], dat_out_bypass_data_w[770], dat_out_bypass_data_w[771], dat_out_bypass_data_w[772], dat_out_bypass_data_w[773], dat_out_bypass_data_w[774], dat_out_bypass_data_w[775], dat_out_bypass_data_w[776], dat_out_bypass_data_w[777], dat_out_bypass_data_w[778], dat_out_bypass_data_w[779], dat_out_bypass_data_w[780], dat_out_bypass_data_w[781], dat_out_bypass_data_w[782], dat_out_bypass_data_w[783] };
  assign dat_rsp_mask_val_int16[99] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16352" *) { dat_out_bypass_data_w[784], dat_out_bypass_data_w[785], dat_out_bypass_data_w[786], dat_out_bypass_data_w[787], dat_out_bypass_data_w[788], dat_out_bypass_data_w[789], dat_out_bypass_data_w[790], dat_out_bypass_data_w[791], dat_out_bypass_data_w[792], dat_out_bypass_data_w[793], dat_out_bypass_data_w[794], dat_out_bypass_data_w[795], dat_out_bypass_data_w[796], dat_out_bypass_data_w[797], dat_out_bypass_data_w[798], dat_out_bypass_data_w[799] };
  assign dat_rsp_mask_val_int16[101] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16352" *) { dat_out_bypass_data_w[800], dat_out_bypass_data_w[801], dat_out_bypass_data_w[802], dat_out_bypass_data_w[803], dat_out_bypass_data_w[804], dat_out_bypass_data_w[805], dat_out_bypass_data_w[806], dat_out_bypass_data_w[807], dat_out_bypass_data_w[808], dat_out_bypass_data_w[809], dat_out_bypass_data_w[810], dat_out_bypass_data_w[811], dat_out_bypass_data_w[812], dat_out_bypass_data_w[813], dat_out_bypass_data_w[814], dat_out_bypass_data_w[815] };
  assign dat_rsp_mask_val_int16[103] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16352" *) { dat_out_bypass_data_w[816], dat_out_bypass_data_w[817], dat_out_bypass_data_w[818], dat_out_bypass_data_w[819], dat_out_bypass_data_w[820], dat_out_bypass_data_w[821], dat_out_bypass_data_w[822], dat_out_bypass_data_w[823], dat_out_bypass_data_w[824], dat_out_bypass_data_w[825], dat_out_bypass_data_w[826], dat_out_bypass_data_w[827], dat_out_bypass_data_w[828], dat_out_bypass_data_w[829], dat_out_bypass_data_w[830], dat_out_bypass_data_w[831] };
  assign dat_rsp_mask_val_int16[105] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16352" *) { dat_out_bypass_data_w[832], dat_out_bypass_data_w[833], dat_out_bypass_data_w[834], dat_out_bypass_data_w[835], dat_out_bypass_data_w[836], dat_out_bypass_data_w[837], dat_out_bypass_data_w[838], dat_out_bypass_data_w[839], dat_out_bypass_data_w[840], dat_out_bypass_data_w[841], dat_out_bypass_data_w[842], dat_out_bypass_data_w[843], dat_out_bypass_data_w[844], dat_out_bypass_data_w[845], dat_out_bypass_data_w[846], dat_out_bypass_data_w[847] };
  assign dat_rsp_mask_val_int16[107] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16352" *) { dat_out_bypass_data_w[848], dat_out_bypass_data_w[849], dat_out_bypass_data_w[850], dat_out_bypass_data_w[851], dat_out_bypass_data_w[852], dat_out_bypass_data_w[853], dat_out_bypass_data_w[854], dat_out_bypass_data_w[855], dat_out_bypass_data_w[856], dat_out_bypass_data_w[857], dat_out_bypass_data_w[858], dat_out_bypass_data_w[859], dat_out_bypass_data_w[860], dat_out_bypass_data_w[861], dat_out_bypass_data_w[862], dat_out_bypass_data_w[863] };
  assign dat_rsp_mask_val_int16[109] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16352" *) { dat_out_bypass_data_w[864], dat_out_bypass_data_w[865], dat_out_bypass_data_w[866], dat_out_bypass_data_w[867], dat_out_bypass_data_w[868], dat_out_bypass_data_w[869], dat_out_bypass_data_w[870], dat_out_bypass_data_w[871], dat_out_bypass_data_w[872], dat_out_bypass_data_w[873], dat_out_bypass_data_w[874], dat_out_bypass_data_w[875], dat_out_bypass_data_w[876], dat_out_bypass_data_w[877], dat_out_bypass_data_w[878], dat_out_bypass_data_w[879] };
  assign dat_rsp_mask_val_int16[111] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16352" *) { dat_out_bypass_data_w[880], dat_out_bypass_data_w[881], dat_out_bypass_data_w[882], dat_out_bypass_data_w[883], dat_out_bypass_data_w[884], dat_out_bypass_data_w[885], dat_out_bypass_data_w[886], dat_out_bypass_data_w[887], dat_out_bypass_data_w[888], dat_out_bypass_data_w[889], dat_out_bypass_data_w[890], dat_out_bypass_data_w[891], dat_out_bypass_data_w[892], dat_out_bypass_data_w[893], dat_out_bypass_data_w[894], dat_out_bypass_data_w[895] };
  assign dat_rsp_mask_val_int16[81] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16353" *) { dat_out_bypass_data_w[640], dat_out_bypass_data_w[641], dat_out_bypass_data_w[642], dat_out_bypass_data_w[643], dat_out_bypass_data_w[644], dat_out_bypass_data_w[645], dat_out_bypass_data_w[646], dat_out_bypass_data_w[647], dat_out_bypass_data_w[648], dat_out_bypass_data_w[649], dat_out_bypass_data_w[650], dat_out_bypass_data_w[651], dat_out_bypass_data_w[652], dat_out_bypass_data_w[653], dat_out_bypass_data_w[654], dat_out_bypass_data_w[655] };
  assign dat_rsp_mask_val_int16[83] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16353" *) { dat_out_bypass_data_w[656], dat_out_bypass_data_w[657], dat_out_bypass_data_w[658], dat_out_bypass_data_w[659], dat_out_bypass_data_w[660], dat_out_bypass_data_w[661], dat_out_bypass_data_w[662], dat_out_bypass_data_w[663], dat_out_bypass_data_w[664], dat_out_bypass_data_w[665], dat_out_bypass_data_w[666], dat_out_bypass_data_w[667], dat_out_bypass_data_w[668], dat_out_bypass_data_w[669], dat_out_bypass_data_w[670], dat_out_bypass_data_w[671] };
  assign dat_rsp_mask_val_int16[85] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16353" *) { dat_out_bypass_data_w[672], dat_out_bypass_data_w[673], dat_out_bypass_data_w[674], dat_out_bypass_data_w[675], dat_out_bypass_data_w[676], dat_out_bypass_data_w[677], dat_out_bypass_data_w[678], dat_out_bypass_data_w[679], dat_out_bypass_data_w[680], dat_out_bypass_data_w[681], dat_out_bypass_data_w[682], dat_out_bypass_data_w[683], dat_out_bypass_data_w[684], dat_out_bypass_data_w[685], dat_out_bypass_data_w[686], dat_out_bypass_data_w[687] };
  assign dat_rsp_mask_val_int16[87] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16353" *) { dat_out_bypass_data_w[688], dat_out_bypass_data_w[689], dat_out_bypass_data_w[690], dat_out_bypass_data_w[691], dat_out_bypass_data_w[692], dat_out_bypass_data_w[693], dat_out_bypass_data_w[694], dat_out_bypass_data_w[695], dat_out_bypass_data_w[696], dat_out_bypass_data_w[697], dat_out_bypass_data_w[698], dat_out_bypass_data_w[699], dat_out_bypass_data_w[700], dat_out_bypass_data_w[701], dat_out_bypass_data_w[702], dat_out_bypass_data_w[703] };
  assign dat_rsp_mask_val_int16[89] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16353" *) { dat_out_bypass_data_w[704], dat_out_bypass_data_w[705], dat_out_bypass_data_w[706], dat_out_bypass_data_w[707], dat_out_bypass_data_w[708], dat_out_bypass_data_w[709], dat_out_bypass_data_w[710], dat_out_bypass_data_w[711], dat_out_bypass_data_w[712], dat_out_bypass_data_w[713], dat_out_bypass_data_w[714], dat_out_bypass_data_w[715], dat_out_bypass_data_w[716], dat_out_bypass_data_w[717], dat_out_bypass_data_w[718], dat_out_bypass_data_w[719] };
  assign dat_rsp_mask_val_int16[91] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16353" *) { dat_out_bypass_data_w[720], dat_out_bypass_data_w[721], dat_out_bypass_data_w[722], dat_out_bypass_data_w[723], dat_out_bypass_data_w[724], dat_out_bypass_data_w[725], dat_out_bypass_data_w[726], dat_out_bypass_data_w[727], dat_out_bypass_data_w[728], dat_out_bypass_data_w[729], dat_out_bypass_data_w[730], dat_out_bypass_data_w[731], dat_out_bypass_data_w[732], dat_out_bypass_data_w[733], dat_out_bypass_data_w[734], dat_out_bypass_data_w[735] };
  assign dat_rsp_mask_val_int16[93] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16353" *) { dat_out_bypass_data_w[736], dat_out_bypass_data_w[737], dat_out_bypass_data_w[738], dat_out_bypass_data_w[739], dat_out_bypass_data_w[740], dat_out_bypass_data_w[741], dat_out_bypass_data_w[742], dat_out_bypass_data_w[743], dat_out_bypass_data_w[744], dat_out_bypass_data_w[745], dat_out_bypass_data_w[746], dat_out_bypass_data_w[747], dat_out_bypass_data_w[748], dat_out_bypass_data_w[749], dat_out_bypass_data_w[750], dat_out_bypass_data_w[751] };
  assign dat_rsp_mask_val_int16[95] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16353" *) { dat_out_bypass_data_w[752], dat_out_bypass_data_w[753], dat_out_bypass_data_w[754], dat_out_bypass_data_w[755], dat_out_bypass_data_w[756], dat_out_bypass_data_w[757], dat_out_bypass_data_w[758], dat_out_bypass_data_w[759], dat_out_bypass_data_w[760], dat_out_bypass_data_w[761], dat_out_bypass_data_w[762], dat_out_bypass_data_w[763], dat_out_bypass_data_w[764], dat_out_bypass_data_w[765], dat_out_bypass_data_w[766], dat_out_bypass_data_w[767] };
  assign dat_rsp_mask_val_int16[65] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16354" *) { dat_out_bypass_data_w[512], dat_out_bypass_data_w[513], dat_out_bypass_data_w[514], dat_out_bypass_data_w[515], dat_out_bypass_data_w[516], dat_out_bypass_data_w[517], dat_out_bypass_data_w[518], dat_out_bypass_data_w[519], dat_out_bypass_data_w[520], dat_out_bypass_data_w[521], dat_out_bypass_data_w[522], dat_out_bypass_data_w[523], dat_out_bypass_data_w[524], dat_out_bypass_data_w[525], dat_out_bypass_data_w[526], dat_out_bypass_data_w[527] };
  assign dat_rsp_mask_val_int16[67] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16354" *) { dat_out_bypass_data_w[528], dat_out_bypass_data_w[529], dat_out_bypass_data_w[530], dat_out_bypass_data_w[531], dat_out_bypass_data_w[532], dat_out_bypass_data_w[533], dat_out_bypass_data_w[534], dat_out_bypass_data_w[535], dat_out_bypass_data_w[536], dat_out_bypass_data_w[537], dat_out_bypass_data_w[538], dat_out_bypass_data_w[539], dat_out_bypass_data_w[540], dat_out_bypass_data_w[541], dat_out_bypass_data_w[542], dat_out_bypass_data_w[543] };
  assign dat_rsp_mask_val_int16[69] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16354" *) { dat_out_bypass_data_w[544], dat_out_bypass_data_w[545], dat_out_bypass_data_w[546], dat_out_bypass_data_w[547], dat_out_bypass_data_w[548], dat_out_bypass_data_w[549], dat_out_bypass_data_w[550], dat_out_bypass_data_w[551], dat_out_bypass_data_w[552], dat_out_bypass_data_w[553], dat_out_bypass_data_w[554], dat_out_bypass_data_w[555], dat_out_bypass_data_w[556], dat_out_bypass_data_w[557], dat_out_bypass_data_w[558], dat_out_bypass_data_w[559] };
  assign dat_rsp_mask_val_int16[71] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16354" *) { dat_out_bypass_data_w[560], dat_out_bypass_data_w[561], dat_out_bypass_data_w[562], dat_out_bypass_data_w[563], dat_out_bypass_data_w[564], dat_out_bypass_data_w[565], dat_out_bypass_data_w[566], dat_out_bypass_data_w[567], dat_out_bypass_data_w[568], dat_out_bypass_data_w[569], dat_out_bypass_data_w[570], dat_out_bypass_data_w[571], dat_out_bypass_data_w[572], dat_out_bypass_data_w[573], dat_out_bypass_data_w[574], dat_out_bypass_data_w[575] };
  assign dat_rsp_mask_val_int16[73] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16354" *) { dat_out_bypass_data_w[576], dat_out_bypass_data_w[577], dat_out_bypass_data_w[578], dat_out_bypass_data_w[579], dat_out_bypass_data_w[580], dat_out_bypass_data_w[581], dat_out_bypass_data_w[582], dat_out_bypass_data_w[583], dat_out_bypass_data_w[584], dat_out_bypass_data_w[585], dat_out_bypass_data_w[586], dat_out_bypass_data_w[587], dat_out_bypass_data_w[588], dat_out_bypass_data_w[589], dat_out_bypass_data_w[590], dat_out_bypass_data_w[591] };
  assign dat_rsp_mask_val_int16[75] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16354" *) { dat_out_bypass_data_w[592], dat_out_bypass_data_w[593], dat_out_bypass_data_w[594], dat_out_bypass_data_w[595], dat_out_bypass_data_w[596], dat_out_bypass_data_w[597], dat_out_bypass_data_w[598], dat_out_bypass_data_w[599], dat_out_bypass_data_w[600], dat_out_bypass_data_w[601], dat_out_bypass_data_w[602], dat_out_bypass_data_w[603], dat_out_bypass_data_w[604], dat_out_bypass_data_w[605], dat_out_bypass_data_w[606], dat_out_bypass_data_w[607] };
  assign dat_rsp_mask_val_int16[77] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16354" *) { dat_out_bypass_data_w[608], dat_out_bypass_data_w[609], dat_out_bypass_data_w[610], dat_out_bypass_data_w[611], dat_out_bypass_data_w[612], dat_out_bypass_data_w[613], dat_out_bypass_data_w[614], dat_out_bypass_data_w[615], dat_out_bypass_data_w[616], dat_out_bypass_data_w[617], dat_out_bypass_data_w[618], dat_out_bypass_data_w[619], dat_out_bypass_data_w[620], dat_out_bypass_data_w[621], dat_out_bypass_data_w[622], dat_out_bypass_data_w[623] };
  assign dat_rsp_mask_val_int16[79] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16354" *) { dat_out_bypass_data_w[624], dat_out_bypass_data_w[625], dat_out_bypass_data_w[626], dat_out_bypass_data_w[627], dat_out_bypass_data_w[628], dat_out_bypass_data_w[629], dat_out_bypass_data_w[630], dat_out_bypass_data_w[631], dat_out_bypass_data_w[632], dat_out_bypass_data_w[633], dat_out_bypass_data_w[634], dat_out_bypass_data_w[635], dat_out_bypass_data_w[636], dat_out_bypass_data_w[637], dat_out_bypass_data_w[638], dat_out_bypass_data_w[639] };
  assign dat_rsp_mask_val_int16[49] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16355" *) { dat_out_bypass_data_w[384], dat_out_bypass_data_w[385], dat_out_bypass_data_w[386], dat_out_bypass_data_w[387], dat_out_bypass_data_w[388], dat_out_bypass_data_w[389], dat_out_bypass_data_w[390], dat_out_bypass_data_w[391], dat_out_bypass_data_w[392], dat_out_bypass_data_w[393], dat_out_bypass_data_w[394], dat_out_bypass_data_w[395], dat_out_bypass_data_w[396], dat_out_bypass_data_w[397], dat_out_bypass_data_w[398], dat_out_bypass_data_w[399] };
  assign dat_rsp_mask_val_int16[51] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16355" *) { dat_out_bypass_data_w[400], dat_out_bypass_data_w[401], dat_out_bypass_data_w[402], dat_out_bypass_data_w[403], dat_out_bypass_data_w[404], dat_out_bypass_data_w[405], dat_out_bypass_data_w[406], dat_out_bypass_data_w[407], dat_out_bypass_data_w[408], dat_out_bypass_data_w[409], dat_out_bypass_data_w[410], dat_out_bypass_data_w[411], dat_out_bypass_data_w[412], dat_out_bypass_data_w[413], dat_out_bypass_data_w[414], dat_out_bypass_data_w[415] };
  assign dat_rsp_mask_val_int16[53] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16355" *) { dat_out_bypass_data_w[416], dat_out_bypass_data_w[417], dat_out_bypass_data_w[418], dat_out_bypass_data_w[419], dat_out_bypass_data_w[420], dat_out_bypass_data_w[421], dat_out_bypass_data_w[422], dat_out_bypass_data_w[423], dat_out_bypass_data_w[424], dat_out_bypass_data_w[425], dat_out_bypass_data_w[426], dat_out_bypass_data_w[427], dat_out_bypass_data_w[428], dat_out_bypass_data_w[429], dat_out_bypass_data_w[430], dat_out_bypass_data_w[431] };
  assign dat_rsp_mask_val_int16[55] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16355" *) { dat_out_bypass_data_w[432], dat_out_bypass_data_w[433], dat_out_bypass_data_w[434], dat_out_bypass_data_w[435], dat_out_bypass_data_w[436], dat_out_bypass_data_w[437], dat_out_bypass_data_w[438], dat_out_bypass_data_w[439], dat_out_bypass_data_w[440], dat_out_bypass_data_w[441], dat_out_bypass_data_w[442], dat_out_bypass_data_w[443], dat_out_bypass_data_w[444], dat_out_bypass_data_w[445], dat_out_bypass_data_w[446], dat_out_bypass_data_w[447] };
  assign dat_rsp_mask_val_int16[57] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16355" *) { dat_out_bypass_data_w[448], dat_out_bypass_data_w[449], dat_out_bypass_data_w[450], dat_out_bypass_data_w[451], dat_out_bypass_data_w[452], dat_out_bypass_data_w[453], dat_out_bypass_data_w[454], dat_out_bypass_data_w[455], dat_out_bypass_data_w[456], dat_out_bypass_data_w[457], dat_out_bypass_data_w[458], dat_out_bypass_data_w[459], dat_out_bypass_data_w[460], dat_out_bypass_data_w[461], dat_out_bypass_data_w[462], dat_out_bypass_data_w[463] };
  assign dat_rsp_mask_val_int16[59] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16355" *) { dat_out_bypass_data_w[464], dat_out_bypass_data_w[465], dat_out_bypass_data_w[466], dat_out_bypass_data_w[467], dat_out_bypass_data_w[468], dat_out_bypass_data_w[469], dat_out_bypass_data_w[470], dat_out_bypass_data_w[471], dat_out_bypass_data_w[472], dat_out_bypass_data_w[473], dat_out_bypass_data_w[474], dat_out_bypass_data_w[475], dat_out_bypass_data_w[476], dat_out_bypass_data_w[477], dat_out_bypass_data_w[478], dat_out_bypass_data_w[479] };
  assign dat_rsp_mask_val_int16[61] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16355" *) { dat_out_bypass_data_w[480], dat_out_bypass_data_w[481], dat_out_bypass_data_w[482], dat_out_bypass_data_w[483], dat_out_bypass_data_w[484], dat_out_bypass_data_w[485], dat_out_bypass_data_w[486], dat_out_bypass_data_w[487], dat_out_bypass_data_w[488], dat_out_bypass_data_w[489], dat_out_bypass_data_w[490], dat_out_bypass_data_w[491], dat_out_bypass_data_w[492], dat_out_bypass_data_w[493], dat_out_bypass_data_w[494], dat_out_bypass_data_w[495] };
  assign dat_rsp_mask_val_int16[63] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16355" *) { dat_out_bypass_data_w[496], dat_out_bypass_data_w[497], dat_out_bypass_data_w[498], dat_out_bypass_data_w[499], dat_out_bypass_data_w[500], dat_out_bypass_data_w[501], dat_out_bypass_data_w[502], dat_out_bypass_data_w[503], dat_out_bypass_data_w[504], dat_out_bypass_data_w[505], dat_out_bypass_data_w[506], dat_out_bypass_data_w[507], dat_out_bypass_data_w[508], dat_out_bypass_data_w[509], dat_out_bypass_data_w[510], dat_out_bypass_data_w[511] };
  assign dat_rsp_mask_val_int16[33] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16356" *) { dat_out_bypass_data_w[256], dat_out_bypass_data_w[257], dat_out_bypass_data_w[258], dat_out_bypass_data_w[259], dat_out_bypass_data_w[260], dat_out_bypass_data_w[261], dat_out_bypass_data_w[262], dat_out_bypass_data_w[263], dat_out_bypass_data_w[264], dat_out_bypass_data_w[265], dat_out_bypass_data_w[266], dat_out_bypass_data_w[267], dat_out_bypass_data_w[268], dat_out_bypass_data_w[269], dat_out_bypass_data_w[270], dat_out_bypass_data_w[271] };
  assign dat_rsp_mask_val_int16[35] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16356" *) { dat_out_bypass_data_w[272], dat_out_bypass_data_w[273], dat_out_bypass_data_w[274], dat_out_bypass_data_w[275], dat_out_bypass_data_w[276], dat_out_bypass_data_w[277], dat_out_bypass_data_w[278], dat_out_bypass_data_w[279], dat_out_bypass_data_w[280], dat_out_bypass_data_w[281], dat_out_bypass_data_w[282], dat_out_bypass_data_w[283], dat_out_bypass_data_w[284], dat_out_bypass_data_w[285], dat_out_bypass_data_w[286], dat_out_bypass_data_w[287] };
  assign dat_rsp_mask_val_int16[37] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16356" *) { dat_out_bypass_data_w[288], dat_out_bypass_data_w[289], dat_out_bypass_data_w[290], dat_out_bypass_data_w[291], dat_out_bypass_data_w[292], dat_out_bypass_data_w[293], dat_out_bypass_data_w[294], dat_out_bypass_data_w[295], dat_out_bypass_data_w[296], dat_out_bypass_data_w[297], dat_out_bypass_data_w[298], dat_out_bypass_data_w[299], dat_out_bypass_data_w[300], dat_out_bypass_data_w[301], dat_out_bypass_data_w[302], dat_out_bypass_data_w[303] };
  assign dat_rsp_mask_val_int16[39] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16356" *) { dat_out_bypass_data_w[304], dat_out_bypass_data_w[305], dat_out_bypass_data_w[306], dat_out_bypass_data_w[307], dat_out_bypass_data_w[308], dat_out_bypass_data_w[309], dat_out_bypass_data_w[310], dat_out_bypass_data_w[311], dat_out_bypass_data_w[312], dat_out_bypass_data_w[313], dat_out_bypass_data_w[314], dat_out_bypass_data_w[315], dat_out_bypass_data_w[316], dat_out_bypass_data_w[317], dat_out_bypass_data_w[318], dat_out_bypass_data_w[319] };
  assign dat_rsp_mask_val_int16[41] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16356" *) { dat_out_bypass_data_w[320], dat_out_bypass_data_w[321], dat_out_bypass_data_w[322], dat_out_bypass_data_w[323], dat_out_bypass_data_w[324], dat_out_bypass_data_w[325], dat_out_bypass_data_w[326], dat_out_bypass_data_w[327], dat_out_bypass_data_w[328], dat_out_bypass_data_w[329], dat_out_bypass_data_w[330], dat_out_bypass_data_w[331], dat_out_bypass_data_w[332], dat_out_bypass_data_w[333], dat_out_bypass_data_w[334], dat_out_bypass_data_w[335] };
  assign dat_rsp_mask_val_int16[43] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16356" *) { dat_out_bypass_data_w[336], dat_out_bypass_data_w[337], dat_out_bypass_data_w[338], dat_out_bypass_data_w[339], dat_out_bypass_data_w[340], dat_out_bypass_data_w[341], dat_out_bypass_data_w[342], dat_out_bypass_data_w[343], dat_out_bypass_data_w[344], dat_out_bypass_data_w[345], dat_out_bypass_data_w[346], dat_out_bypass_data_w[347], dat_out_bypass_data_w[348], dat_out_bypass_data_w[349], dat_out_bypass_data_w[350], dat_out_bypass_data_w[351] };
  assign dat_rsp_mask_val_int16[45] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16356" *) { dat_out_bypass_data_w[352], dat_out_bypass_data_w[353], dat_out_bypass_data_w[354], dat_out_bypass_data_w[355], dat_out_bypass_data_w[356], dat_out_bypass_data_w[357], dat_out_bypass_data_w[358], dat_out_bypass_data_w[359], dat_out_bypass_data_w[360], dat_out_bypass_data_w[361], dat_out_bypass_data_w[362], dat_out_bypass_data_w[363], dat_out_bypass_data_w[364], dat_out_bypass_data_w[365], dat_out_bypass_data_w[366], dat_out_bypass_data_w[367] };
  assign dat_rsp_mask_val_int16[47] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16356" *) { dat_out_bypass_data_w[368], dat_out_bypass_data_w[369], dat_out_bypass_data_w[370], dat_out_bypass_data_w[371], dat_out_bypass_data_w[372], dat_out_bypass_data_w[373], dat_out_bypass_data_w[374], dat_out_bypass_data_w[375], dat_out_bypass_data_w[376], dat_out_bypass_data_w[377], dat_out_bypass_data_w[378], dat_out_bypass_data_w[379], dat_out_bypass_data_w[380], dat_out_bypass_data_w[381], dat_out_bypass_data_w[382], dat_out_bypass_data_w[383] };
  assign dat_rsp_mask_val_int16[17] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16357" *) { dat_out_bypass_data_w[128], dat_out_bypass_data_w[129], dat_out_bypass_data_w[130], dat_out_bypass_data_w[131], dat_out_bypass_data_w[132], dat_out_bypass_data_w[133], dat_out_bypass_data_w[134], dat_out_bypass_data_w[135], dat_out_bypass_data_w[136], dat_out_bypass_data_w[137], dat_out_bypass_data_w[138], dat_out_bypass_data_w[139], dat_out_bypass_data_w[140], dat_out_bypass_data_w[141], dat_out_bypass_data_w[142], dat_out_bypass_data_w[143] };
  assign dat_rsp_mask_val_int16[19] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16357" *) { dat_out_bypass_data_w[144], dat_out_bypass_data_w[145], dat_out_bypass_data_w[146], dat_out_bypass_data_w[147], dat_out_bypass_data_w[148], dat_out_bypass_data_w[149], dat_out_bypass_data_w[150], dat_out_bypass_data_w[151], dat_out_bypass_data_w[152], dat_out_bypass_data_w[153], dat_out_bypass_data_w[154], dat_out_bypass_data_w[155], dat_out_bypass_data_w[156], dat_out_bypass_data_w[157], dat_out_bypass_data_w[158], dat_out_bypass_data_w[159] };
  assign dat_rsp_mask_val_int16[21] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16357" *) { dat_out_bypass_data_w[160], dat_out_bypass_data_w[161], dat_out_bypass_data_w[162], dat_out_bypass_data_w[163], dat_out_bypass_data_w[164], dat_out_bypass_data_w[165], dat_out_bypass_data_w[166], dat_out_bypass_data_w[167], dat_out_bypass_data_w[168], dat_out_bypass_data_w[169], dat_out_bypass_data_w[170], dat_out_bypass_data_w[171], dat_out_bypass_data_w[172], dat_out_bypass_data_w[173], dat_out_bypass_data_w[174], dat_out_bypass_data_w[175] };
  assign dat_rsp_mask_val_int16[23] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16357" *) { dat_out_bypass_data_w[176], dat_out_bypass_data_w[177], dat_out_bypass_data_w[178], dat_out_bypass_data_w[179], dat_out_bypass_data_w[180], dat_out_bypass_data_w[181], dat_out_bypass_data_w[182], dat_out_bypass_data_w[183], dat_out_bypass_data_w[184], dat_out_bypass_data_w[185], dat_out_bypass_data_w[186], dat_out_bypass_data_w[187], dat_out_bypass_data_w[188], dat_out_bypass_data_w[189], dat_out_bypass_data_w[190], dat_out_bypass_data_w[191] };
  assign dat_rsp_mask_val_int16[25] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16357" *) { dat_out_bypass_data_w[192], dat_out_bypass_data_w[193], dat_out_bypass_data_w[194], dat_out_bypass_data_w[195], dat_out_bypass_data_w[196], dat_out_bypass_data_w[197], dat_out_bypass_data_w[198], dat_out_bypass_data_w[199], dat_out_bypass_data_w[200], dat_out_bypass_data_w[201], dat_out_bypass_data_w[202], dat_out_bypass_data_w[203], dat_out_bypass_data_w[204], dat_out_bypass_data_w[205], dat_out_bypass_data_w[206], dat_out_bypass_data_w[207] };
  assign dat_rsp_mask_val_int16[27] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16357" *) { dat_out_bypass_data_w[208], dat_out_bypass_data_w[209], dat_out_bypass_data_w[210], dat_out_bypass_data_w[211], dat_out_bypass_data_w[212], dat_out_bypass_data_w[213], dat_out_bypass_data_w[214], dat_out_bypass_data_w[215], dat_out_bypass_data_w[216], dat_out_bypass_data_w[217], dat_out_bypass_data_w[218], dat_out_bypass_data_w[219], dat_out_bypass_data_w[220], dat_out_bypass_data_w[221], dat_out_bypass_data_w[222], dat_out_bypass_data_w[223] };
  assign dat_rsp_mask_val_int16[29] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16357" *) { dat_out_bypass_data_w[224], dat_out_bypass_data_w[225], dat_out_bypass_data_w[226], dat_out_bypass_data_w[227], dat_out_bypass_data_w[228], dat_out_bypass_data_w[229], dat_out_bypass_data_w[230], dat_out_bypass_data_w[231], dat_out_bypass_data_w[232], dat_out_bypass_data_w[233], dat_out_bypass_data_w[234], dat_out_bypass_data_w[235], dat_out_bypass_data_w[236], dat_out_bypass_data_w[237], dat_out_bypass_data_w[238], dat_out_bypass_data_w[239] };
  assign dat_rsp_mask_val_int16[31] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16357" *) { dat_out_bypass_data_w[240], dat_out_bypass_data_w[241], dat_out_bypass_data_w[242], dat_out_bypass_data_w[243], dat_out_bypass_data_w[244], dat_out_bypass_data_w[245], dat_out_bypass_data_w[246], dat_out_bypass_data_w[247], dat_out_bypass_data_w[248], dat_out_bypass_data_w[249], dat_out_bypass_data_w[250], dat_out_bypass_data_w[251], dat_out_bypass_data_w[252], dat_out_bypass_data_w[253], dat_out_bypass_data_w[254], dat_out_bypass_data_w[255] };
  assign dat_rsp_mask_val_int16[1] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16358" *) { dat_out_bypass_data_w[0], dat_out_bypass_data_w[1], dat_out_bypass_data_w[2], dat_out_bypass_data_w[3], dat_out_bypass_data_w[4], dat_out_bypass_data_w[5], dat_out_bypass_data_w[6], dat_out_bypass_data_w[7], dat_out_bypass_data_w[8], dat_out_bypass_data_w[9], dat_out_bypass_data_w[10], dat_out_bypass_data_w[11], dat_out_bypass_data_w[12], dat_out_bypass_data_w[13], dat_out_bypass_data_w[14], dat_out_bypass_data_w[15] };
  assign dat_rsp_mask_val_int16[3] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16358" *) { dat_out_bypass_data_w[16], dat_out_bypass_data_w[17], dat_out_bypass_data_w[18], dat_out_bypass_data_w[19], dat_out_bypass_data_w[20], dat_out_bypass_data_w[21], dat_out_bypass_data_w[22], dat_out_bypass_data_w[23], dat_out_bypass_data_w[24], dat_out_bypass_data_w[25], dat_out_bypass_data_w[26], dat_out_bypass_data_w[27], dat_out_bypass_data_w[28], dat_out_bypass_data_w[29], dat_out_bypass_data_w[30], dat_out_bypass_data_w[31] };
  assign dat_rsp_mask_val_int16[5] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16358" *) { dat_out_bypass_data_w[32], dat_out_bypass_data_w[33], dat_out_bypass_data_w[34], dat_out_bypass_data_w[35], dat_out_bypass_data_w[36], dat_out_bypass_data_w[37], dat_out_bypass_data_w[38], dat_out_bypass_data_w[39], dat_out_bypass_data_w[40], dat_out_bypass_data_w[41], dat_out_bypass_data_w[42], dat_out_bypass_data_w[43], dat_out_bypass_data_w[44], dat_out_bypass_data_w[45], dat_out_bypass_data_w[46], dat_out_bypass_data_w[47] };
  assign dat_rsp_mask_val_int16[7] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16358" *) { dat_out_bypass_data_w[48], dat_out_bypass_data_w[49], dat_out_bypass_data_w[50], dat_out_bypass_data_w[51], dat_out_bypass_data_w[52], dat_out_bypass_data_w[53], dat_out_bypass_data_w[54], dat_out_bypass_data_w[55], dat_out_bypass_data_w[56], dat_out_bypass_data_w[57], dat_out_bypass_data_w[58], dat_out_bypass_data_w[59], dat_out_bypass_data_w[60], dat_out_bypass_data_w[61], dat_out_bypass_data_w[62], dat_out_bypass_data_w[63] };
  assign dat_rsp_mask_val_int16[9] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16358" *) { dat_out_bypass_data_w[64], dat_out_bypass_data_w[65], dat_out_bypass_data_w[66], dat_out_bypass_data_w[67], dat_out_bypass_data_w[68], dat_out_bypass_data_w[69], dat_out_bypass_data_w[70], dat_out_bypass_data_w[71], dat_out_bypass_data_w[72], dat_out_bypass_data_w[73], dat_out_bypass_data_w[74], dat_out_bypass_data_w[75], dat_out_bypass_data_w[76], dat_out_bypass_data_w[77], dat_out_bypass_data_w[78], dat_out_bypass_data_w[79] };
  assign dat_rsp_mask_val_int16[11] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16358" *) { dat_out_bypass_data_w[80], dat_out_bypass_data_w[81], dat_out_bypass_data_w[82], dat_out_bypass_data_w[83], dat_out_bypass_data_w[84], dat_out_bypass_data_w[85], dat_out_bypass_data_w[86], dat_out_bypass_data_w[87], dat_out_bypass_data_w[88], dat_out_bypass_data_w[89], dat_out_bypass_data_w[90], dat_out_bypass_data_w[91], dat_out_bypass_data_w[92], dat_out_bypass_data_w[93], dat_out_bypass_data_w[94], dat_out_bypass_data_w[95] };
  assign dat_rsp_mask_val_int16[13] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16358" *) { dat_out_bypass_data_w[96], dat_out_bypass_data_w[97], dat_out_bypass_data_w[98], dat_out_bypass_data_w[99], dat_out_bypass_data_w[100], dat_out_bypass_data_w[101], dat_out_bypass_data_w[102], dat_out_bypass_data_w[103], dat_out_bypass_data_w[104], dat_out_bypass_data_w[105], dat_out_bypass_data_w[106], dat_out_bypass_data_w[107], dat_out_bypass_data_w[108], dat_out_bypass_data_w[109], dat_out_bypass_data_w[110], dat_out_bypass_data_w[111] };
  assign dat_rsp_mask_val_int16[15] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16358" *) { dat_out_bypass_data_w[112], dat_out_bypass_data_w[113], dat_out_bypass_data_w[114], dat_out_bypass_data_w[115], dat_out_bypass_data_w[116], dat_out_bypass_data_w[117], dat_out_bypass_data_w[118], dat_out_bypass_data_w[119], dat_out_bypass_data_w[120], dat_out_bypass_data_w[121], dat_out_bypass_data_w[122], dat_out_bypass_data_w[123], dat_out_bypass_data_w[124], dat_out_bypass_data_w[125], dat_out_bypass_data_w[126], dat_out_bypass_data_w[127] };
  assign dat_out_wg_mask_int8[56] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18382" *) { dat_out_wg_data[448], dat_out_wg_data[449], dat_out_wg_data[450], dat_out_wg_data[451], dat_out_wg_data[452], dat_out_wg_data[453], dat_out_wg_data[454], dat_out_wg_data[455] };
  assign dat_out_wg_mask_int8[57] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18382" *) { dat_out_wg_data[456], dat_out_wg_data[457], dat_out_wg_data[458], dat_out_wg_data[459], dat_out_wg_data[460], dat_out_wg_data[461], dat_out_wg_data[462], dat_out_wg_data[463] };
  assign dat_out_wg_mask_int8[58] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18382" *) { dat_out_wg_data[464], dat_out_wg_data[465], dat_out_wg_data[466], dat_out_wg_data[467], dat_out_wg_data[468], dat_out_wg_data[469], dat_out_wg_data[470], dat_out_wg_data[471] };
  assign dat_out_wg_mask_int8[59] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18382" *) { dat_out_wg_data[472], dat_out_wg_data[473], dat_out_wg_data[474], dat_out_wg_data[475], dat_out_wg_data[476], dat_out_wg_data[477], dat_out_wg_data[478], dat_out_wg_data[479] };
  assign dat_out_wg_mask_int8[60] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18382" *) { dat_out_wg_data[480], dat_out_wg_data[481], dat_out_wg_data[482], dat_out_wg_data[483], dat_out_wg_data[484], dat_out_wg_data[485], dat_out_wg_data[486], dat_out_wg_data[487] };
  assign dat_out_wg_mask_int8[61] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18382" *) { dat_out_wg_data[488], dat_out_wg_data[489], dat_out_wg_data[490], dat_out_wg_data[491], dat_out_wg_data[492], dat_out_wg_data[493], dat_out_wg_data[494], dat_out_wg_data[495] };
  assign dat_out_wg_mask_int8[62] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18382" *) { dat_out_wg_data[496], dat_out_wg_data[497], dat_out_wg_data[498], dat_out_wg_data[499], dat_out_wg_data[500], dat_out_wg_data[501], dat_out_wg_data[502], dat_out_wg_data[503] };
  assign dat_out_wg_mask_int8[63] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18382" *) { dat_out_wg_data[504], dat_out_wg_data[505], dat_out_wg_data[506], dat_out_wg_data[507], dat_out_wg_data[508], dat_out_wg_data[509], dat_out_wg_data[510], dat_out_wg_data[511] };
  assign dat_out_wg_mask_int8[48] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18383" *) { dat_out_wg_data[384], dat_out_wg_data[385], dat_out_wg_data[386], dat_out_wg_data[387], dat_out_wg_data[388], dat_out_wg_data[389], dat_out_wg_data[390], dat_out_wg_data[391] };
  assign dat_out_wg_mask_int8[49] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18383" *) { dat_out_wg_data[392], dat_out_wg_data[393], dat_out_wg_data[394], dat_out_wg_data[395], dat_out_wg_data[396], dat_out_wg_data[397], dat_out_wg_data[398], dat_out_wg_data[399] };
  assign dat_out_wg_mask_int8[50] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18383" *) { dat_out_wg_data[400], dat_out_wg_data[401], dat_out_wg_data[402], dat_out_wg_data[403], dat_out_wg_data[404], dat_out_wg_data[405], dat_out_wg_data[406], dat_out_wg_data[407] };
  assign dat_out_wg_mask_int8[51] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18383" *) { dat_out_wg_data[408], dat_out_wg_data[409], dat_out_wg_data[410], dat_out_wg_data[411], dat_out_wg_data[412], dat_out_wg_data[413], dat_out_wg_data[414], dat_out_wg_data[415] };
  assign dat_out_wg_mask_int8[52] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18383" *) { dat_out_wg_data[416], dat_out_wg_data[417], dat_out_wg_data[418], dat_out_wg_data[419], dat_out_wg_data[420], dat_out_wg_data[421], dat_out_wg_data[422], dat_out_wg_data[423] };
  assign dat_out_wg_mask_int8[53] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18383" *) { dat_out_wg_data[424], dat_out_wg_data[425], dat_out_wg_data[426], dat_out_wg_data[427], dat_out_wg_data[428], dat_out_wg_data[429], dat_out_wg_data[430], dat_out_wg_data[431] };
  assign dat_out_wg_mask_int8[54] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18383" *) { dat_out_wg_data[432], dat_out_wg_data[433], dat_out_wg_data[434], dat_out_wg_data[435], dat_out_wg_data[436], dat_out_wg_data[437], dat_out_wg_data[438], dat_out_wg_data[439] };
  assign dat_out_wg_mask_int8[55] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18383" *) { dat_out_wg_data[440], dat_out_wg_data[441], dat_out_wg_data[442], dat_out_wg_data[443], dat_out_wg_data[444], dat_out_wg_data[445], dat_out_wg_data[446], dat_out_wg_data[447] };
  assign dat_out_wg_mask_int8[40] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18384" *) { dat_out_wg_data[320], dat_out_wg_data[321], dat_out_wg_data[322], dat_out_wg_data[323], dat_out_wg_data[324], dat_out_wg_data[325], dat_out_wg_data[326], dat_out_wg_data[327] };
  assign dat_out_wg_mask_int8[41] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18384" *) { dat_out_wg_data[328], dat_out_wg_data[329], dat_out_wg_data[330], dat_out_wg_data[331], dat_out_wg_data[332], dat_out_wg_data[333], dat_out_wg_data[334], dat_out_wg_data[335] };
  assign dat_out_wg_mask_int8[42] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18384" *) { dat_out_wg_data[336], dat_out_wg_data[337], dat_out_wg_data[338], dat_out_wg_data[339], dat_out_wg_data[340], dat_out_wg_data[341], dat_out_wg_data[342], dat_out_wg_data[343] };
  assign dat_out_wg_mask_int8[43] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18384" *) { dat_out_wg_data[344], dat_out_wg_data[345], dat_out_wg_data[346], dat_out_wg_data[347], dat_out_wg_data[348], dat_out_wg_data[349], dat_out_wg_data[350], dat_out_wg_data[351] };
  assign dat_out_wg_mask_int8[44] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18384" *) { dat_out_wg_data[352], dat_out_wg_data[353], dat_out_wg_data[354], dat_out_wg_data[355], dat_out_wg_data[356], dat_out_wg_data[357], dat_out_wg_data[358], dat_out_wg_data[359] };
  assign dat_out_wg_mask_int8[45] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18384" *) { dat_out_wg_data[360], dat_out_wg_data[361], dat_out_wg_data[362], dat_out_wg_data[363], dat_out_wg_data[364], dat_out_wg_data[365], dat_out_wg_data[366], dat_out_wg_data[367] };
  assign dat_out_wg_mask_int8[46] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18384" *) { dat_out_wg_data[368], dat_out_wg_data[369], dat_out_wg_data[370], dat_out_wg_data[371], dat_out_wg_data[372], dat_out_wg_data[373], dat_out_wg_data[374], dat_out_wg_data[375] };
  assign dat_out_wg_mask_int8[47] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18384" *) { dat_out_wg_data[376], dat_out_wg_data[377], dat_out_wg_data[378], dat_out_wg_data[379], dat_out_wg_data[380], dat_out_wg_data[381], dat_out_wg_data[382], dat_out_wg_data[383] };
  assign dat_out_wg_mask_int8[32] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18385" *) { dat_out_wg_data[256], dat_out_wg_data[257], dat_out_wg_data[258], dat_out_wg_data[259], dat_out_wg_data[260], dat_out_wg_data[261], dat_out_wg_data[262], dat_out_wg_data[263] };
  assign dat_out_wg_mask_int8[33] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18385" *) { dat_out_wg_data[264], dat_out_wg_data[265], dat_out_wg_data[266], dat_out_wg_data[267], dat_out_wg_data[268], dat_out_wg_data[269], dat_out_wg_data[270], dat_out_wg_data[271] };
  assign dat_out_wg_mask_int8[34] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18385" *) { dat_out_wg_data[272], dat_out_wg_data[273], dat_out_wg_data[274], dat_out_wg_data[275], dat_out_wg_data[276], dat_out_wg_data[277], dat_out_wg_data[278], dat_out_wg_data[279] };
  assign dat_out_wg_mask_int8[35] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18385" *) { dat_out_wg_data[280], dat_out_wg_data[281], dat_out_wg_data[282], dat_out_wg_data[283], dat_out_wg_data[284], dat_out_wg_data[285], dat_out_wg_data[286], dat_out_wg_data[287] };
  assign dat_out_wg_mask_int8[36] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18385" *) { dat_out_wg_data[288], dat_out_wg_data[289], dat_out_wg_data[290], dat_out_wg_data[291], dat_out_wg_data[292], dat_out_wg_data[293], dat_out_wg_data[294], dat_out_wg_data[295] };
  assign dat_out_wg_mask_int8[37] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18385" *) { dat_out_wg_data[296], dat_out_wg_data[297], dat_out_wg_data[298], dat_out_wg_data[299], dat_out_wg_data[300], dat_out_wg_data[301], dat_out_wg_data[302], dat_out_wg_data[303] };
  assign dat_out_wg_mask_int8[38] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18385" *) { dat_out_wg_data[304], dat_out_wg_data[305], dat_out_wg_data[306], dat_out_wg_data[307], dat_out_wg_data[308], dat_out_wg_data[309], dat_out_wg_data[310], dat_out_wg_data[311] };
  assign dat_out_wg_mask_int8[39] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18385" *) { dat_out_wg_data[312], dat_out_wg_data[313], dat_out_wg_data[314], dat_out_wg_data[315], dat_out_wg_data[316], dat_out_wg_data[317], dat_out_wg_data[318], dat_out_wg_data[319] };
  assign dat_out_wg_mask_int8[24] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18386" *) { dat_out_wg_data[192], dat_out_wg_data[193], dat_out_wg_data[194], dat_out_wg_data[195], dat_out_wg_data[196], dat_out_wg_data[197], dat_out_wg_data[198], dat_out_wg_data[199] };
  assign dat_out_wg_mask_int8[25] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18386" *) { dat_out_wg_data[200], dat_out_wg_data[201], dat_out_wg_data[202], dat_out_wg_data[203], dat_out_wg_data[204], dat_out_wg_data[205], dat_out_wg_data[206], dat_out_wg_data[207] };
  assign dat_out_wg_mask_int8[26] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18386" *) { dat_out_wg_data[208], dat_out_wg_data[209], dat_out_wg_data[210], dat_out_wg_data[211], dat_out_wg_data[212], dat_out_wg_data[213], dat_out_wg_data[214], dat_out_wg_data[215] };
  assign dat_out_wg_mask_int8[27] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18386" *) { dat_out_wg_data[216], dat_out_wg_data[217], dat_out_wg_data[218], dat_out_wg_data[219], dat_out_wg_data[220], dat_out_wg_data[221], dat_out_wg_data[222], dat_out_wg_data[223] };
  assign dat_out_wg_mask_int8[28] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18386" *) { dat_out_wg_data[224], dat_out_wg_data[225], dat_out_wg_data[226], dat_out_wg_data[227], dat_out_wg_data[228], dat_out_wg_data[229], dat_out_wg_data[230], dat_out_wg_data[231] };
  assign dat_out_wg_mask_int8[29] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18386" *) { dat_out_wg_data[232], dat_out_wg_data[233], dat_out_wg_data[234], dat_out_wg_data[235], dat_out_wg_data[236], dat_out_wg_data[237], dat_out_wg_data[238], dat_out_wg_data[239] };
  assign dat_out_wg_mask_int8[30] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18386" *) { dat_out_wg_data[240], dat_out_wg_data[241], dat_out_wg_data[242], dat_out_wg_data[243], dat_out_wg_data[244], dat_out_wg_data[245], dat_out_wg_data[246], dat_out_wg_data[247] };
  assign dat_out_wg_mask_int8[31] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18386" *) { dat_out_wg_data[248], dat_out_wg_data[249], dat_out_wg_data[250], dat_out_wg_data[251], dat_out_wg_data[252], dat_out_wg_data[253], dat_out_wg_data[254], dat_out_wg_data[255] };
  assign dat_out_wg_mask_int8[16] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18387" *) { dat_out_wg_data[128], dat_out_wg_data[129], dat_out_wg_data[130], dat_out_wg_data[131], dat_out_wg_data[132], dat_out_wg_data[133], dat_out_wg_data[134], dat_out_wg_data[135] };
  assign dat_out_wg_mask_int8[17] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18387" *) { dat_out_wg_data[136], dat_out_wg_data[137], dat_out_wg_data[138], dat_out_wg_data[139], dat_out_wg_data[140], dat_out_wg_data[141], dat_out_wg_data[142], dat_out_wg_data[143] };
  assign dat_out_wg_mask_int8[18] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18387" *) { dat_out_wg_data[144], dat_out_wg_data[145], dat_out_wg_data[146], dat_out_wg_data[147], dat_out_wg_data[148], dat_out_wg_data[149], dat_out_wg_data[150], dat_out_wg_data[151] };
  assign dat_out_wg_mask_int8[19] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18387" *) { dat_out_wg_data[152], dat_out_wg_data[153], dat_out_wg_data[154], dat_out_wg_data[155], dat_out_wg_data[156], dat_out_wg_data[157], dat_out_wg_data[158], dat_out_wg_data[159] };
  assign dat_out_wg_mask_int8[20] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18387" *) { dat_out_wg_data[160], dat_out_wg_data[161], dat_out_wg_data[162], dat_out_wg_data[163], dat_out_wg_data[164], dat_out_wg_data[165], dat_out_wg_data[166], dat_out_wg_data[167] };
  assign dat_out_wg_mask_int8[21] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18387" *) { dat_out_wg_data[168], dat_out_wg_data[169], dat_out_wg_data[170], dat_out_wg_data[171], dat_out_wg_data[172], dat_out_wg_data[173], dat_out_wg_data[174], dat_out_wg_data[175] };
  assign dat_out_wg_mask_int8[22] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18387" *) { dat_out_wg_data[176], dat_out_wg_data[177], dat_out_wg_data[178], dat_out_wg_data[179], dat_out_wg_data[180], dat_out_wg_data[181], dat_out_wg_data[182], dat_out_wg_data[183] };
  assign dat_out_wg_mask_int8[23] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18387" *) { dat_out_wg_data[184], dat_out_wg_data[185], dat_out_wg_data[186], dat_out_wg_data[187], dat_out_wg_data[188], dat_out_wg_data[189], dat_out_wg_data[190], dat_out_wg_data[191] };
  assign dat_out_wg_mask_int8[8] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18388" *) { dat_out_wg_data[64], dat_out_wg_data[65], dat_out_wg_data[66], dat_out_wg_data[67], dat_out_wg_data[68], dat_out_wg_data[69], dat_out_wg_data[70], dat_out_wg_data[71] };
  assign dat_out_wg_mask_int8[9] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18388" *) { dat_out_wg_data[72], dat_out_wg_data[73], dat_out_wg_data[74], dat_out_wg_data[75], dat_out_wg_data[76], dat_out_wg_data[77], dat_out_wg_data[78], dat_out_wg_data[79] };
  assign dat_out_wg_mask_int8[10] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18388" *) { dat_out_wg_data[80], dat_out_wg_data[81], dat_out_wg_data[82], dat_out_wg_data[83], dat_out_wg_data[84], dat_out_wg_data[85], dat_out_wg_data[86], dat_out_wg_data[87] };
  assign dat_out_wg_mask_int8[11] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18388" *) { dat_out_wg_data[88], dat_out_wg_data[89], dat_out_wg_data[90], dat_out_wg_data[91], dat_out_wg_data[92], dat_out_wg_data[93], dat_out_wg_data[94], dat_out_wg_data[95] };
  assign dat_out_wg_mask_int8[12] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18388" *) { dat_out_wg_data[96], dat_out_wg_data[97], dat_out_wg_data[98], dat_out_wg_data[99], dat_out_wg_data[100], dat_out_wg_data[101], dat_out_wg_data[102], dat_out_wg_data[103] };
  assign dat_out_wg_mask_int8[13] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18388" *) { dat_out_wg_data[104], dat_out_wg_data[105], dat_out_wg_data[106], dat_out_wg_data[107], dat_out_wg_data[108], dat_out_wg_data[109], dat_out_wg_data[110], dat_out_wg_data[111] };
  assign dat_out_wg_mask_int8[14] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18388" *) { dat_out_wg_data[112], dat_out_wg_data[113], dat_out_wg_data[114], dat_out_wg_data[115], dat_out_wg_data[116], dat_out_wg_data[117], dat_out_wg_data[118], dat_out_wg_data[119] };
  assign dat_out_wg_mask_int8[15] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18388" *) { dat_out_wg_data[120], dat_out_wg_data[121], dat_out_wg_data[122], dat_out_wg_data[123], dat_out_wg_data[124], dat_out_wg_data[125], dat_out_wg_data[126], dat_out_wg_data[127] };
  assign dat_out_wg_mask_int8[0] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18389" *) { dat_out_wg_data[0], dat_out_wg_data[1], dat_out_wg_data[2], dat_out_wg_data[3], dat_out_wg_data[4], dat_out_wg_data[5], dat_out_wg_data[6], dat_out_wg_data[7] };
  assign dat_out_wg_mask_int8[1] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18389" *) { dat_out_wg_data[8], dat_out_wg_data[9], dat_out_wg_data[10], dat_out_wg_data[11], dat_out_wg_data[12], dat_out_wg_data[13], dat_out_wg_data[14], dat_out_wg_data[15] };
  assign dat_out_wg_mask_int8[2] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18389" *) { dat_out_wg_data[16], dat_out_wg_data[17], dat_out_wg_data[18], dat_out_wg_data[19], dat_out_wg_data[20], dat_out_wg_data[21], dat_out_wg_data[22], dat_out_wg_data[23] };
  assign dat_out_wg_mask_int8[3] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18389" *) { dat_out_wg_data[24], dat_out_wg_data[25], dat_out_wg_data[26], dat_out_wg_data[27], dat_out_wg_data[28], dat_out_wg_data[29], dat_out_wg_data[30], dat_out_wg_data[31] };
  assign dat_out_wg_mask_int8[4] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18389" *) { dat_out_wg_data[32], dat_out_wg_data[33], dat_out_wg_data[34], dat_out_wg_data[35], dat_out_wg_data[36], dat_out_wg_data[37], dat_out_wg_data[38], dat_out_wg_data[39] };
  assign dat_out_wg_mask_int8[5] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18389" *) { dat_out_wg_data[40], dat_out_wg_data[41], dat_out_wg_data[42], dat_out_wg_data[43], dat_out_wg_data[44], dat_out_wg_data[45], dat_out_wg_data[46], dat_out_wg_data[47] };
  assign dat_out_wg_mask_int8[6] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18389" *) { dat_out_wg_data[48], dat_out_wg_data[49], dat_out_wg_data[50], dat_out_wg_data[51], dat_out_wg_data[52], dat_out_wg_data[53], dat_out_wg_data[54], dat_out_wg_data[55] };
  assign dat_out_wg_mask_int8[7] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18389" *) { dat_out_wg_data[56], dat_out_wg_data[57], dat_out_wg_data[58], dat_out_wg_data[59], dat_out_wg_data[60], dat_out_wg_data[61], dat_out_wg_data[62], dat_out_wg_data[63] };
  assign dat_out_wg_mask_fp16[113] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18394" *) { dat_out_wg_data[896], dat_out_wg_data[897], dat_out_wg_data[898], dat_out_wg_data[899], dat_out_wg_data[900], dat_out_wg_data[901], dat_out_wg_data[902], dat_out_wg_data[903], dat_out_wg_data[904], dat_out_wg_data[905], dat_out_wg_data[906], dat_out_wg_data[907], dat_out_wg_data[908], dat_out_wg_data[909], dat_out_wg_data[910] };
  assign dat_out_wg_mask_fp16[115] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18394" *) { dat_out_wg_data[912], dat_out_wg_data[913], dat_out_wg_data[914], dat_out_wg_data[915], dat_out_wg_data[916], dat_out_wg_data[917], dat_out_wg_data[918], dat_out_wg_data[919], dat_out_wg_data[920], dat_out_wg_data[921], dat_out_wg_data[922], dat_out_wg_data[923], dat_out_wg_data[924], dat_out_wg_data[925], dat_out_wg_data[926] };
  assign dat_out_wg_mask_fp16[117] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18394" *) { dat_out_wg_data[928], dat_out_wg_data[929], dat_out_wg_data[930], dat_out_wg_data[931], dat_out_wg_data[932], dat_out_wg_data[933], dat_out_wg_data[934], dat_out_wg_data[935], dat_out_wg_data[936], dat_out_wg_data[937], dat_out_wg_data[938], dat_out_wg_data[939], dat_out_wg_data[940], dat_out_wg_data[941], dat_out_wg_data[942] };
  assign dat_out_wg_mask_fp16[119] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18394" *) { dat_out_wg_data[944], dat_out_wg_data[945], dat_out_wg_data[946], dat_out_wg_data[947], dat_out_wg_data[948], dat_out_wg_data[949], dat_out_wg_data[950], dat_out_wg_data[951], dat_out_wg_data[952], dat_out_wg_data[953], dat_out_wg_data[954], dat_out_wg_data[955], dat_out_wg_data[956], dat_out_wg_data[957], dat_out_wg_data[958] };
  assign dat_out_wg_mask_fp16[121] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18394" *) { dat_out_wg_data[960], dat_out_wg_data[961], dat_out_wg_data[962], dat_out_wg_data[963], dat_out_wg_data[964], dat_out_wg_data[965], dat_out_wg_data[966], dat_out_wg_data[967], dat_out_wg_data[968], dat_out_wg_data[969], dat_out_wg_data[970], dat_out_wg_data[971], dat_out_wg_data[972], dat_out_wg_data[973], dat_out_wg_data[974] };
  assign dat_out_wg_mask_fp16[123] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18394" *) { dat_out_wg_data[976], dat_out_wg_data[977], dat_out_wg_data[978], dat_out_wg_data[979], dat_out_wg_data[980], dat_out_wg_data[981], dat_out_wg_data[982], dat_out_wg_data[983], dat_out_wg_data[984], dat_out_wg_data[985], dat_out_wg_data[986], dat_out_wg_data[987], dat_out_wg_data[988], dat_out_wg_data[989], dat_out_wg_data[990] };
  assign dat_out_wg_mask_fp16[125] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18394" *) { dat_out_wg_data[992], dat_out_wg_data[993], dat_out_wg_data[994], dat_out_wg_data[995], dat_out_wg_data[996], dat_out_wg_data[997], dat_out_wg_data[998], dat_out_wg_data[999], dat_out_wg_data[1000], dat_out_wg_data[1001], dat_out_wg_data[1002], dat_out_wg_data[1003], dat_out_wg_data[1004], dat_out_wg_data[1005], dat_out_wg_data[1006] };
  assign dat_out_wg_mask_fp16[127] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18394" *) { dat_out_wg_data[1008], dat_out_wg_data[1009], dat_out_wg_data[1010], dat_out_wg_data[1011], dat_out_wg_data[1012], dat_out_wg_data[1013], dat_out_wg_data[1014], dat_out_wg_data[1015], dat_out_wg_data[1016], dat_out_wg_data[1017], dat_out_wg_data[1018], dat_out_wg_data[1019], dat_out_wg_data[1020], dat_out_wg_data[1021], dat_out_wg_data[1022] };
  assign dat_out_wg_mask_fp16[97] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18395" *) { dat_out_wg_data[768], dat_out_wg_data[769], dat_out_wg_data[770], dat_out_wg_data[771], dat_out_wg_data[772], dat_out_wg_data[773], dat_out_wg_data[774], dat_out_wg_data[775], dat_out_wg_data[776], dat_out_wg_data[777], dat_out_wg_data[778], dat_out_wg_data[779], dat_out_wg_data[780], dat_out_wg_data[781], dat_out_wg_data[782] };
  assign dat_out_wg_mask_fp16[99] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18395" *) { dat_out_wg_data[784], dat_out_wg_data[785], dat_out_wg_data[786], dat_out_wg_data[787], dat_out_wg_data[788], dat_out_wg_data[789], dat_out_wg_data[790], dat_out_wg_data[791], dat_out_wg_data[792], dat_out_wg_data[793], dat_out_wg_data[794], dat_out_wg_data[795], dat_out_wg_data[796], dat_out_wg_data[797], dat_out_wg_data[798] };
  assign dat_out_wg_mask_fp16[101] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18395" *) { dat_out_wg_data[800], dat_out_wg_data[801], dat_out_wg_data[802], dat_out_wg_data[803], dat_out_wg_data[804], dat_out_wg_data[805], dat_out_wg_data[806], dat_out_wg_data[807], dat_out_wg_data[808], dat_out_wg_data[809], dat_out_wg_data[810], dat_out_wg_data[811], dat_out_wg_data[812], dat_out_wg_data[813], dat_out_wg_data[814] };
  assign dat_out_wg_mask_fp16[103] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18395" *) { dat_out_wg_data[816], dat_out_wg_data[817], dat_out_wg_data[818], dat_out_wg_data[819], dat_out_wg_data[820], dat_out_wg_data[821], dat_out_wg_data[822], dat_out_wg_data[823], dat_out_wg_data[824], dat_out_wg_data[825], dat_out_wg_data[826], dat_out_wg_data[827], dat_out_wg_data[828], dat_out_wg_data[829], dat_out_wg_data[830] };
  assign dat_out_wg_mask_fp16[105] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18395" *) { dat_out_wg_data[832], dat_out_wg_data[833], dat_out_wg_data[834], dat_out_wg_data[835], dat_out_wg_data[836], dat_out_wg_data[837], dat_out_wg_data[838], dat_out_wg_data[839], dat_out_wg_data[840], dat_out_wg_data[841], dat_out_wg_data[842], dat_out_wg_data[843], dat_out_wg_data[844], dat_out_wg_data[845], dat_out_wg_data[846] };
  assign dat_out_wg_mask_fp16[107] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18395" *) { dat_out_wg_data[848], dat_out_wg_data[849], dat_out_wg_data[850], dat_out_wg_data[851], dat_out_wg_data[852], dat_out_wg_data[853], dat_out_wg_data[854], dat_out_wg_data[855], dat_out_wg_data[856], dat_out_wg_data[857], dat_out_wg_data[858], dat_out_wg_data[859], dat_out_wg_data[860], dat_out_wg_data[861], dat_out_wg_data[862] };
  assign dat_out_wg_mask_fp16[109] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18395" *) { dat_out_wg_data[864], dat_out_wg_data[865], dat_out_wg_data[866], dat_out_wg_data[867], dat_out_wg_data[868], dat_out_wg_data[869], dat_out_wg_data[870], dat_out_wg_data[871], dat_out_wg_data[872], dat_out_wg_data[873], dat_out_wg_data[874], dat_out_wg_data[875], dat_out_wg_data[876], dat_out_wg_data[877], dat_out_wg_data[878] };
  assign dat_out_wg_mask_fp16[111] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18395" *) { dat_out_wg_data[880], dat_out_wg_data[881], dat_out_wg_data[882], dat_out_wg_data[883], dat_out_wg_data[884], dat_out_wg_data[885], dat_out_wg_data[886], dat_out_wg_data[887], dat_out_wg_data[888], dat_out_wg_data[889], dat_out_wg_data[890], dat_out_wg_data[891], dat_out_wg_data[892], dat_out_wg_data[893], dat_out_wg_data[894] };
  assign dat_out_wg_mask_fp16[81] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18396" *) { dat_out_wg_data[640], dat_out_wg_data[641], dat_out_wg_data[642], dat_out_wg_data[643], dat_out_wg_data[644], dat_out_wg_data[645], dat_out_wg_data[646], dat_out_wg_data[647], dat_out_wg_data[648], dat_out_wg_data[649], dat_out_wg_data[650], dat_out_wg_data[651], dat_out_wg_data[652], dat_out_wg_data[653], dat_out_wg_data[654] };
  assign dat_out_wg_mask_fp16[83] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18396" *) { dat_out_wg_data[656], dat_out_wg_data[657], dat_out_wg_data[658], dat_out_wg_data[659], dat_out_wg_data[660], dat_out_wg_data[661], dat_out_wg_data[662], dat_out_wg_data[663], dat_out_wg_data[664], dat_out_wg_data[665], dat_out_wg_data[666], dat_out_wg_data[667], dat_out_wg_data[668], dat_out_wg_data[669], dat_out_wg_data[670] };
  assign dat_out_wg_mask_fp16[85] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18396" *) { dat_out_wg_data[672], dat_out_wg_data[673], dat_out_wg_data[674], dat_out_wg_data[675], dat_out_wg_data[676], dat_out_wg_data[677], dat_out_wg_data[678], dat_out_wg_data[679], dat_out_wg_data[680], dat_out_wg_data[681], dat_out_wg_data[682], dat_out_wg_data[683], dat_out_wg_data[684], dat_out_wg_data[685], dat_out_wg_data[686] };
  assign dat_out_wg_mask_fp16[87] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18396" *) { dat_out_wg_data[688], dat_out_wg_data[689], dat_out_wg_data[690], dat_out_wg_data[691], dat_out_wg_data[692], dat_out_wg_data[693], dat_out_wg_data[694], dat_out_wg_data[695], dat_out_wg_data[696], dat_out_wg_data[697], dat_out_wg_data[698], dat_out_wg_data[699], dat_out_wg_data[700], dat_out_wg_data[701], dat_out_wg_data[702] };
  assign dat_out_wg_mask_fp16[89] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18396" *) { dat_out_wg_data[704], dat_out_wg_data[705], dat_out_wg_data[706], dat_out_wg_data[707], dat_out_wg_data[708], dat_out_wg_data[709], dat_out_wg_data[710], dat_out_wg_data[711], dat_out_wg_data[712], dat_out_wg_data[713], dat_out_wg_data[714], dat_out_wg_data[715], dat_out_wg_data[716], dat_out_wg_data[717], dat_out_wg_data[718] };
  assign dat_out_wg_mask_fp16[91] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18396" *) { dat_out_wg_data[720], dat_out_wg_data[721], dat_out_wg_data[722], dat_out_wg_data[723], dat_out_wg_data[724], dat_out_wg_data[725], dat_out_wg_data[726], dat_out_wg_data[727], dat_out_wg_data[728], dat_out_wg_data[729], dat_out_wg_data[730], dat_out_wg_data[731], dat_out_wg_data[732], dat_out_wg_data[733], dat_out_wg_data[734] };
  assign dat_out_wg_mask_fp16[93] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18396" *) { dat_out_wg_data[736], dat_out_wg_data[737], dat_out_wg_data[738], dat_out_wg_data[739], dat_out_wg_data[740], dat_out_wg_data[741], dat_out_wg_data[742], dat_out_wg_data[743], dat_out_wg_data[744], dat_out_wg_data[745], dat_out_wg_data[746], dat_out_wg_data[747], dat_out_wg_data[748], dat_out_wg_data[749], dat_out_wg_data[750] };
  assign dat_out_wg_mask_fp16[95] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18396" *) { dat_out_wg_data[752], dat_out_wg_data[753], dat_out_wg_data[754], dat_out_wg_data[755], dat_out_wg_data[756], dat_out_wg_data[757], dat_out_wg_data[758], dat_out_wg_data[759], dat_out_wg_data[760], dat_out_wg_data[761], dat_out_wg_data[762], dat_out_wg_data[763], dat_out_wg_data[764], dat_out_wg_data[765], dat_out_wg_data[766] };
  assign dat_out_wg_mask_fp16[65] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18397" *) { dat_out_wg_data[512], dat_out_wg_data[513], dat_out_wg_data[514], dat_out_wg_data[515], dat_out_wg_data[516], dat_out_wg_data[517], dat_out_wg_data[518], dat_out_wg_data[519], dat_out_wg_data[520], dat_out_wg_data[521], dat_out_wg_data[522], dat_out_wg_data[523], dat_out_wg_data[524], dat_out_wg_data[525], dat_out_wg_data[526] };
  assign dat_out_wg_mask_fp16[67] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18397" *) { dat_out_wg_data[528], dat_out_wg_data[529], dat_out_wg_data[530], dat_out_wg_data[531], dat_out_wg_data[532], dat_out_wg_data[533], dat_out_wg_data[534], dat_out_wg_data[535], dat_out_wg_data[536], dat_out_wg_data[537], dat_out_wg_data[538], dat_out_wg_data[539], dat_out_wg_data[540], dat_out_wg_data[541], dat_out_wg_data[542] };
  assign dat_out_wg_mask_fp16[69] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18397" *) { dat_out_wg_data[544], dat_out_wg_data[545], dat_out_wg_data[546], dat_out_wg_data[547], dat_out_wg_data[548], dat_out_wg_data[549], dat_out_wg_data[550], dat_out_wg_data[551], dat_out_wg_data[552], dat_out_wg_data[553], dat_out_wg_data[554], dat_out_wg_data[555], dat_out_wg_data[556], dat_out_wg_data[557], dat_out_wg_data[558] };
  assign dat_out_wg_mask_fp16[71] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18397" *) { dat_out_wg_data[560], dat_out_wg_data[561], dat_out_wg_data[562], dat_out_wg_data[563], dat_out_wg_data[564], dat_out_wg_data[565], dat_out_wg_data[566], dat_out_wg_data[567], dat_out_wg_data[568], dat_out_wg_data[569], dat_out_wg_data[570], dat_out_wg_data[571], dat_out_wg_data[572], dat_out_wg_data[573], dat_out_wg_data[574] };
  assign dat_out_wg_mask_fp16[73] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18397" *) { dat_out_wg_data[576], dat_out_wg_data[577], dat_out_wg_data[578], dat_out_wg_data[579], dat_out_wg_data[580], dat_out_wg_data[581], dat_out_wg_data[582], dat_out_wg_data[583], dat_out_wg_data[584], dat_out_wg_data[585], dat_out_wg_data[586], dat_out_wg_data[587], dat_out_wg_data[588], dat_out_wg_data[589], dat_out_wg_data[590] };
  assign dat_out_wg_mask_fp16[75] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18397" *) { dat_out_wg_data[592], dat_out_wg_data[593], dat_out_wg_data[594], dat_out_wg_data[595], dat_out_wg_data[596], dat_out_wg_data[597], dat_out_wg_data[598], dat_out_wg_data[599], dat_out_wg_data[600], dat_out_wg_data[601], dat_out_wg_data[602], dat_out_wg_data[603], dat_out_wg_data[604], dat_out_wg_data[605], dat_out_wg_data[606] };
  assign dat_out_wg_mask_fp16[77] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18397" *) { dat_out_wg_data[608], dat_out_wg_data[609], dat_out_wg_data[610], dat_out_wg_data[611], dat_out_wg_data[612], dat_out_wg_data[613], dat_out_wg_data[614], dat_out_wg_data[615], dat_out_wg_data[616], dat_out_wg_data[617], dat_out_wg_data[618], dat_out_wg_data[619], dat_out_wg_data[620], dat_out_wg_data[621], dat_out_wg_data[622] };
  assign dat_out_wg_mask_fp16[79] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18397" *) { dat_out_wg_data[624], dat_out_wg_data[625], dat_out_wg_data[626], dat_out_wg_data[627], dat_out_wg_data[628], dat_out_wg_data[629], dat_out_wg_data[630], dat_out_wg_data[631], dat_out_wg_data[632], dat_out_wg_data[633], dat_out_wg_data[634], dat_out_wg_data[635], dat_out_wg_data[636], dat_out_wg_data[637], dat_out_wg_data[638] };
  assign dat_out_wg_mask_fp16[49] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18398" *) { dat_out_wg_data[384], dat_out_wg_data[385], dat_out_wg_data[386], dat_out_wg_data[387], dat_out_wg_data[388], dat_out_wg_data[389], dat_out_wg_data[390], dat_out_wg_data[391], dat_out_wg_data[392], dat_out_wg_data[393], dat_out_wg_data[394], dat_out_wg_data[395], dat_out_wg_data[396], dat_out_wg_data[397], dat_out_wg_data[398] };
  assign dat_out_wg_mask_fp16[51] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18398" *) { dat_out_wg_data[400], dat_out_wg_data[401], dat_out_wg_data[402], dat_out_wg_data[403], dat_out_wg_data[404], dat_out_wg_data[405], dat_out_wg_data[406], dat_out_wg_data[407], dat_out_wg_data[408], dat_out_wg_data[409], dat_out_wg_data[410], dat_out_wg_data[411], dat_out_wg_data[412], dat_out_wg_data[413], dat_out_wg_data[414] };
  assign dat_out_wg_mask_fp16[53] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18398" *) { dat_out_wg_data[416], dat_out_wg_data[417], dat_out_wg_data[418], dat_out_wg_data[419], dat_out_wg_data[420], dat_out_wg_data[421], dat_out_wg_data[422], dat_out_wg_data[423], dat_out_wg_data[424], dat_out_wg_data[425], dat_out_wg_data[426], dat_out_wg_data[427], dat_out_wg_data[428], dat_out_wg_data[429], dat_out_wg_data[430] };
  assign dat_out_wg_mask_fp16[55] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18398" *) { dat_out_wg_data[432], dat_out_wg_data[433], dat_out_wg_data[434], dat_out_wg_data[435], dat_out_wg_data[436], dat_out_wg_data[437], dat_out_wg_data[438], dat_out_wg_data[439], dat_out_wg_data[440], dat_out_wg_data[441], dat_out_wg_data[442], dat_out_wg_data[443], dat_out_wg_data[444], dat_out_wg_data[445], dat_out_wg_data[446] };
  assign dat_out_wg_mask_fp16[57] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18398" *) { dat_out_wg_data[448], dat_out_wg_data[449], dat_out_wg_data[450], dat_out_wg_data[451], dat_out_wg_data[452], dat_out_wg_data[453], dat_out_wg_data[454], dat_out_wg_data[455], dat_out_wg_data[456], dat_out_wg_data[457], dat_out_wg_data[458], dat_out_wg_data[459], dat_out_wg_data[460], dat_out_wg_data[461], dat_out_wg_data[462] };
  assign dat_out_wg_mask_fp16[59] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18398" *) { dat_out_wg_data[464], dat_out_wg_data[465], dat_out_wg_data[466], dat_out_wg_data[467], dat_out_wg_data[468], dat_out_wg_data[469], dat_out_wg_data[470], dat_out_wg_data[471], dat_out_wg_data[472], dat_out_wg_data[473], dat_out_wg_data[474], dat_out_wg_data[475], dat_out_wg_data[476], dat_out_wg_data[477], dat_out_wg_data[478] };
  assign dat_out_wg_mask_fp16[61] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18398" *) { dat_out_wg_data[480], dat_out_wg_data[481], dat_out_wg_data[482], dat_out_wg_data[483], dat_out_wg_data[484], dat_out_wg_data[485], dat_out_wg_data[486], dat_out_wg_data[487], dat_out_wg_data[488], dat_out_wg_data[489], dat_out_wg_data[490], dat_out_wg_data[491], dat_out_wg_data[492], dat_out_wg_data[493], dat_out_wg_data[494] };
  assign dat_out_wg_mask_fp16[63] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18398" *) { dat_out_wg_data[496], dat_out_wg_data[497], dat_out_wg_data[498], dat_out_wg_data[499], dat_out_wg_data[500], dat_out_wg_data[501], dat_out_wg_data[502], dat_out_wg_data[503], dat_out_wg_data[504], dat_out_wg_data[505], dat_out_wg_data[506], dat_out_wg_data[507], dat_out_wg_data[508], dat_out_wg_data[509], dat_out_wg_data[510] };
  assign dat_out_wg_mask_fp16[33] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18399" *) { dat_out_wg_data[256], dat_out_wg_data[257], dat_out_wg_data[258], dat_out_wg_data[259], dat_out_wg_data[260], dat_out_wg_data[261], dat_out_wg_data[262], dat_out_wg_data[263], dat_out_wg_data[264], dat_out_wg_data[265], dat_out_wg_data[266], dat_out_wg_data[267], dat_out_wg_data[268], dat_out_wg_data[269], dat_out_wg_data[270] };
  assign dat_out_wg_mask_fp16[35] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18399" *) { dat_out_wg_data[272], dat_out_wg_data[273], dat_out_wg_data[274], dat_out_wg_data[275], dat_out_wg_data[276], dat_out_wg_data[277], dat_out_wg_data[278], dat_out_wg_data[279], dat_out_wg_data[280], dat_out_wg_data[281], dat_out_wg_data[282], dat_out_wg_data[283], dat_out_wg_data[284], dat_out_wg_data[285], dat_out_wg_data[286] };
  assign dat_out_wg_mask_fp16[37] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18399" *) { dat_out_wg_data[288], dat_out_wg_data[289], dat_out_wg_data[290], dat_out_wg_data[291], dat_out_wg_data[292], dat_out_wg_data[293], dat_out_wg_data[294], dat_out_wg_data[295], dat_out_wg_data[296], dat_out_wg_data[297], dat_out_wg_data[298], dat_out_wg_data[299], dat_out_wg_data[300], dat_out_wg_data[301], dat_out_wg_data[302] };
  assign dat_out_wg_mask_fp16[39] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18399" *) { dat_out_wg_data[304], dat_out_wg_data[305], dat_out_wg_data[306], dat_out_wg_data[307], dat_out_wg_data[308], dat_out_wg_data[309], dat_out_wg_data[310], dat_out_wg_data[311], dat_out_wg_data[312], dat_out_wg_data[313], dat_out_wg_data[314], dat_out_wg_data[315], dat_out_wg_data[316], dat_out_wg_data[317], dat_out_wg_data[318] };
  assign dat_out_wg_mask_fp16[41] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18399" *) { dat_out_wg_data[320], dat_out_wg_data[321], dat_out_wg_data[322], dat_out_wg_data[323], dat_out_wg_data[324], dat_out_wg_data[325], dat_out_wg_data[326], dat_out_wg_data[327], dat_out_wg_data[328], dat_out_wg_data[329], dat_out_wg_data[330], dat_out_wg_data[331], dat_out_wg_data[332], dat_out_wg_data[333], dat_out_wg_data[334] };
  assign dat_out_wg_mask_fp16[43] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18399" *) { dat_out_wg_data[336], dat_out_wg_data[337], dat_out_wg_data[338], dat_out_wg_data[339], dat_out_wg_data[340], dat_out_wg_data[341], dat_out_wg_data[342], dat_out_wg_data[343], dat_out_wg_data[344], dat_out_wg_data[345], dat_out_wg_data[346], dat_out_wg_data[347], dat_out_wg_data[348], dat_out_wg_data[349], dat_out_wg_data[350] };
  assign dat_out_wg_mask_fp16[45] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18399" *) { dat_out_wg_data[352], dat_out_wg_data[353], dat_out_wg_data[354], dat_out_wg_data[355], dat_out_wg_data[356], dat_out_wg_data[357], dat_out_wg_data[358], dat_out_wg_data[359], dat_out_wg_data[360], dat_out_wg_data[361], dat_out_wg_data[362], dat_out_wg_data[363], dat_out_wg_data[364], dat_out_wg_data[365], dat_out_wg_data[366] };
  assign dat_out_wg_mask_fp16[47] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18399" *) { dat_out_wg_data[368], dat_out_wg_data[369], dat_out_wg_data[370], dat_out_wg_data[371], dat_out_wg_data[372], dat_out_wg_data[373], dat_out_wg_data[374], dat_out_wg_data[375], dat_out_wg_data[376], dat_out_wg_data[377], dat_out_wg_data[378], dat_out_wg_data[379], dat_out_wg_data[380], dat_out_wg_data[381], dat_out_wg_data[382] };
  assign dat_out_wg_mask_fp16[17] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18400" *) { dat_out_wg_data[128], dat_out_wg_data[129], dat_out_wg_data[130], dat_out_wg_data[131], dat_out_wg_data[132], dat_out_wg_data[133], dat_out_wg_data[134], dat_out_wg_data[135], dat_out_wg_data[136], dat_out_wg_data[137], dat_out_wg_data[138], dat_out_wg_data[139], dat_out_wg_data[140], dat_out_wg_data[141], dat_out_wg_data[142] };
  assign dat_out_wg_mask_fp16[19] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18400" *) { dat_out_wg_data[144], dat_out_wg_data[145], dat_out_wg_data[146], dat_out_wg_data[147], dat_out_wg_data[148], dat_out_wg_data[149], dat_out_wg_data[150], dat_out_wg_data[151], dat_out_wg_data[152], dat_out_wg_data[153], dat_out_wg_data[154], dat_out_wg_data[155], dat_out_wg_data[156], dat_out_wg_data[157], dat_out_wg_data[158] };
  assign dat_out_wg_mask_fp16[21] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18400" *) { dat_out_wg_data[160], dat_out_wg_data[161], dat_out_wg_data[162], dat_out_wg_data[163], dat_out_wg_data[164], dat_out_wg_data[165], dat_out_wg_data[166], dat_out_wg_data[167], dat_out_wg_data[168], dat_out_wg_data[169], dat_out_wg_data[170], dat_out_wg_data[171], dat_out_wg_data[172], dat_out_wg_data[173], dat_out_wg_data[174] };
  assign dat_out_wg_mask_fp16[23] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18400" *) { dat_out_wg_data[176], dat_out_wg_data[177], dat_out_wg_data[178], dat_out_wg_data[179], dat_out_wg_data[180], dat_out_wg_data[181], dat_out_wg_data[182], dat_out_wg_data[183], dat_out_wg_data[184], dat_out_wg_data[185], dat_out_wg_data[186], dat_out_wg_data[187], dat_out_wg_data[188], dat_out_wg_data[189], dat_out_wg_data[190] };
  assign dat_out_wg_mask_fp16[25] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18400" *) { dat_out_wg_data[192], dat_out_wg_data[193], dat_out_wg_data[194], dat_out_wg_data[195], dat_out_wg_data[196], dat_out_wg_data[197], dat_out_wg_data[198], dat_out_wg_data[199], dat_out_wg_data[200], dat_out_wg_data[201], dat_out_wg_data[202], dat_out_wg_data[203], dat_out_wg_data[204], dat_out_wg_data[205], dat_out_wg_data[206] };
  assign dat_out_wg_mask_fp16[27] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18400" *) { dat_out_wg_data[208], dat_out_wg_data[209], dat_out_wg_data[210], dat_out_wg_data[211], dat_out_wg_data[212], dat_out_wg_data[213], dat_out_wg_data[214], dat_out_wg_data[215], dat_out_wg_data[216], dat_out_wg_data[217], dat_out_wg_data[218], dat_out_wg_data[219], dat_out_wg_data[220], dat_out_wg_data[221], dat_out_wg_data[222] };
  assign dat_out_wg_mask_fp16[29] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18400" *) { dat_out_wg_data[224], dat_out_wg_data[225], dat_out_wg_data[226], dat_out_wg_data[227], dat_out_wg_data[228], dat_out_wg_data[229], dat_out_wg_data[230], dat_out_wg_data[231], dat_out_wg_data[232], dat_out_wg_data[233], dat_out_wg_data[234], dat_out_wg_data[235], dat_out_wg_data[236], dat_out_wg_data[237], dat_out_wg_data[238] };
  assign dat_out_wg_mask_fp16[31] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18400" *) { dat_out_wg_data[240], dat_out_wg_data[241], dat_out_wg_data[242], dat_out_wg_data[243], dat_out_wg_data[244], dat_out_wg_data[245], dat_out_wg_data[246], dat_out_wg_data[247], dat_out_wg_data[248], dat_out_wg_data[249], dat_out_wg_data[250], dat_out_wg_data[251], dat_out_wg_data[252], dat_out_wg_data[253], dat_out_wg_data[254] };
  assign dat_out_wg_mask_fp16[1] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18401" *) { dat_out_wg_data[0], dat_out_wg_data[1], dat_out_wg_data[2], dat_out_wg_data[3], dat_out_wg_data[4], dat_out_wg_data[5], dat_out_wg_data[6], dat_out_wg_data[7], dat_out_wg_data[8], dat_out_wg_data[9], dat_out_wg_data[10], dat_out_wg_data[11], dat_out_wg_data[12], dat_out_wg_data[13], dat_out_wg_data[14] };
  assign dat_out_wg_mask_fp16[3] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18401" *) { dat_out_wg_data[16], dat_out_wg_data[17], dat_out_wg_data[18], dat_out_wg_data[19], dat_out_wg_data[20], dat_out_wg_data[21], dat_out_wg_data[22], dat_out_wg_data[23], dat_out_wg_data[24], dat_out_wg_data[25], dat_out_wg_data[26], dat_out_wg_data[27], dat_out_wg_data[28], dat_out_wg_data[29], dat_out_wg_data[30] };
  assign dat_out_wg_mask_fp16[5] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18401" *) { dat_out_wg_data[32], dat_out_wg_data[33], dat_out_wg_data[34], dat_out_wg_data[35], dat_out_wg_data[36], dat_out_wg_data[37], dat_out_wg_data[38], dat_out_wg_data[39], dat_out_wg_data[40], dat_out_wg_data[41], dat_out_wg_data[42], dat_out_wg_data[43], dat_out_wg_data[44], dat_out_wg_data[45], dat_out_wg_data[46] };
  assign dat_out_wg_mask_fp16[7] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18401" *) { dat_out_wg_data[48], dat_out_wg_data[49], dat_out_wg_data[50], dat_out_wg_data[51], dat_out_wg_data[52], dat_out_wg_data[53], dat_out_wg_data[54], dat_out_wg_data[55], dat_out_wg_data[56], dat_out_wg_data[57], dat_out_wg_data[58], dat_out_wg_data[59], dat_out_wg_data[60], dat_out_wg_data[61], dat_out_wg_data[62] };
  assign dat_out_wg_mask_fp16[9] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18401" *) { dat_out_wg_data[64], dat_out_wg_data[65], dat_out_wg_data[66], dat_out_wg_data[67], dat_out_wg_data[68], dat_out_wg_data[69], dat_out_wg_data[70], dat_out_wg_data[71], dat_out_wg_data[72], dat_out_wg_data[73], dat_out_wg_data[74], dat_out_wg_data[75], dat_out_wg_data[76], dat_out_wg_data[77], dat_out_wg_data[78] };
  assign dat_out_wg_mask_fp16[11] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18401" *) { dat_out_wg_data[80], dat_out_wg_data[81], dat_out_wg_data[82], dat_out_wg_data[83], dat_out_wg_data[84], dat_out_wg_data[85], dat_out_wg_data[86], dat_out_wg_data[87], dat_out_wg_data[88], dat_out_wg_data[89], dat_out_wg_data[90], dat_out_wg_data[91], dat_out_wg_data[92], dat_out_wg_data[93], dat_out_wg_data[94] };
  assign dat_out_wg_mask_fp16[13] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18401" *) { dat_out_wg_data[96], dat_out_wg_data[97], dat_out_wg_data[98], dat_out_wg_data[99], dat_out_wg_data[100], dat_out_wg_data[101], dat_out_wg_data[102], dat_out_wg_data[103], dat_out_wg_data[104], dat_out_wg_data[105], dat_out_wg_data[106], dat_out_wg_data[107], dat_out_wg_data[108], dat_out_wg_data[109], dat_out_wg_data[110] };
  assign dat_out_wg_mask_fp16[15] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18401" *) { dat_out_wg_data[112], dat_out_wg_data[113], dat_out_wg_data[114], dat_out_wg_data[115], dat_out_wg_data[116], dat_out_wg_data[117], dat_out_wg_data[118], dat_out_wg_data[119], dat_out_wg_data[120], dat_out_wg_data[121], dat_out_wg_data[122], dat_out_wg_data[123], dat_out_wg_data[124], dat_out_wg_data[125], dat_out_wg_data[126] };
  assign dat_out_wg_mask_int16[113] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18406" *) { dat_out_wg_data[896], dat_out_wg_data[897], dat_out_wg_data[898], dat_out_wg_data[899], dat_out_wg_data[900], dat_out_wg_data[901], dat_out_wg_data[902], dat_out_wg_data[903], dat_out_wg_data[904], dat_out_wg_data[905], dat_out_wg_data[906], dat_out_wg_data[907], dat_out_wg_data[908], dat_out_wg_data[909], dat_out_wg_data[910], dat_out_wg_data[911] };
  assign dat_out_wg_mask_int16[115] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18406" *) { dat_out_wg_data[912], dat_out_wg_data[913], dat_out_wg_data[914], dat_out_wg_data[915], dat_out_wg_data[916], dat_out_wg_data[917], dat_out_wg_data[918], dat_out_wg_data[919], dat_out_wg_data[920], dat_out_wg_data[921], dat_out_wg_data[922], dat_out_wg_data[923], dat_out_wg_data[924], dat_out_wg_data[925], dat_out_wg_data[926], dat_out_wg_data[927] };
  assign dat_out_wg_mask_int16[117] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18406" *) { dat_out_wg_data[928], dat_out_wg_data[929], dat_out_wg_data[930], dat_out_wg_data[931], dat_out_wg_data[932], dat_out_wg_data[933], dat_out_wg_data[934], dat_out_wg_data[935], dat_out_wg_data[936], dat_out_wg_data[937], dat_out_wg_data[938], dat_out_wg_data[939], dat_out_wg_data[940], dat_out_wg_data[941], dat_out_wg_data[942], dat_out_wg_data[943] };
  assign dat_out_wg_mask_int16[119] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18406" *) { dat_out_wg_data[944], dat_out_wg_data[945], dat_out_wg_data[946], dat_out_wg_data[947], dat_out_wg_data[948], dat_out_wg_data[949], dat_out_wg_data[950], dat_out_wg_data[951], dat_out_wg_data[952], dat_out_wg_data[953], dat_out_wg_data[954], dat_out_wg_data[955], dat_out_wg_data[956], dat_out_wg_data[957], dat_out_wg_data[958], dat_out_wg_data[959] };
  assign dat_out_wg_mask_int16[121] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18406" *) { dat_out_wg_data[960], dat_out_wg_data[961], dat_out_wg_data[962], dat_out_wg_data[963], dat_out_wg_data[964], dat_out_wg_data[965], dat_out_wg_data[966], dat_out_wg_data[967], dat_out_wg_data[968], dat_out_wg_data[969], dat_out_wg_data[970], dat_out_wg_data[971], dat_out_wg_data[972], dat_out_wg_data[973], dat_out_wg_data[974], dat_out_wg_data[975] };
  assign dat_out_wg_mask_int16[123] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18406" *) { dat_out_wg_data[976], dat_out_wg_data[977], dat_out_wg_data[978], dat_out_wg_data[979], dat_out_wg_data[980], dat_out_wg_data[981], dat_out_wg_data[982], dat_out_wg_data[983], dat_out_wg_data[984], dat_out_wg_data[985], dat_out_wg_data[986], dat_out_wg_data[987], dat_out_wg_data[988], dat_out_wg_data[989], dat_out_wg_data[990], dat_out_wg_data[991] };
  assign dat_out_wg_mask_int16[125] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18406" *) { dat_out_wg_data[992], dat_out_wg_data[993], dat_out_wg_data[994], dat_out_wg_data[995], dat_out_wg_data[996], dat_out_wg_data[997], dat_out_wg_data[998], dat_out_wg_data[999], dat_out_wg_data[1000], dat_out_wg_data[1001], dat_out_wg_data[1002], dat_out_wg_data[1003], dat_out_wg_data[1004], dat_out_wg_data[1005], dat_out_wg_data[1006], dat_out_wg_data[1007] };
  assign dat_out_wg_mask_int16[127] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18406" *) { dat_out_wg_data[1008], dat_out_wg_data[1009], dat_out_wg_data[1010], dat_out_wg_data[1011], dat_out_wg_data[1012], dat_out_wg_data[1013], dat_out_wg_data[1014], dat_out_wg_data[1015], dat_out_wg_data[1016], dat_out_wg_data[1017], dat_out_wg_data[1018], dat_out_wg_data[1019], dat_out_wg_data[1020], dat_out_wg_data[1021], dat_out_wg_data[1022], dat_out_wg_data[1023] };
  assign dat_out_wg_mask_int16[97] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18407" *) { dat_out_wg_data[768], dat_out_wg_data[769], dat_out_wg_data[770], dat_out_wg_data[771], dat_out_wg_data[772], dat_out_wg_data[773], dat_out_wg_data[774], dat_out_wg_data[775], dat_out_wg_data[776], dat_out_wg_data[777], dat_out_wg_data[778], dat_out_wg_data[779], dat_out_wg_data[780], dat_out_wg_data[781], dat_out_wg_data[782], dat_out_wg_data[783] };
  assign dat_out_wg_mask_int16[99] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18407" *) { dat_out_wg_data[784], dat_out_wg_data[785], dat_out_wg_data[786], dat_out_wg_data[787], dat_out_wg_data[788], dat_out_wg_data[789], dat_out_wg_data[790], dat_out_wg_data[791], dat_out_wg_data[792], dat_out_wg_data[793], dat_out_wg_data[794], dat_out_wg_data[795], dat_out_wg_data[796], dat_out_wg_data[797], dat_out_wg_data[798], dat_out_wg_data[799] };
  assign dat_out_wg_mask_int16[101] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18407" *) { dat_out_wg_data[800], dat_out_wg_data[801], dat_out_wg_data[802], dat_out_wg_data[803], dat_out_wg_data[804], dat_out_wg_data[805], dat_out_wg_data[806], dat_out_wg_data[807], dat_out_wg_data[808], dat_out_wg_data[809], dat_out_wg_data[810], dat_out_wg_data[811], dat_out_wg_data[812], dat_out_wg_data[813], dat_out_wg_data[814], dat_out_wg_data[815] };
  assign dat_out_wg_mask_int16[103] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18407" *) { dat_out_wg_data[816], dat_out_wg_data[817], dat_out_wg_data[818], dat_out_wg_data[819], dat_out_wg_data[820], dat_out_wg_data[821], dat_out_wg_data[822], dat_out_wg_data[823], dat_out_wg_data[824], dat_out_wg_data[825], dat_out_wg_data[826], dat_out_wg_data[827], dat_out_wg_data[828], dat_out_wg_data[829], dat_out_wg_data[830], dat_out_wg_data[831] };
  assign dat_out_wg_mask_int16[105] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18407" *) { dat_out_wg_data[832], dat_out_wg_data[833], dat_out_wg_data[834], dat_out_wg_data[835], dat_out_wg_data[836], dat_out_wg_data[837], dat_out_wg_data[838], dat_out_wg_data[839], dat_out_wg_data[840], dat_out_wg_data[841], dat_out_wg_data[842], dat_out_wg_data[843], dat_out_wg_data[844], dat_out_wg_data[845], dat_out_wg_data[846], dat_out_wg_data[847] };
  assign dat_out_wg_mask_int16[107] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18407" *) { dat_out_wg_data[848], dat_out_wg_data[849], dat_out_wg_data[850], dat_out_wg_data[851], dat_out_wg_data[852], dat_out_wg_data[853], dat_out_wg_data[854], dat_out_wg_data[855], dat_out_wg_data[856], dat_out_wg_data[857], dat_out_wg_data[858], dat_out_wg_data[859], dat_out_wg_data[860], dat_out_wg_data[861], dat_out_wg_data[862], dat_out_wg_data[863] };
  assign dat_out_wg_mask_int16[109] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18407" *) { dat_out_wg_data[864], dat_out_wg_data[865], dat_out_wg_data[866], dat_out_wg_data[867], dat_out_wg_data[868], dat_out_wg_data[869], dat_out_wg_data[870], dat_out_wg_data[871], dat_out_wg_data[872], dat_out_wg_data[873], dat_out_wg_data[874], dat_out_wg_data[875], dat_out_wg_data[876], dat_out_wg_data[877], dat_out_wg_data[878], dat_out_wg_data[879] };
  assign dat_out_wg_mask_int16[111] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18407" *) { dat_out_wg_data[880], dat_out_wg_data[881], dat_out_wg_data[882], dat_out_wg_data[883], dat_out_wg_data[884], dat_out_wg_data[885], dat_out_wg_data[886], dat_out_wg_data[887], dat_out_wg_data[888], dat_out_wg_data[889], dat_out_wg_data[890], dat_out_wg_data[891], dat_out_wg_data[892], dat_out_wg_data[893], dat_out_wg_data[894], dat_out_wg_data[895] };
  assign dat_out_wg_mask_int16[81] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18408" *) { dat_out_wg_data[640], dat_out_wg_data[641], dat_out_wg_data[642], dat_out_wg_data[643], dat_out_wg_data[644], dat_out_wg_data[645], dat_out_wg_data[646], dat_out_wg_data[647], dat_out_wg_data[648], dat_out_wg_data[649], dat_out_wg_data[650], dat_out_wg_data[651], dat_out_wg_data[652], dat_out_wg_data[653], dat_out_wg_data[654], dat_out_wg_data[655] };
  assign dat_out_wg_mask_int16[83] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18408" *) { dat_out_wg_data[656], dat_out_wg_data[657], dat_out_wg_data[658], dat_out_wg_data[659], dat_out_wg_data[660], dat_out_wg_data[661], dat_out_wg_data[662], dat_out_wg_data[663], dat_out_wg_data[664], dat_out_wg_data[665], dat_out_wg_data[666], dat_out_wg_data[667], dat_out_wg_data[668], dat_out_wg_data[669], dat_out_wg_data[670], dat_out_wg_data[671] };
  assign dat_out_wg_mask_int16[85] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18408" *) { dat_out_wg_data[672], dat_out_wg_data[673], dat_out_wg_data[674], dat_out_wg_data[675], dat_out_wg_data[676], dat_out_wg_data[677], dat_out_wg_data[678], dat_out_wg_data[679], dat_out_wg_data[680], dat_out_wg_data[681], dat_out_wg_data[682], dat_out_wg_data[683], dat_out_wg_data[684], dat_out_wg_data[685], dat_out_wg_data[686], dat_out_wg_data[687] };
  assign dat_out_wg_mask_int16[87] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18408" *) { dat_out_wg_data[688], dat_out_wg_data[689], dat_out_wg_data[690], dat_out_wg_data[691], dat_out_wg_data[692], dat_out_wg_data[693], dat_out_wg_data[694], dat_out_wg_data[695], dat_out_wg_data[696], dat_out_wg_data[697], dat_out_wg_data[698], dat_out_wg_data[699], dat_out_wg_data[700], dat_out_wg_data[701], dat_out_wg_data[702], dat_out_wg_data[703] };
  assign dat_out_wg_mask_int16[89] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18408" *) { dat_out_wg_data[704], dat_out_wg_data[705], dat_out_wg_data[706], dat_out_wg_data[707], dat_out_wg_data[708], dat_out_wg_data[709], dat_out_wg_data[710], dat_out_wg_data[711], dat_out_wg_data[712], dat_out_wg_data[713], dat_out_wg_data[714], dat_out_wg_data[715], dat_out_wg_data[716], dat_out_wg_data[717], dat_out_wg_data[718], dat_out_wg_data[719] };
  assign dat_out_wg_mask_int16[91] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18408" *) { dat_out_wg_data[720], dat_out_wg_data[721], dat_out_wg_data[722], dat_out_wg_data[723], dat_out_wg_data[724], dat_out_wg_data[725], dat_out_wg_data[726], dat_out_wg_data[727], dat_out_wg_data[728], dat_out_wg_data[729], dat_out_wg_data[730], dat_out_wg_data[731], dat_out_wg_data[732], dat_out_wg_data[733], dat_out_wg_data[734], dat_out_wg_data[735] };
  assign dat_out_wg_mask_int16[93] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18408" *) { dat_out_wg_data[736], dat_out_wg_data[737], dat_out_wg_data[738], dat_out_wg_data[739], dat_out_wg_data[740], dat_out_wg_data[741], dat_out_wg_data[742], dat_out_wg_data[743], dat_out_wg_data[744], dat_out_wg_data[745], dat_out_wg_data[746], dat_out_wg_data[747], dat_out_wg_data[748], dat_out_wg_data[749], dat_out_wg_data[750], dat_out_wg_data[751] };
  assign dat_out_wg_mask_int16[95] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18408" *) { dat_out_wg_data[752], dat_out_wg_data[753], dat_out_wg_data[754], dat_out_wg_data[755], dat_out_wg_data[756], dat_out_wg_data[757], dat_out_wg_data[758], dat_out_wg_data[759], dat_out_wg_data[760], dat_out_wg_data[761], dat_out_wg_data[762], dat_out_wg_data[763], dat_out_wg_data[764], dat_out_wg_data[765], dat_out_wg_data[766], dat_out_wg_data[767] };
  assign dat_out_wg_mask_int16[65] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18409" *) { dat_out_wg_data[512], dat_out_wg_data[513], dat_out_wg_data[514], dat_out_wg_data[515], dat_out_wg_data[516], dat_out_wg_data[517], dat_out_wg_data[518], dat_out_wg_data[519], dat_out_wg_data[520], dat_out_wg_data[521], dat_out_wg_data[522], dat_out_wg_data[523], dat_out_wg_data[524], dat_out_wg_data[525], dat_out_wg_data[526], dat_out_wg_data[527] };
  assign dat_out_wg_mask_int16[67] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18409" *) { dat_out_wg_data[528], dat_out_wg_data[529], dat_out_wg_data[530], dat_out_wg_data[531], dat_out_wg_data[532], dat_out_wg_data[533], dat_out_wg_data[534], dat_out_wg_data[535], dat_out_wg_data[536], dat_out_wg_data[537], dat_out_wg_data[538], dat_out_wg_data[539], dat_out_wg_data[540], dat_out_wg_data[541], dat_out_wg_data[542], dat_out_wg_data[543] };
  assign dat_out_wg_mask_int16[69] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18409" *) { dat_out_wg_data[544], dat_out_wg_data[545], dat_out_wg_data[546], dat_out_wg_data[547], dat_out_wg_data[548], dat_out_wg_data[549], dat_out_wg_data[550], dat_out_wg_data[551], dat_out_wg_data[552], dat_out_wg_data[553], dat_out_wg_data[554], dat_out_wg_data[555], dat_out_wg_data[556], dat_out_wg_data[557], dat_out_wg_data[558], dat_out_wg_data[559] };
  assign dat_out_wg_mask_int16[71] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18409" *) { dat_out_wg_data[560], dat_out_wg_data[561], dat_out_wg_data[562], dat_out_wg_data[563], dat_out_wg_data[564], dat_out_wg_data[565], dat_out_wg_data[566], dat_out_wg_data[567], dat_out_wg_data[568], dat_out_wg_data[569], dat_out_wg_data[570], dat_out_wg_data[571], dat_out_wg_data[572], dat_out_wg_data[573], dat_out_wg_data[574], dat_out_wg_data[575] };
  assign dat_out_wg_mask_int16[73] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18409" *) { dat_out_wg_data[576], dat_out_wg_data[577], dat_out_wg_data[578], dat_out_wg_data[579], dat_out_wg_data[580], dat_out_wg_data[581], dat_out_wg_data[582], dat_out_wg_data[583], dat_out_wg_data[584], dat_out_wg_data[585], dat_out_wg_data[586], dat_out_wg_data[587], dat_out_wg_data[588], dat_out_wg_data[589], dat_out_wg_data[590], dat_out_wg_data[591] };
  assign dat_out_wg_mask_int16[75] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18409" *) { dat_out_wg_data[592], dat_out_wg_data[593], dat_out_wg_data[594], dat_out_wg_data[595], dat_out_wg_data[596], dat_out_wg_data[597], dat_out_wg_data[598], dat_out_wg_data[599], dat_out_wg_data[600], dat_out_wg_data[601], dat_out_wg_data[602], dat_out_wg_data[603], dat_out_wg_data[604], dat_out_wg_data[605], dat_out_wg_data[606], dat_out_wg_data[607] };
  assign dat_out_wg_mask_int16[77] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18409" *) { dat_out_wg_data[608], dat_out_wg_data[609], dat_out_wg_data[610], dat_out_wg_data[611], dat_out_wg_data[612], dat_out_wg_data[613], dat_out_wg_data[614], dat_out_wg_data[615], dat_out_wg_data[616], dat_out_wg_data[617], dat_out_wg_data[618], dat_out_wg_data[619], dat_out_wg_data[620], dat_out_wg_data[621], dat_out_wg_data[622], dat_out_wg_data[623] };
  assign dat_out_wg_mask_int16[79] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18409" *) { dat_out_wg_data[624], dat_out_wg_data[625], dat_out_wg_data[626], dat_out_wg_data[627], dat_out_wg_data[628], dat_out_wg_data[629], dat_out_wg_data[630], dat_out_wg_data[631], dat_out_wg_data[632], dat_out_wg_data[633], dat_out_wg_data[634], dat_out_wg_data[635], dat_out_wg_data[636], dat_out_wg_data[637], dat_out_wg_data[638], dat_out_wg_data[639] };
  assign dat_out_wg_mask_int16[49] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18410" *) { dat_out_wg_data[384], dat_out_wg_data[385], dat_out_wg_data[386], dat_out_wg_data[387], dat_out_wg_data[388], dat_out_wg_data[389], dat_out_wg_data[390], dat_out_wg_data[391], dat_out_wg_data[392], dat_out_wg_data[393], dat_out_wg_data[394], dat_out_wg_data[395], dat_out_wg_data[396], dat_out_wg_data[397], dat_out_wg_data[398], dat_out_wg_data[399] };
  assign dat_out_wg_mask_int16[51] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18410" *) { dat_out_wg_data[400], dat_out_wg_data[401], dat_out_wg_data[402], dat_out_wg_data[403], dat_out_wg_data[404], dat_out_wg_data[405], dat_out_wg_data[406], dat_out_wg_data[407], dat_out_wg_data[408], dat_out_wg_data[409], dat_out_wg_data[410], dat_out_wg_data[411], dat_out_wg_data[412], dat_out_wg_data[413], dat_out_wg_data[414], dat_out_wg_data[415] };
  assign dat_out_wg_mask_int16[53] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18410" *) { dat_out_wg_data[416], dat_out_wg_data[417], dat_out_wg_data[418], dat_out_wg_data[419], dat_out_wg_data[420], dat_out_wg_data[421], dat_out_wg_data[422], dat_out_wg_data[423], dat_out_wg_data[424], dat_out_wg_data[425], dat_out_wg_data[426], dat_out_wg_data[427], dat_out_wg_data[428], dat_out_wg_data[429], dat_out_wg_data[430], dat_out_wg_data[431] };
  assign dat_out_wg_mask_int16[55] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18410" *) { dat_out_wg_data[432], dat_out_wg_data[433], dat_out_wg_data[434], dat_out_wg_data[435], dat_out_wg_data[436], dat_out_wg_data[437], dat_out_wg_data[438], dat_out_wg_data[439], dat_out_wg_data[440], dat_out_wg_data[441], dat_out_wg_data[442], dat_out_wg_data[443], dat_out_wg_data[444], dat_out_wg_data[445], dat_out_wg_data[446], dat_out_wg_data[447] };
  assign dat_out_wg_mask_int16[57] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18410" *) { dat_out_wg_data[448], dat_out_wg_data[449], dat_out_wg_data[450], dat_out_wg_data[451], dat_out_wg_data[452], dat_out_wg_data[453], dat_out_wg_data[454], dat_out_wg_data[455], dat_out_wg_data[456], dat_out_wg_data[457], dat_out_wg_data[458], dat_out_wg_data[459], dat_out_wg_data[460], dat_out_wg_data[461], dat_out_wg_data[462], dat_out_wg_data[463] };
  assign dat_out_wg_mask_int16[59] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18410" *) { dat_out_wg_data[464], dat_out_wg_data[465], dat_out_wg_data[466], dat_out_wg_data[467], dat_out_wg_data[468], dat_out_wg_data[469], dat_out_wg_data[470], dat_out_wg_data[471], dat_out_wg_data[472], dat_out_wg_data[473], dat_out_wg_data[474], dat_out_wg_data[475], dat_out_wg_data[476], dat_out_wg_data[477], dat_out_wg_data[478], dat_out_wg_data[479] };
  assign dat_out_wg_mask_int16[61] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18410" *) { dat_out_wg_data[480], dat_out_wg_data[481], dat_out_wg_data[482], dat_out_wg_data[483], dat_out_wg_data[484], dat_out_wg_data[485], dat_out_wg_data[486], dat_out_wg_data[487], dat_out_wg_data[488], dat_out_wg_data[489], dat_out_wg_data[490], dat_out_wg_data[491], dat_out_wg_data[492], dat_out_wg_data[493], dat_out_wg_data[494], dat_out_wg_data[495] };
  assign dat_out_wg_mask_int16[63] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18410" *) { dat_out_wg_data[496], dat_out_wg_data[497], dat_out_wg_data[498], dat_out_wg_data[499], dat_out_wg_data[500], dat_out_wg_data[501], dat_out_wg_data[502], dat_out_wg_data[503], dat_out_wg_data[504], dat_out_wg_data[505], dat_out_wg_data[506], dat_out_wg_data[507], dat_out_wg_data[508], dat_out_wg_data[509], dat_out_wg_data[510], dat_out_wg_data[511] };
  assign dat_out_wg_mask_int16[33] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18411" *) { dat_out_wg_data[256], dat_out_wg_data[257], dat_out_wg_data[258], dat_out_wg_data[259], dat_out_wg_data[260], dat_out_wg_data[261], dat_out_wg_data[262], dat_out_wg_data[263], dat_out_wg_data[264], dat_out_wg_data[265], dat_out_wg_data[266], dat_out_wg_data[267], dat_out_wg_data[268], dat_out_wg_data[269], dat_out_wg_data[270], dat_out_wg_data[271] };
  assign dat_out_wg_mask_int16[35] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18411" *) { dat_out_wg_data[272], dat_out_wg_data[273], dat_out_wg_data[274], dat_out_wg_data[275], dat_out_wg_data[276], dat_out_wg_data[277], dat_out_wg_data[278], dat_out_wg_data[279], dat_out_wg_data[280], dat_out_wg_data[281], dat_out_wg_data[282], dat_out_wg_data[283], dat_out_wg_data[284], dat_out_wg_data[285], dat_out_wg_data[286], dat_out_wg_data[287] };
  assign dat_out_wg_mask_int16[37] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18411" *) { dat_out_wg_data[288], dat_out_wg_data[289], dat_out_wg_data[290], dat_out_wg_data[291], dat_out_wg_data[292], dat_out_wg_data[293], dat_out_wg_data[294], dat_out_wg_data[295], dat_out_wg_data[296], dat_out_wg_data[297], dat_out_wg_data[298], dat_out_wg_data[299], dat_out_wg_data[300], dat_out_wg_data[301], dat_out_wg_data[302], dat_out_wg_data[303] };
  assign dat_out_wg_mask_int16[39] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18411" *) { dat_out_wg_data[304], dat_out_wg_data[305], dat_out_wg_data[306], dat_out_wg_data[307], dat_out_wg_data[308], dat_out_wg_data[309], dat_out_wg_data[310], dat_out_wg_data[311], dat_out_wg_data[312], dat_out_wg_data[313], dat_out_wg_data[314], dat_out_wg_data[315], dat_out_wg_data[316], dat_out_wg_data[317], dat_out_wg_data[318], dat_out_wg_data[319] };
  assign dat_out_wg_mask_int16[41] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18411" *) { dat_out_wg_data[320], dat_out_wg_data[321], dat_out_wg_data[322], dat_out_wg_data[323], dat_out_wg_data[324], dat_out_wg_data[325], dat_out_wg_data[326], dat_out_wg_data[327], dat_out_wg_data[328], dat_out_wg_data[329], dat_out_wg_data[330], dat_out_wg_data[331], dat_out_wg_data[332], dat_out_wg_data[333], dat_out_wg_data[334], dat_out_wg_data[335] };
  assign dat_out_wg_mask_int16[43] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18411" *) { dat_out_wg_data[336], dat_out_wg_data[337], dat_out_wg_data[338], dat_out_wg_data[339], dat_out_wg_data[340], dat_out_wg_data[341], dat_out_wg_data[342], dat_out_wg_data[343], dat_out_wg_data[344], dat_out_wg_data[345], dat_out_wg_data[346], dat_out_wg_data[347], dat_out_wg_data[348], dat_out_wg_data[349], dat_out_wg_data[350], dat_out_wg_data[351] };
  assign dat_out_wg_mask_int16[45] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18411" *) { dat_out_wg_data[352], dat_out_wg_data[353], dat_out_wg_data[354], dat_out_wg_data[355], dat_out_wg_data[356], dat_out_wg_data[357], dat_out_wg_data[358], dat_out_wg_data[359], dat_out_wg_data[360], dat_out_wg_data[361], dat_out_wg_data[362], dat_out_wg_data[363], dat_out_wg_data[364], dat_out_wg_data[365], dat_out_wg_data[366], dat_out_wg_data[367] };
  assign dat_out_wg_mask_int16[47] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18411" *) { dat_out_wg_data[368], dat_out_wg_data[369], dat_out_wg_data[370], dat_out_wg_data[371], dat_out_wg_data[372], dat_out_wg_data[373], dat_out_wg_data[374], dat_out_wg_data[375], dat_out_wg_data[376], dat_out_wg_data[377], dat_out_wg_data[378], dat_out_wg_data[379], dat_out_wg_data[380], dat_out_wg_data[381], dat_out_wg_data[382], dat_out_wg_data[383] };
  assign dat_out_wg_mask_int16[17] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18412" *) { dat_out_wg_data[128], dat_out_wg_data[129], dat_out_wg_data[130], dat_out_wg_data[131], dat_out_wg_data[132], dat_out_wg_data[133], dat_out_wg_data[134], dat_out_wg_data[135], dat_out_wg_data[136], dat_out_wg_data[137], dat_out_wg_data[138], dat_out_wg_data[139], dat_out_wg_data[140], dat_out_wg_data[141], dat_out_wg_data[142], dat_out_wg_data[143] };
  assign dat_out_wg_mask_int16[19] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18412" *) { dat_out_wg_data[144], dat_out_wg_data[145], dat_out_wg_data[146], dat_out_wg_data[147], dat_out_wg_data[148], dat_out_wg_data[149], dat_out_wg_data[150], dat_out_wg_data[151], dat_out_wg_data[152], dat_out_wg_data[153], dat_out_wg_data[154], dat_out_wg_data[155], dat_out_wg_data[156], dat_out_wg_data[157], dat_out_wg_data[158], dat_out_wg_data[159] };
  assign dat_out_wg_mask_int16[21] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18412" *) { dat_out_wg_data[160], dat_out_wg_data[161], dat_out_wg_data[162], dat_out_wg_data[163], dat_out_wg_data[164], dat_out_wg_data[165], dat_out_wg_data[166], dat_out_wg_data[167], dat_out_wg_data[168], dat_out_wg_data[169], dat_out_wg_data[170], dat_out_wg_data[171], dat_out_wg_data[172], dat_out_wg_data[173], dat_out_wg_data[174], dat_out_wg_data[175] };
  assign dat_out_wg_mask_int16[23] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18412" *) { dat_out_wg_data[176], dat_out_wg_data[177], dat_out_wg_data[178], dat_out_wg_data[179], dat_out_wg_data[180], dat_out_wg_data[181], dat_out_wg_data[182], dat_out_wg_data[183], dat_out_wg_data[184], dat_out_wg_data[185], dat_out_wg_data[186], dat_out_wg_data[187], dat_out_wg_data[188], dat_out_wg_data[189], dat_out_wg_data[190], dat_out_wg_data[191] };
  assign dat_out_wg_mask_int16[25] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18412" *) { dat_out_wg_data[192], dat_out_wg_data[193], dat_out_wg_data[194], dat_out_wg_data[195], dat_out_wg_data[196], dat_out_wg_data[197], dat_out_wg_data[198], dat_out_wg_data[199], dat_out_wg_data[200], dat_out_wg_data[201], dat_out_wg_data[202], dat_out_wg_data[203], dat_out_wg_data[204], dat_out_wg_data[205], dat_out_wg_data[206], dat_out_wg_data[207] };
  assign dat_out_wg_mask_int16[27] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18412" *) { dat_out_wg_data[208], dat_out_wg_data[209], dat_out_wg_data[210], dat_out_wg_data[211], dat_out_wg_data[212], dat_out_wg_data[213], dat_out_wg_data[214], dat_out_wg_data[215], dat_out_wg_data[216], dat_out_wg_data[217], dat_out_wg_data[218], dat_out_wg_data[219], dat_out_wg_data[220], dat_out_wg_data[221], dat_out_wg_data[222], dat_out_wg_data[223] };
  assign dat_out_wg_mask_int16[29] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18412" *) { dat_out_wg_data[224], dat_out_wg_data[225], dat_out_wg_data[226], dat_out_wg_data[227], dat_out_wg_data[228], dat_out_wg_data[229], dat_out_wg_data[230], dat_out_wg_data[231], dat_out_wg_data[232], dat_out_wg_data[233], dat_out_wg_data[234], dat_out_wg_data[235], dat_out_wg_data[236], dat_out_wg_data[237], dat_out_wg_data[238], dat_out_wg_data[239] };
  assign dat_out_wg_mask_int16[31] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18412" *) { dat_out_wg_data[240], dat_out_wg_data[241], dat_out_wg_data[242], dat_out_wg_data[243], dat_out_wg_data[244], dat_out_wg_data[245], dat_out_wg_data[246], dat_out_wg_data[247], dat_out_wg_data[248], dat_out_wg_data[249], dat_out_wg_data[250], dat_out_wg_data[251], dat_out_wg_data[252], dat_out_wg_data[253], dat_out_wg_data[254], dat_out_wg_data[255] };
  assign dat_out_wg_mask_int16[1] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18413" *) { dat_out_wg_data[0], dat_out_wg_data[1], dat_out_wg_data[2], dat_out_wg_data[3], dat_out_wg_data[4], dat_out_wg_data[5], dat_out_wg_data[6], dat_out_wg_data[7], dat_out_wg_data[8], dat_out_wg_data[9], dat_out_wg_data[10], dat_out_wg_data[11], dat_out_wg_data[12], dat_out_wg_data[13], dat_out_wg_data[14], dat_out_wg_data[15] };
  assign dat_out_wg_mask_int16[3] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18413" *) { dat_out_wg_data[16], dat_out_wg_data[17], dat_out_wg_data[18], dat_out_wg_data[19], dat_out_wg_data[20], dat_out_wg_data[21], dat_out_wg_data[22], dat_out_wg_data[23], dat_out_wg_data[24], dat_out_wg_data[25], dat_out_wg_data[26], dat_out_wg_data[27], dat_out_wg_data[28], dat_out_wg_data[29], dat_out_wg_data[30], dat_out_wg_data[31] };
  assign dat_out_wg_mask_int16[5] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18413" *) { dat_out_wg_data[32], dat_out_wg_data[33], dat_out_wg_data[34], dat_out_wg_data[35], dat_out_wg_data[36], dat_out_wg_data[37], dat_out_wg_data[38], dat_out_wg_data[39], dat_out_wg_data[40], dat_out_wg_data[41], dat_out_wg_data[42], dat_out_wg_data[43], dat_out_wg_data[44], dat_out_wg_data[45], dat_out_wg_data[46], dat_out_wg_data[47] };
  assign dat_out_wg_mask_int16[7] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18413" *) { dat_out_wg_data[48], dat_out_wg_data[49], dat_out_wg_data[50], dat_out_wg_data[51], dat_out_wg_data[52], dat_out_wg_data[53], dat_out_wg_data[54], dat_out_wg_data[55], dat_out_wg_data[56], dat_out_wg_data[57], dat_out_wg_data[58], dat_out_wg_data[59], dat_out_wg_data[60], dat_out_wg_data[61], dat_out_wg_data[62], dat_out_wg_data[63] };
  assign dat_out_wg_mask_int16[9] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18413" *) { dat_out_wg_data[64], dat_out_wg_data[65], dat_out_wg_data[66], dat_out_wg_data[67], dat_out_wg_data[68], dat_out_wg_data[69], dat_out_wg_data[70], dat_out_wg_data[71], dat_out_wg_data[72], dat_out_wg_data[73], dat_out_wg_data[74], dat_out_wg_data[75], dat_out_wg_data[76], dat_out_wg_data[77], dat_out_wg_data[78], dat_out_wg_data[79] };
  assign dat_out_wg_mask_int16[11] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18413" *) { dat_out_wg_data[80], dat_out_wg_data[81], dat_out_wg_data[82], dat_out_wg_data[83], dat_out_wg_data[84], dat_out_wg_data[85], dat_out_wg_data[86], dat_out_wg_data[87], dat_out_wg_data[88], dat_out_wg_data[89], dat_out_wg_data[90], dat_out_wg_data[91], dat_out_wg_data[92], dat_out_wg_data[93], dat_out_wg_data[94], dat_out_wg_data[95] };
  assign dat_out_wg_mask_int16[13] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18413" *) { dat_out_wg_data[96], dat_out_wg_data[97], dat_out_wg_data[98], dat_out_wg_data[99], dat_out_wg_data[100], dat_out_wg_data[101], dat_out_wg_data[102], dat_out_wg_data[103], dat_out_wg_data[104], dat_out_wg_data[105], dat_out_wg_data[106], dat_out_wg_data[107], dat_out_wg_data[108], dat_out_wg_data[109], dat_out_wg_data[110], dat_out_wg_data[111] };
  assign dat_out_wg_mask_int16[15] = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18413" *) { dat_out_wg_data[112], dat_out_wg_data[113], dat_out_wg_data[114], dat_out_wg_data[115], dat_out_wg_data[116], dat_out_wg_data[117], dat_out_wg_data[118], dat_out_wg_data[119], dat_out_wg_data[120], dat_out_wg_data[121], dat_out_wg_data[122], dat_out_wg_data[123], dat_out_wg_data[124], dat_out_wg_data[125], dat_out_wg_data[126], dat_out_wg_data[127] };
  assign _1160_ = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:7446" *) { last_slices[0], last_slices[1], last_slices[2], last_slices[3], last_slices[4], last_slices[5], last_slices[6], last_slices[7], last_slices[8], last_slices[9], last_slices[10], last_slices[11] };
  assign _1161_ = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:7446" *) { rls_slices[0], rls_slices[1], rls_slices[2], rls_slices[3], rls_slices[4], rls_slices[5], rls_slices[6], rls_slices[7], rls_slices[8], rls_slices[9], rls_slices[10], rls_slices[11] };
  assign _1162_ = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:8728" *) { reg2dp_y_extension[0], reg2dp_y_extension[1] };
  assign _1163_ = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:9100" *) { stripe_cnt[0], stripe_cnt[1], stripe_cnt[2], stripe_cnt[3], stripe_cnt[4], stripe_cnt[5], stripe_cnt[6] };
  assign _1164_ = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:9100" *) { sub_h_cnt[0], sub_h_cnt[1] };
  assign _1165_ = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:9100" *) { batch_cnt[0], batch_cnt[1], batch_cnt[2], batch_cnt[3], batch_cnt[4] };
  assign _1166_ = 128'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111 << (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16271" *) dat_rsp_pd[14:7];
  assign _1167_ = 4'b1001 << (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1989" *) reg2dp_y_extension;
  assign dat_rsp_l0_sft = dat_rsp_l0_sft_in >> (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16087" *) { rsp_sft_cnt_l0[6:0], 3'b000 };
  assign dat_rsp_l1_sft = dat_rsp_l1_sft_in >> (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16088" *) { rsp_sft_cnt_l1[5:0], 3'b000 };
  assign dat_rsp_l2_sft = dat_rsp_l2_sft_in >> (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16089" *) { rsp_sft_cnt_l2[5:0], 3'b000 };
  assign dat_rsp_l3_sft = dat_rsp_l3_sft_in >> (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16090" *) { rsp_sft_cnt_l3[5:0], 3'b000 };
  assign { _1168_[13], _1168_[4:0] } = 1'b0 - (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:10224" *) reg2dp_pad_top;
  assign dat_req_addr_wrap = dat_req_addr_sum[11:0] - (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:12170" *) { data_bank, 8'b00000000 };
  assign rsp_sft_cnt_l0_inc = _0709_ - (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15136" *) rsp_sft_cnt_l0_sub;
  assign rsp_sft_cnt_l1_inc = _0710_ - (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15144" *) rsp_sft_cnt_l1_sub;
  assign rsp_sft_cnt_l2_inc = _0711_ - (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15152" *) rsp_sft_cnt_l2_sub;
  assign rsp_sft_cnt_l3_inc = _0712_ - (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15160" *) rsp_sft_cnt_l3_sub;
  assign { dataout_w_init[12], dataout_w_init[2:0] } = sub_h_cmp_w - (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:2004" *) 1'b1;
  assign _1020_[11:0] = reg2dp_datain_height_ext[11:0] - (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:2134" *) reg2dp_rls_slices;
  assign dat_entry_st_inc_wrap = dat_entry_st_inc[11:0] - (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:6709" *) { data_bank, 8'b00000000 };
  assign { _1169_[13], _1169_[4:0] } = 1'b0 - (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:9608" *) reg2dp_pad_left;
  assign datain_h_cnt_st = reg2dp_conv_mode ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:10224" *) 14'b00000000000000 : { _1168_[13], _1168_[13], _1168_[13], _1168_[13], _1168_[13], _1168_[13], _1168_[13], _1168_[13], _1168_[13], _1168_[4:0] };
  assign _1170_ = is_w_end ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:10247" *) datain_h_cnt_inc : datain_h_cnt;
  assign _1171_ = _0733_ ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:10247" *) datain_h_ori : _1170_;
  assign datain_h_cnt_w = _1123_ ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:10247" *) datain_h_cnt_st : _1171_;
  assign _1172_ = is_winograd_d1[4] ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:10440" *) 1'b0 : dat_conv_req_dummy;
  assign dat_req_dummy = is_img_d1[5] ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:10440" *) dat_img_req_dummy : _1172_;
  assign dat_req_sub_c_w = is_img_d1[7] ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:10465" *) dl_pd[26] : _0741_;
  assign dat_req_sub_w_w = is_winograd_d1[6] ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:10472" *) { 1'b0, _1081_ } : datain_w_cur[1:0];
  assign c_bias_add = _0744_ ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:11331" *) datain_width[11:0] : 12'b000000000000;
  assign _1173_[11:0] = _0745_ ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:11343" *) 12'b000000000000 : _0704_;
  assign c_bias_w = layer_st ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:11343" *) 12'b000000000000 : _1173_[11:0];
  assign h_bias_3_w = layer_st ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:11388" *) 12'b000000000000 : _1019_[11:0];
  assign _1021_[13:0] = _1069_ ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:11407" *) { datain_w_cur[12:0], 1'b0 } : { 1'b0, datain_w_cur[12:0] };
  assign _1022_[13:0] = _1130_ ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:11407" *) { datain_w_cur[11:0], 2'b00 } : _1021_[13:0];
  assign _1023_[13:0] = is_winograd_d1[8] ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:11407" *) datain_w_cnt : _1022_[13:0];
  assign w_bias_int8 = is_img_d1[10] ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:11407" *) { 3'b000, pixel_w_cnt[15:6], 1'b0 } : _1023_[13:0];
  assign _1024_[13:0] = _1131_ ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:11421" *) { datain_w_cur[11:0], 2'b00 } : _1021_[13:0];
  assign _1025_[13:0] = is_winograd_d1[9] ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:11421" *) datain_w_cnt : _1024_[13:0];
  assign w_bias_16 = is_img_d1[11] ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:11421" *) { 2'b00, pixel_w_cnt[15:6], 2'b00 } : _1025_[13:0];
  assign w_bias_w = is_int8_d1[4] ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:11428" *) w_bias_int8 : w_bias_16;
  assign _1174_ = is_dat_req_addr_wrap ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:12180" *) dat_req_addr_wrap : dat_req_addr_sum[11:0];
  assign dat_req_addr_w = _1132_ ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:12180" *) 12'b111111111111 : _1174_;
  assign _1175_ = _1029_ ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:12193" *) dat_req_sub_h_2_addr : dat_req_sub_h_3_addr;
  assign _1176_ = _1028_ ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:12193" *) dat_req_sub_h_1_addr : _1175_;
  assign dat_req_addr_last = _1027_ ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:12193" *) dat_req_sub_h_0_addr : _1176_;
  assign _1177_ = dat_dummy_l0_en ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:14567" *) 1'b1 : dat_l0c0_dummy;
  assign dat_l0c0_dummy_w = dat_l0c0_en ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:14567" *) 1'b0 : _1177_;
  assign _1178_ = dat_dummy_l1_en ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:14570" *) 1'b1 : dat_l1c0_dummy;
  assign dat_l1c0_dummy_w = dat_l1c0_en ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:14570" *) 1'b0 : _1178_;
  assign _1179_ = dat_dummy_l2_en ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:14573" *) 1'b1 : dat_l2c0_dummy;
  assign dat_l2c0_dummy_w = dat_l2c0_en ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:14573" *) 1'b0 : _1179_;
  assign _1180_ = dat_dummy_l3_en ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:14576" *) 1'b1 : dat_l3c0_dummy;
  assign dat_l3c0_dummy_w = dat_l3c0_en ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:14576" *) 1'b0 : _1180_;
  assign _1181_ = dat_l0_set ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:14579" *) dat_l0c0_dummy : dat_l0c1_dummy;
  assign dat_l0c1_dummy_w = dat_l0c1_en ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:14579" *) 1'b0 : _1181_;
  assign _1182_ = _0763_ ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:14582" *) dat_l1c0_dummy : dat_l1c1_dummy;
  assign dat_l1c1_dummy_w = dat_l1c1_en ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:14582" *) 1'b0 : _1182_;
  assign _1183_ = _0764_ ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:14585" *) dat_l2c0_dummy : dat_l2c1_dummy;
  assign dat_l2c1_dummy_w = dat_l2c1_en ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:14585" *) 1'b0 : _1183_;
  assign _1184_ = _0765_ ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:14588" *) dat_l3c0_dummy : dat_l3c1_dummy;
  assign dat_l3c1_dummy_w = dat_l3c1_en ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:14588" *) 1'b0 : _1184_;
  assign rsp_sft_cnt_l0_sub = dat_l0c0_en ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15126" *) 8'b10000000 : 8'b00000000;
  assign rsp_sft_cnt_l1_sub = dat_l1c0_en ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15127" *) 8'b10000000 : 8'b00000000;
  assign rsp_sft_cnt_l2_sub = dat_l2c0_en ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15128" *) 8'b10000000 : 8'b00000000;
  assign rsp_sft_cnt_l3_sub = dat_l3c0_en ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15129" *) 8'b10000000 : 8'b00000000;
  assign _1185_ = dat_dummy_l0_en ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15180" *) _0776_ : rsp_sft_cnt_l0_inc;
  assign _1186_ = _0775_ ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15180" *) 8'b10000000 : _1185_;
  assign _1187_ = _0774_ ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15180" *) 8'b11000000 : _1186_;
  assign _1188_ = _0772_ ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15180" *) rsp_sft_cnt_l0_ori : _1187_;
  assign rsp_sft_cnt_l0_w = layer_st ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15180" *) 8'b10000000 : _1188_;
  assign _1189_ = dat_dummy_l1_en ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15196" *) _0781_ : rsp_sft_cnt_l1_inc;
  assign _1190_ = _0780_ ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15196" *) 8'b10000000 : _1189_;
  assign _1191_ = _0779_ ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15196" *) 8'b11000000 : _1190_;
  assign _1192_ = _0777_ ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15196" *) rsp_sft_cnt_l1_ori : _1191_;
  assign rsp_sft_cnt_l1_w = layer_st ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15196" *) 8'b10000000 : _1192_;
  assign _1193_ = dat_dummy_l2_en ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15212" *) _0786_ : rsp_sft_cnt_l2_inc;
  assign _1194_ = _0785_ ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15212" *) 8'b10000000 : _1193_;
  assign _1195_ = _0784_ ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15212" *) 8'b11000000 : _1194_;
  assign _1196_ = _0782_ ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15212" *) rsp_sft_cnt_l2_ori : _1195_;
  assign rsp_sft_cnt_l2_w = layer_st ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15212" *) 8'b10000000 : _1196_;
  assign _1197_ = dat_dummy_l3_en ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15228" *) _0791_ : rsp_sft_cnt_l3_inc;
  assign _1198_ = _0790_ ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15228" *) 8'b10000000 : _1197_;
  assign _1199_ = _0789_ ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15228" *) 8'b11000000 : _1198_;
  assign _1200_ = _0787_ ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15228" *) rsp_sft_cnt_l3_ori : _1199_;
  assign rsp_sft_cnt_l3_w = layer_st ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15228" *) 8'b10000000 : _1200_;
  assign dat_wg = is_winograd_d1[12] ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15774" *) { dat_l1c0_lo[511:256], dat_l1c1_lo[511:384], dat_l1c0_lo[255:0], dat_l1c1_lo[255:128], dat_l0c0_hi[511:256], dat_l0c1_hi[511:384], dat_l0c0_hi[255:0], dat_l0c1_hi[255:128], dat_l0c0_lo[511:256], dat_l0c1_lo[511:384], dat_l0c0_lo[255:0], dat_l0c1_lo[255:128] } : 2304'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
  assign dat_rsp_pad_value = is_int8_d1[8] ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15901" *) { pad_value[7:0], pad_value[7:0], pad_value[7:0], pad_value[7:0], pad_value[7:0], pad_value[7:0], pad_value[7:0], pad_value[7:0], pad_value[7:0], pad_value[7:0], pad_value[7:0], pad_value[7:0], pad_value[7:0], pad_value[7:0], pad_value[7:0], pad_value[7:0], pad_value[7:0], pad_value[7:0], pad_value[7:0], pad_value[7:0], pad_value[7:0], pad_value[7:0], pad_value[7:0], pad_value[7:0], pad_value[7:0], pad_value[7:0], pad_value[7:0], pad_value[7:0], pad_value[7:0], pad_value[7:0], pad_value[7:0], pad_value[7:0], pad_value[7:0], pad_value[7:0], pad_value[7:0], pad_value[7:0], pad_value[7:0], pad_value[7:0], pad_value[7:0], pad_value[7:0], pad_value[7:0], pad_value[7:0], pad_value[7:0], pad_value[7:0], pad_value[7:0], pad_value[7:0], pad_value[7:0], pad_value[7:0], pad_value[7:0], pad_value[7:0], pad_value[7:0], pad_value[7:0], pad_value[7:0], pad_value[7:0], pad_value[7:0], pad_value[7:0], pad_value[7:0], pad_value[7:0], pad_value[7:0], pad_value[7:0], pad_value[7:0], pad_value[7:0], pad_value[7:0], pad_value[7:0] } : { pad_value, pad_value, pad_value, pad_value, pad_value, pad_value, pad_value, pad_value, pad_value, pad_value, pad_value, pad_value, pad_value, pad_value, pad_value, pad_value, pad_value, pad_value, pad_value, pad_value, pad_value, pad_value, pad_value, pad_value, pad_value, pad_value, pad_value, pad_value, pad_value, pad_value, pad_value, pad_value };
  assign dat_rsp_l0c0_lo = dat_l0c0_dummy ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15918" *) dat_rsp_pad_value : dat_l0c0_lo;
  assign dat_rsp_l0c0_hi = dat_l0c0_dummy ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15919" *) dat_rsp_pad_value : dat_l0c0_hi;
  assign dat_rsp_l1c0_lo = dat_l1c0_dummy ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15920" *) dat_rsp_pad_value : dat_l1c0_lo;
  assign dat_rsp_l1c0_hi = dat_l1c0_dummy ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15921" *) dat_rsp_pad_value : dat_l1c0_hi;
  assign dat_rsp_l2c0_lo = dat_l2c0_dummy ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15922" *) dat_rsp_pad_value : dat_l2c0_lo;
  assign dat_rsp_l2c0_hi = dat_l2c0_dummy ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15923" *) dat_rsp_pad_value : dat_l2c0_hi;
  assign dat_rsp_l3c0_lo = dat_l3c0_dummy ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15924" *) dat_rsp_pad_value : dat_l3c0_lo;
  assign dat_rsp_l3c0_hi = dat_l3c0_dummy ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15925" *) dat_rsp_pad_value : dat_l3c0_hi;
  assign dat_rsp_l0c1_lo = dat_l0c1_dummy ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15942" *) dat_rsp_pad_value : dat_l0c1_lo;
  assign dat_rsp_l0c1_hi = dat_l0c1_dummy ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15943" *) dat_rsp_pad_value : dat_l0c1_hi;
  assign dat_rsp_l1c1_lo = dat_l1c1_dummy ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15944" *) dat_rsp_pad_value : dat_l1c1_lo;
  assign dat_rsp_l1c1_hi = dat_l1c1_dummy ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15945" *) dat_rsp_pad_value : dat_l1c1_hi;
  assign dat_rsp_l2c1_lo = dat_l2c1_dummy ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15946" *) dat_rsp_pad_value : dat_l2c1_lo;
  assign dat_rsp_l2c1_hi = dat_l2c1_dummy ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15947" *) dat_rsp_pad_value : dat_l2c1_hi;
  assign dat_rsp_l3c1_lo = dat_l3c1_dummy ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15948" *) dat_rsp_pad_value : dat_l3c1_lo;
  assign dat_rsp_l3c1_hi = dat_l3c1_dummy ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15949" *) dat_rsp_pad_value : dat_l3c1_hi;
  assign _1201_ = _0836_ ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15967" *) { 768'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, dat_rsp_l0c0_hi[511:256] } : { dat_rsp_l0c0_hi, dat_rsp_l0c0_lo };
  assign _1202_ = _0835_ ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15967" *) { 768'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, dat_rsp_l0c0_hi[255:0] } : _1201_;
  assign _1203_ = _0834_ ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15967" *) { 768'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, dat_rsp_l0c0_lo[511:256] } : _1202_;
  assign _1204_ = _0833_ ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15967" *) { 768'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, dat_rsp_l0c0_lo[255:0] } : _1203_;
  assign _1205_ = _0832_ ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15967" *) { 512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, dat_rsp_l0c0_hi } : _1204_;
  assign _1206_ = _0831_ ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15967" *) { 512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, dat_rsp_l0c0_lo } : _1205_;
  assign dat_rsp_conv_16b = _1144_ ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15967" *) 1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 : _1206_;
  assign _1207_ = _1147_ ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15987" *) dat_rsp_l0c0_hi : dat_rsp_l0c0_lo;
  assign _1208_ = _0836_ ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15987" *) { 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, dat_rsp_l0c0_hi[511:256] } : _1207_;
  assign _1209_ = _0835_ ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15987" *) { 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, dat_rsp_l0c0_hi[255:0] } : _1208_;
  assign _1210_ = _0834_ ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15987" *) { 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, dat_rsp_l0c0_lo[511:256] } : _1209_;
  assign _1211_ = _0833_ ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15987" *) { 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, dat_rsp_l0c0_lo[255:0] } : _1210_;
  assign _1212_ = _0837_ ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15987" *) { 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, dat_rsp_l0c0_hi[255:0] } : _1211_;
  assign dat_rsp_conv_8b = _1146_ ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:15987" *) 512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 : _1212_;
  assign _1213_ = rsp_sft_cnt_l0[7] ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16027" *) { 1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, dat_rsp_l0c0_hi, dat_rsp_l0c0_lo } : { dat_rsp_l0c0_hi, dat_rsp_l0c0_lo, dat_rsp_l0c1_hi, dat_rsp_l0c1_lo };
  assign dat_rsp_l0_sft_in = is_img_d1[27] ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16027" *) _1213_ : 2048'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
  assign _1214_ = rsp_sft_l1_sel_1 ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16043" *) { dat_rsp_l1c0_lo, dat_rsp_l1c1_hi } : { dat_rsp_l1c1_hi, dat_rsp_l1c1_lo };
  assign _1215_ = rsp_sft_l1_sel_2 ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16043" *) { dat_rsp_l1c0_hi, dat_rsp_l1c0_lo } : _1214_;
  assign _1216_ = rsp_sft_l1_sel_3 ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16043" *) { 512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, dat_rsp_l1c0_hi } : _1215_;
  assign dat_rsp_l1_sft_in = is_img_d1[28] ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16043" *) _1216_ : 1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
  assign _1217_ = rsp_sft_l2_sel_1 ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16059" *) { dat_rsp_l2c0_lo, dat_rsp_l2c1_hi } : { dat_rsp_l2c1_hi, dat_rsp_l2c1_lo };
  assign _1218_ = rsp_sft_l2_sel_2 ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16059" *) { dat_rsp_l2c0_hi, dat_rsp_l2c0_lo } : _1217_;
  assign _1219_ = rsp_sft_l2_sel_3 ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16059" *) { 512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, dat_rsp_l2c0_hi } : _1218_;
  assign dat_rsp_l2_sft_in = is_img_d1[29] ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16059" *) _1219_ : 1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
  assign _1220_ = rsp_sft_l3_sel_1 ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16075" *) { dat_rsp_l3c0_lo, dat_rsp_l3c1_hi } : { dat_rsp_l3c1_hi, dat_rsp_l3c1_lo };
  assign _1221_ = rsp_sft_l3_sel_2 ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16075" *) { dat_rsp_l3c0_hi, dat_rsp_l3c0_lo } : _1220_;
  assign _1222_ = rsp_sft_l3_sel_3 ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16075" *) { 512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, dat_rsp_l3c0_hi } : _1221_;
  assign dat_rsp_l3_sft_in = is_img_d1[30] ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16075" *) _1222_ : 1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
  assign _1223_ = _1044_ ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16107" *) { dat_rsp_l1_sft, dat_rsp_l0_sft_d1 } : dat_rsp_l0_sft;
  assign _1224_ = _1043_ ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16107" *) { dat_rsp_l3_sft, dat_rsp_l2_sft_d3, dat_rsp_l1_sft_d3, dat_rsp_l0_sft_d3 } : _1223_;
  assign dat_rsp_img_16b = _1148_ ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16107" *) 1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 : _1224_;
  assign _1225_ = _1046_ ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16124" *) { dat_rsp_l1_sft[255:0], dat_rsp_l0_sft_d1[255:0] } : dat_rsp_l0_sft[511:0];
  assign _1226_ = _1045_ ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16124" *) { dat_rsp_l3_sft[127:0], dat_rsp_l2_sft_d3[127:0], dat_rsp_l1_sft_d3[127:0], dat_rsp_l0_sft_d3[127:0] } : _1225_;
  assign dat_rsp_img_8b = _1149_ ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16124" *) 512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 : _1226_;
  assign dat_rsp_img = is_int8_d1[13] ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16131" *) { dat_rsp_img_8b, dat_rsp_img_8b } : dat_rsp_img_16b;
  assign dat_rsp_cur_h_mask_p1 = _1063_ ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16276" *) 64'b1111111111111111111111111111111111111111111111111111111111111111 : 64'b0000000000000000000000000000000000000000000000000000000000000000;
  assign dat_rsp_cur_h_mask_p2 = _1064_ ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16277" *) 32'd4294967295 : 32'd0;
  assign dat_rsp_cur_h_mask_p3 = _1048_ ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16278" *) 32'd4294967295 : 32'd0;
  assign _1227_ = _1050_ ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16304" *) _0840_ : dat_rsp_ori_mask;
  assign dat_rsp_mask_16b = _1049_ ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16304" *) _0839_ : _1227_;
  assign _1228_ = _1052_ ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16314" *) _0842_ : dat_rsp_ori_mask[63:0];
  assign dat_rsp_mask_8b = _1051_ ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16314" *) _0841_ : _1228_;
  assign dat_out_bypass_data_w = is_img_d1[33] ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16322" *) dat_rsp_img : dat_rsp_conv;
  assign _1229_ = is_fp16_d1[0] ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16371" *) _0844_ : _0845_;
  assign dat_out_bypass_mask_w = is_int8_d1[17] ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16371" *) { 64'b0000000000000000000000000000000000000000000000000000000000000000, _0843_ } : _1229_;
  assign dat_out_pvld_w = is_winograd_d1[17] ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16726" *) dat_out_pvld_l5 : dat_rsp_pvld;
  assign dat_out_flag_w = is_winograd_d1[18] ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:16727" *) dat_out_flag_l5 : dat_rsp_pd[26:18];
  assign dat_out_wg_data = is_int8_d1[19] ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18377" *) { dat_pra_dat_ch3[247:240], dat_pra_dat_ch2[247:240], dat_pra_dat_ch1[247:240], dat_pra_dat_ch0[247:240], dat_pra_dat_ch3[231:224], dat_pra_dat_ch2[231:224], dat_pra_dat_ch1[231:224], dat_pra_dat_ch0[231:224], dat_pra_dat_ch3[215:208], dat_pra_dat_ch2[215:208], dat_pra_dat_ch1[215:208], dat_pra_dat_ch0[215:208], dat_pra_dat_ch3[199:192], dat_pra_dat_ch2[199:192], dat_pra_dat_ch1[199:192], dat_pra_dat_ch0[199:192], dat_pra_dat_ch3[183:176], dat_pra_dat_ch2[183:176], dat_pra_dat_ch1[183:176], dat_pra_dat_ch0[183:176], dat_pra_dat_ch3[167:160], dat_pra_dat_ch2[167:160], dat_pra_dat_ch1[167:160], dat_pra_dat_ch0[167:160], dat_pra_dat_ch3[151:144], dat_pra_dat_ch2[151:144], dat_pra_dat_ch1[151:144], dat_pra_dat_ch0[151:144], dat_pra_dat_ch3[135:128], dat_pra_dat_ch2[135:128], dat_pra_dat_ch1[135:128], dat_pra_dat_ch0[135:128], dat_pra_dat_ch3[119:112], dat_pra_dat_ch2[119:112], dat_pra_dat_ch1[119:112], dat_pra_dat_ch0[119:112], dat_pra_dat_ch3[103:96], dat_pra_dat_ch2[103:96], dat_pra_dat_ch1[103:96], dat_pra_dat_ch0[103:96], dat_pra_dat_ch3[87:80], dat_pra_dat_ch2[87:80], dat_pra_dat_ch1[87:80], dat_pra_dat_ch0[87:80], dat_pra_dat_ch3[71:64], dat_pra_dat_ch2[71:64], dat_pra_dat_ch1[71:64], dat_pra_dat_ch0[71:64], dat_pra_dat_ch3[55:48], dat_pra_dat_ch2[55:48], dat_pra_dat_ch1[55:48], dat_pra_dat_ch0[55:48], dat_pra_dat_ch3[39:32], dat_pra_dat_ch2[39:32], dat_pra_dat_ch1[39:32], dat_pra_dat_ch0[39:32], dat_pra_dat_ch3[23:16], dat_pra_dat_ch2[23:16], dat_pra_dat_ch1[23:16], dat_pra_dat_ch0[23:16], dat_pra_dat_ch3[7:0], dat_pra_dat_ch2[7:0], dat_pra_dat_ch1[7:0], dat_pra_dat_ch0[7:0], dat_pra_dat_ch3[247:240], dat_pra_dat_ch2[247:240], dat_pra_dat_ch1[247:240], dat_pra_dat_ch0[247:240], dat_pra_dat_ch3[231:224], dat_pra_dat_ch2[231:224], dat_pra_dat_ch1[231:224], dat_pra_dat_ch0[231:224], dat_pra_dat_ch3[215:208], dat_pra_dat_ch2[215:208], dat_pra_dat_ch1[215:208], dat_pra_dat_ch0[215:208], dat_pra_dat_ch3[199:192], dat_pra_dat_ch2[199:192], dat_pra_dat_ch1[199:192], dat_pra_dat_ch0[199:192], dat_pra_dat_ch3[183:176], dat_pra_dat_ch2[183:176], dat_pra_dat_ch1[183:176], dat_pra_dat_ch0[183:176], dat_pra_dat_ch3[167:160], dat_pra_dat_ch2[167:160], dat_pra_dat_ch1[167:160], dat_pra_dat_ch0[167:160], dat_pra_dat_ch3[151:144], dat_pra_dat_ch2[151:144], dat_pra_dat_ch1[151:144], dat_pra_dat_ch0[151:144], dat_pra_dat_ch3[135:128], dat_pra_dat_ch2[135:128], dat_pra_dat_ch1[135:128], dat_pra_dat_ch0[135:128], dat_pra_dat_ch3[119:112], dat_pra_dat_ch2[119:112], dat_pra_dat_ch1[119:112], dat_pra_dat_ch0[119:112], dat_pra_dat_ch3[103:96], dat_pra_dat_ch2[103:96], dat_pra_dat_ch1[103:96], dat_pra_dat_ch0[103:96], dat_pra_dat_ch3[87:80], dat_pra_dat_ch2[87:80], dat_pra_dat_ch1[87:80], dat_pra_dat_ch0[87:80], dat_pra_dat_ch3[71:64], dat_pra_dat_ch2[71:64], dat_pra_dat_ch1[71:64], dat_pra_dat_ch0[71:64], dat_pra_dat_ch3[55:48], dat_pra_dat_ch2[55:48], dat_pra_dat_ch1[55:48], dat_pra_dat_ch0[55:48], dat_pra_dat_ch3[39:32], dat_pra_dat_ch2[39:32], dat_pra_dat_ch1[39:32], dat_pra_dat_ch0[39:32], dat_pra_dat_ch3[23:16], dat_pra_dat_ch2[23:16], dat_pra_dat_ch1[23:16], dat_pra_dat_ch0[23:16], dat_pra_dat_ch3[7:0], dat_pra_dat_ch2[7:0], dat_pra_dat_ch1[7:0], dat_pra_dat_ch0[7:0] } : { dat_pra_dat_ch3[255:240], dat_pra_dat_ch2[255:240], dat_pra_dat_ch1[255:240], dat_pra_dat_ch0[255:240], dat_pra_dat_ch3[239:224], dat_pra_dat_ch2[239:224], dat_pra_dat_ch1[239:224], dat_pra_dat_ch0[239:224], dat_pra_dat_ch3[223:208], dat_pra_dat_ch2[223:208], dat_pra_dat_ch1[223:208], dat_pra_dat_ch0[223:208], dat_pra_dat_ch3[207:192], dat_pra_dat_ch2[207:192], dat_pra_dat_ch1[207:192], dat_pra_dat_ch0[207:192], dat_pra_dat_ch3[191:176], dat_pra_dat_ch2[191:176], dat_pra_dat_ch1[191:176], dat_pra_dat_ch0[191:176], dat_pra_dat_ch3[175:160], dat_pra_dat_ch2[175:160], dat_pra_dat_ch1[175:160], dat_pra_dat_ch0[175:160], dat_pra_dat_ch3[159:144], dat_pra_dat_ch2[159:144], dat_pra_dat_ch1[159:144], dat_pra_dat_ch0[159:144], dat_pra_dat_ch3[143:128], dat_pra_dat_ch2[143:128], dat_pra_dat_ch1[143:128], dat_pra_dat_ch0[143:128], dat_pra_dat_ch3[127:112], dat_pra_dat_ch2[127:112], dat_pra_dat_ch1[127:112], dat_pra_dat_ch0[127:112], dat_pra_dat_ch3[111:96], dat_pra_dat_ch2[111:96], dat_pra_dat_ch1[111:96], dat_pra_dat_ch0[111:96], dat_pra_dat_ch3[95:80], dat_pra_dat_ch2[95:80], dat_pra_dat_ch1[95:80], dat_pra_dat_ch0[95:80], dat_pra_dat_ch3[79:64], dat_pra_dat_ch2[79:64], dat_pra_dat_ch1[79:64], dat_pra_dat_ch0[79:64], dat_pra_dat_ch3[63:48], dat_pra_dat_ch2[63:48], dat_pra_dat_ch1[63:48], dat_pra_dat_ch0[63:48], dat_pra_dat_ch3[47:32], dat_pra_dat_ch2[47:32], dat_pra_dat_ch1[47:32], dat_pra_dat_ch0[47:32], dat_pra_dat_ch3[31:16], dat_pra_dat_ch2[31:16], dat_pra_dat_ch1[31:16], dat_pra_dat_ch0[31:16], dat_pra_dat_ch3[15:0], dat_pra_dat_ch2[15:0], dat_pra_dat_ch1[15:0], dat_pra_dat_ch0[15:0] };
  assign _1230_ = is_fp16_d1[1] ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18424" *) { dat_out_wg_mask_fp16[127], dat_out_wg_mask_fp16[127], dat_out_wg_mask_fp16[125], dat_out_wg_mask_fp16[125], dat_out_wg_mask_fp16[123], dat_out_wg_mask_fp16[123], dat_out_wg_mask_fp16[121], dat_out_wg_mask_fp16[121], dat_out_wg_mask_fp16[119], dat_out_wg_mask_fp16[119], dat_out_wg_mask_fp16[117], dat_out_wg_mask_fp16[117], dat_out_wg_mask_fp16[115], dat_out_wg_mask_fp16[115], dat_out_wg_mask_fp16[113], dat_out_wg_mask_fp16[113], dat_out_wg_mask_fp16[111], dat_out_wg_mask_fp16[111], dat_out_wg_mask_fp16[109], dat_out_wg_mask_fp16[109], dat_out_wg_mask_fp16[107], dat_out_wg_mask_fp16[107], dat_out_wg_mask_fp16[105], dat_out_wg_mask_fp16[105], dat_out_wg_mask_fp16[103], dat_out_wg_mask_fp16[103], dat_out_wg_mask_fp16[101], dat_out_wg_mask_fp16[101], dat_out_wg_mask_fp16[99], dat_out_wg_mask_fp16[99], dat_out_wg_mask_fp16[97], dat_out_wg_mask_fp16[97], dat_out_wg_mask_fp16[95], dat_out_wg_mask_fp16[95], dat_out_wg_mask_fp16[93], dat_out_wg_mask_fp16[93], dat_out_wg_mask_fp16[91], dat_out_wg_mask_fp16[91], dat_out_wg_mask_fp16[89], dat_out_wg_mask_fp16[89], dat_out_wg_mask_fp16[87], dat_out_wg_mask_fp16[87], dat_out_wg_mask_fp16[85], dat_out_wg_mask_fp16[85], dat_out_wg_mask_fp16[83], dat_out_wg_mask_fp16[83], dat_out_wg_mask_fp16[81], dat_out_wg_mask_fp16[81], dat_out_wg_mask_fp16[79], dat_out_wg_mask_fp16[79], dat_out_wg_mask_fp16[77], dat_out_wg_mask_fp16[77], dat_out_wg_mask_fp16[75], dat_out_wg_mask_fp16[75], dat_out_wg_mask_fp16[73], dat_out_wg_mask_fp16[73], dat_out_wg_mask_fp16[71], dat_out_wg_mask_fp16[71], dat_out_wg_mask_fp16[69], dat_out_wg_mask_fp16[69], dat_out_wg_mask_fp16[67], dat_out_wg_mask_fp16[67], dat_out_wg_mask_fp16[65], dat_out_wg_mask_fp16[65], dat_out_wg_mask_fp16[63], dat_out_wg_mask_fp16[63], dat_out_wg_mask_fp16[61], dat_out_wg_mask_fp16[61], dat_out_wg_mask_fp16[59], dat_out_wg_mask_fp16[59], dat_out_wg_mask_fp16[57], dat_out_wg_mask_fp16[57], dat_out_wg_mask_fp16[55], dat_out_wg_mask_fp16[55], dat_out_wg_mask_fp16[53], dat_out_wg_mask_fp16[53], dat_out_wg_mask_fp16[51], dat_out_wg_mask_fp16[51], dat_out_wg_mask_fp16[49], dat_out_wg_mask_fp16[49], dat_out_wg_mask_fp16[47], dat_out_wg_mask_fp16[47], dat_out_wg_mask_fp16[45], dat_out_wg_mask_fp16[45], dat_out_wg_mask_fp16[43], dat_out_wg_mask_fp16[43], dat_out_wg_mask_fp16[41], dat_out_wg_mask_fp16[41], dat_out_wg_mask_fp16[39], dat_out_wg_mask_fp16[39], dat_out_wg_mask_fp16[37], dat_out_wg_mask_fp16[37], dat_out_wg_mask_fp16[35], dat_out_wg_mask_fp16[35], dat_out_wg_mask_fp16[33], dat_out_wg_mask_fp16[33], dat_out_wg_mask_fp16[31], dat_out_wg_mask_fp16[31], dat_out_wg_mask_fp16[29], dat_out_wg_mask_fp16[29], dat_out_wg_mask_fp16[27], dat_out_wg_mask_fp16[27], dat_out_wg_mask_fp16[25], dat_out_wg_mask_fp16[25], dat_out_wg_mask_fp16[23], dat_out_wg_mask_fp16[23], dat_out_wg_mask_fp16[21], dat_out_wg_mask_fp16[21], dat_out_wg_mask_fp16[19], dat_out_wg_mask_fp16[19], dat_out_wg_mask_fp16[17], dat_out_wg_mask_fp16[17], dat_out_wg_mask_fp16[15], dat_out_wg_mask_fp16[15], dat_out_wg_mask_fp16[13], dat_out_wg_mask_fp16[13], dat_out_wg_mask_fp16[11], dat_out_wg_mask_fp16[11], dat_out_wg_mask_fp16[9], dat_out_wg_mask_fp16[9], dat_out_wg_mask_fp16[7], dat_out_wg_mask_fp16[7], dat_out_wg_mask_fp16[5], dat_out_wg_mask_fp16[5], dat_out_wg_mask_fp16[3], dat_out_wg_mask_fp16[3], dat_out_wg_mask_fp16[1], dat_out_wg_mask_fp16[1] } : { dat_out_wg_mask_int16[127], dat_out_wg_mask_int16[127], dat_out_wg_mask_int16[125], dat_out_wg_mask_int16[125], dat_out_wg_mask_int16[123], dat_out_wg_mask_int16[123], dat_out_wg_mask_int16[121], dat_out_wg_mask_int16[121], dat_out_wg_mask_int16[119], dat_out_wg_mask_int16[119], dat_out_wg_mask_int16[117], dat_out_wg_mask_int16[117], dat_out_wg_mask_int16[115], dat_out_wg_mask_int16[115], dat_out_wg_mask_int16[113], dat_out_wg_mask_int16[113], dat_out_wg_mask_int16[111], dat_out_wg_mask_int16[111], dat_out_wg_mask_int16[109], dat_out_wg_mask_int16[109], dat_out_wg_mask_int16[107], dat_out_wg_mask_int16[107], dat_out_wg_mask_int16[105], dat_out_wg_mask_int16[105], dat_out_wg_mask_int16[103], dat_out_wg_mask_int16[103], dat_out_wg_mask_int16[101], dat_out_wg_mask_int16[101], dat_out_wg_mask_int16[99], dat_out_wg_mask_int16[99], dat_out_wg_mask_int16[97], dat_out_wg_mask_int16[97], dat_out_wg_mask_int16[95], dat_out_wg_mask_int16[95], dat_out_wg_mask_int16[93], dat_out_wg_mask_int16[93], dat_out_wg_mask_int16[91], dat_out_wg_mask_int16[91], dat_out_wg_mask_int16[89], dat_out_wg_mask_int16[89], dat_out_wg_mask_int16[87], dat_out_wg_mask_int16[87], dat_out_wg_mask_int16[85], dat_out_wg_mask_int16[85], dat_out_wg_mask_int16[83], dat_out_wg_mask_int16[83], dat_out_wg_mask_int16[81], dat_out_wg_mask_int16[81], dat_out_wg_mask_int16[79], dat_out_wg_mask_int16[79], dat_out_wg_mask_int16[77], dat_out_wg_mask_int16[77], dat_out_wg_mask_int16[75], dat_out_wg_mask_int16[75], dat_out_wg_mask_int16[73], dat_out_wg_mask_int16[73], dat_out_wg_mask_int16[71], dat_out_wg_mask_int16[71], dat_out_wg_mask_int16[69], dat_out_wg_mask_int16[69], dat_out_wg_mask_int16[67], dat_out_wg_mask_int16[67], dat_out_wg_mask_int16[65], dat_out_wg_mask_int16[65], dat_out_wg_mask_int16[63], dat_out_wg_mask_int16[63], dat_out_wg_mask_int16[61], dat_out_wg_mask_int16[61], dat_out_wg_mask_int16[59], dat_out_wg_mask_int16[59], dat_out_wg_mask_int16[57], dat_out_wg_mask_int16[57], dat_out_wg_mask_int16[55], dat_out_wg_mask_int16[55], dat_out_wg_mask_int16[53], dat_out_wg_mask_int16[53], dat_out_wg_mask_int16[51], dat_out_wg_mask_int16[51], dat_out_wg_mask_int16[49], dat_out_wg_mask_int16[49], dat_out_wg_mask_int16[47], dat_out_wg_mask_int16[47], dat_out_wg_mask_int16[45], dat_out_wg_mask_int16[45], dat_out_wg_mask_int16[43], dat_out_wg_mask_int16[43], dat_out_wg_mask_int16[41], dat_out_wg_mask_int16[41], dat_out_wg_mask_int16[39], dat_out_wg_mask_int16[39], dat_out_wg_mask_int16[37], dat_out_wg_mask_int16[37], dat_out_wg_mask_int16[35], dat_out_wg_mask_int16[35], dat_out_wg_mask_int16[33], dat_out_wg_mask_int16[33], dat_out_wg_mask_int16[31], dat_out_wg_mask_int16[31], dat_out_wg_mask_int16[29], dat_out_wg_mask_int16[29], dat_out_wg_mask_int16[27], dat_out_wg_mask_int16[27], dat_out_wg_mask_int16[25], dat_out_wg_mask_int16[25], dat_out_wg_mask_int16[23], dat_out_wg_mask_int16[23], dat_out_wg_mask_int16[21], dat_out_wg_mask_int16[21], dat_out_wg_mask_int16[19], dat_out_wg_mask_int16[19], dat_out_wg_mask_int16[17], dat_out_wg_mask_int16[17], dat_out_wg_mask_int16[15], dat_out_wg_mask_int16[15], dat_out_wg_mask_int16[13], dat_out_wg_mask_int16[13], dat_out_wg_mask_int16[11], dat_out_wg_mask_int16[11], dat_out_wg_mask_int16[9], dat_out_wg_mask_int16[9], dat_out_wg_mask_int16[7], dat_out_wg_mask_int16[7], dat_out_wg_mask_int16[5], dat_out_wg_mask_int16[5], dat_out_wg_mask_int16[3], dat_out_wg_mask_int16[3], dat_out_wg_mask_int16[1], dat_out_wg_mask_int16[1] };
  assign dat_out_wg_mask = is_int8_d1[20] ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18424" *) { dat_out_wg_mask_int8, dat_out_wg_mask_int8 } : _1230_;
  assign _1231_ = is_int8_d1[21] ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18484" *) { dat_out_bypass_data[511:0], dat_out_bypass_data[511:0] } : dat_out_bypass_data;
  assign dat_out_data = is_winograd_d1[20] ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18484" *) dat_out_wg_data : _1231_;
  assign _1232_ = is_int8_d1[22] ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18496" *) { dat_out_bypass_mask[63:0], dat_out_bypass_mask[63:0] } : dat_out_bypass_mask;
  assign _1233_ = is_winograd_d1[21] ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18496" *) dat_out_wg_mask : _1232_;
  assign dat_out_mask = dat_out_pvld ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18496" *) _1233_ : 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
  assign data_batch_w = _1150_ ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1941" *) 6'b000001 : _0713_;
  assign batch_cmp_w = _1150_ ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1948" *) 5'b00000 : reg2dp_batches;
  assign datain_width_w = reg2dp_conv_mode ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1965" *) { 2'b00, _0714_ } : _0715_;
  assign datain_channel_cmp_w = reg2dp_conv_mode ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1982" *) reg2dp_weight_channel_ext[12:2] : { 4'b0000, reg2dp_weight_channel_ext[12:6] };
  assign { sub_h_total_w, mon_sub_h_total_w } = is_img ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1990" *) _1167_ : 6'b001000;
  assign sc2mac_dat_pd_w = dl_out_pvld ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:19914" *) dl_out_flag : 9'b000000000;
  assign _1234_[1:0] = reg2dp_conv_mode ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1999" *) 2'b10 : 2'b01;
  assign sub_h_cmp_w = is_img ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:1999" *) sub_h_total_w : { 1'b0, _1234_[1:0] };
  assign conv_x_stride_w = reg2dp_conv_mode ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:2011" *) 4'b0001 : _0716_;
  assign _1235_ = _1056_ ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:2019" *) _0717_ : { 2'b00, conv_x_stride_w };
  assign pixel_x_stride_w = _1055_ ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:2019" *) { conv_x_stride_w, 2'b00 } : _1235_;
  assign _1236_ = _1065_ ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:2030" *) 6'b111111 : reg2dp_weight_channel_ext[5:0];
  assign _1237_[5:0] = _1058_ ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:2030" *) _0720_ : _1236_;
  assign pixel_x_init_w = _1057_ ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:2030" *) _0719_ : _1237_[5:0];
  assign _1238_[6:0] = _1058_ ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:2043" *) { pixel_x_stride_w, 1'b0 } : { 1'b0, pixel_x_stride_w };
  assign pixel_x_add_w = _1057_ ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:2043" *) { pixel_x_stride_w[4:0], 2'b00 } : _1238_[6:0];
  assign pixel_x_byte_stride_w = is_int8 ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:2049" *) { 1'b0, pixel_x_stride_w } : { pixel_x_stride_w, 1'b0 };
  assign conv_y_stride_w = reg2dp_conv_mode ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:2061" *) 4'b0001 : _0721_;
  assign x_dilate_w = _1150_ ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:2069" *) 6'b000001 : _0722_;
  assign y_dilate_w = _1150_ ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:2077" *) 6'b000001 : _0723_;
  assign entries_w = reg2dp_conv_mode ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:2099" *) _0724_ : entries_single_w;
  assign slice_left_w = reg2dp_skip_data_rls ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:2134" *) _0725_ : _1020_[11:0];
  assign slices_oprand = layer_st_d1 ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:2142" *) rls_slices : slice_left;
  assign pra_truncate_w = _1059_ ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:2160" *) 2'b10 : reg2dp_pra_truncate;
  assign dat_entry_avl_sub = dat_rls ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:6685" *) sc2cdma_dat_entries_w : 12'b000000000000;
  assign _1239_ = is_dat_entry_st_wrap ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:6725" *) dat_entry_st_inc_wrap : dat_entry_st_inc[11:0];
  assign dat_entry_st_w = sc2cdma_dat_pending_req ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:6725" *) 12'b000000000000 : _1239_;
  assign sc2cdma_dat_slices_w = sub_rls ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:7454" *) rls_slices : last_slices;
  assign sc2cdma_dat_entries_w = sub_rls ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:7462" *) rls_entries : last_entries;
  assign dl_in_pvld = is_winograd_d1[0] ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:8223" *) sg2dl_pvld : dl_in_pvld_d5;
  assign dl_pd_d0 = is_winograd_d1[1] ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:8224" *) sg2dl_pd : dl_in_pd_d5;
  assign _1240_[4:0] = is_batch_end ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:8539" *) 5'b00000 : _0726_[4:0];
  assign batch_cnt_w = layer_st ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:8539" *) 5'b00000 : _1240_[4:0];
  assign sub_h_cnt_w = _1153_ ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:8714" *) 2'b00 : sub_h_cnt_inc[1:0];
  assign _1241_ = is_stripe_end ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:8809" *) 7'b0000000 : stripe_cnt_inc;
  assign _1242_ = _0984_ ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:8809" *) stripe_cnt : _1241_;
  assign stripe_cnt_w = layer_st ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:8809" *) 7'b0000000 : _1242_;
  assign _1243_ = dat_req_stripe_st ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:9089" *) 1'b1 : dat_pipe_local_valid;
  assign dat_pipe_local_valid_w = dat_req_stripe_end ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:9089" *) 1'b0 : _1243_;
  assign _1244_ = _0987_ ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:9101" *) 1'b0 : dat_exec_valid_d1;
  assign dat_exec_valid = dat_req_stripe_st ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:9101" *) 1'b1 : _1244_;
  assign dat_req_bytes = is_int8_d1[0] ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:9176" *) { 1'b0, dl_pd[16:10] } : { dl_pd[16:10], 1'b0 };
  assign _1245_ = is_w_end ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:9369" *) { dataout_w_init[12], dataout_w_init[12], dataout_w_init[12], dataout_w_init[12], dataout_w_init[12], dataout_w_init[12], dataout_w_init[12], dataout_w_init[12], dataout_w_init[12], dataout_w_init[12], dataout_w_init[2:0] } : dataout_w_cnt_inc;
  assign _1246_ = _0733_ ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:9369" *) dataout_w_ori : _1245_;
  assign dataout_w_cnt_w = layer_st ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:9369" *) { dataout_w_init[12], dataout_w_init[12], dataout_w_init[12], dataout_w_init[12], dataout_w_init[12], dataout_w_init[12], dataout_w_init[12], dataout_w_init[12], dataout_w_init[12], dataout_w_init[12], dataout_w_init[2:0] } : _1246_;
  assign _1247_ = dl_pd[27] ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:9529" *) 11'b00000000000 : datain_c_cnt_inc;
  assign datain_c_cnt_w = layer_st ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:9529" *) 11'b00000000000 : _1247_;
  assign _1248_ = reg2dp_conv_mode ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:9608" *) 14'b00000000000010 : { _1169_[13], _1169_[13], _1169_[13], _1169_[13], _1169_[13], _1169_[13], _1169_[13], _1169_[13], _1169_[13], _1169_[4:0] };
  assign datain_w_cnt_st = is_img ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:9608" *) 14'b00000000000000 : _1248_;
  assign datain_w_cnt_inc = is_winograd_d1[3] ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:9617" *) _0727_[13:0] : _0728_[13:0];
  assign _1249_ = is_w_end ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:9631" *) datain_w_cnt_st : datain_w_cnt_inc;
  assign _1250_ = _0733_ ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:9631" *) datain_w_ori : _1249_;
  assign datain_w_cnt_w = layer_st ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:9631" *) datain_w_cnt_st : _1250_;
  assign pixel_x_cnt_add = is_sub_h_end ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:9637" *) pixel_x_add : 7'b0000000;
  assign _1251_[15:0] = _0995_ ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:9659" *) pixel_w_ori : _0731_[15:0];
  assign _1252_[15:0] = _0994_ ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:9659" *) _0730_[15:0] : _1251_[15:0];
  assign _1253_[15:0] = _0993_ ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:9659" *) _0729_[15:0] : _1252_[15:0];
  assign _1254_[15:0] = _0992_ ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:9659" *) { 10'b0000000000, pixel_x_init } : _1253_[15:0];
  assign pixel_w_cnt_w = layer_st_d1 ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:9659" *) { 10'b0000000000, pixel_x_init } : _1254_[15:0];
  assign _1255_ = _1014_ ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:9736" *) _1122_ : pixel_req_ch_odd;
  assign _1256_ = _1013_ ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:9736" *) pixel_req_ch_odd_ori : _1255_;
  assign _1257_ = _1012_ ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:9736" *) _1120_ : _1256_;
  assign _1258_ = _1009_ ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:9736" *) 1'b0 : _1257_;
  assign pixel_req_ch_odd_w = layer_st_d1 ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:9736" *) 1'b0 : _1258_;
  assign _1259_ = pixel_force_clr_d1 ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:9742" *) 1'b0 : pixel_force_fetch_d1;
  assign pixel_force_fetch = _1015_ ? (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:9742" *) 1'b1 : _1259_;
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18260" *)
  NV_NVDLA_CSC_pra_cell u_pra_cell_0 (
    .cfg_precision(pra_precision[1:0]),
    .cfg_truncate_rsc_z(pra_truncate[1:0]),
    .chn_data_in_rsc_lz(mon_dat_rsp_pra_rdy[0]),
    .chn_data_in_rsc_vz(dat_rsp_pra_en_d1[0]),
    .chn_data_in_rsc_z(dat_rsp_wg_ch0_d1),
    .chn_data_out_rsc_lz(mon_dat_out_pra_vld[0]),
    .chn_data_out_rsc_vz(1'b1),
    .chn_data_out_rsc_z(dat_pra_dat_ch0),
    .nvdla_core_clk(nvdla_wg_clk),
    .nvdla_core_rstn(nvdla_core_rstn)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18276" *)
  NV_NVDLA_CSC_pra_cell u_pra_cell_1 (
    .cfg_precision(pra_precision[3:2]),
    .cfg_truncate_rsc_z(pra_truncate[3:2]),
    .chn_data_in_rsc_lz(mon_dat_rsp_pra_rdy[1]),
    .chn_data_in_rsc_vz(dat_rsp_pra_en_d1[0]),
    .chn_data_in_rsc_z(dat_rsp_wg_ch1_d1),
    .chn_data_out_rsc_lz(mon_dat_out_pra_vld[1]),
    .chn_data_out_rsc_vz(1'b1),
    .chn_data_out_rsc_z(dat_pra_dat_ch1),
    .nvdla_core_clk(nvdla_wg_clk),
    .nvdla_core_rstn(nvdla_core_rstn)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18292" *)
  NV_NVDLA_CSC_pra_cell u_pra_cell_2 (
    .cfg_precision(pra_precision[5:4]),
    .cfg_truncate_rsc_z(pra_truncate[5:4]),
    .chn_data_in_rsc_lz(mon_dat_rsp_pra_rdy[2]),
    .chn_data_in_rsc_vz(dat_rsp_pra_en_d1[0]),
    .chn_data_in_rsc_z(dat_rsp_wg_ch2_d1),
    .chn_data_out_rsc_lz(mon_dat_out_pra_vld[2]),
    .chn_data_out_rsc_vz(1'b1),
    .chn_data_out_rsc_z(dat_pra_dat_ch2),
    .nvdla_core_clk(nvdla_wg_clk),
    .nvdla_core_rstn(nvdla_core_rstn)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_dl.v:18308" *)
  NV_NVDLA_CSC_pra_cell u_pra_cell_3 (
    .cfg_precision(pra_precision[7:6]),
    .cfg_truncate_rsc_z(pra_truncate[7:6]),
    .chn_data_in_rsc_lz(mon_dat_rsp_pra_rdy[3]),
    .chn_data_in_rsc_vz(dat_rsp_pra_en_d1[0]),
    .chn_data_in_rsc_z(dat_rsp_wg_ch3_d1),
    .chn_data_out_rsc_lz(mon_dat_out_pra_vld[3]),
    .chn_data_out_rsc_vz(1'b1),
    .chn_data_out_rsc_z(dat_pra_dat_ch3),
    .nvdla_core_clk(nvdla_wg_clk),
    .nvdla_core_rstn(nvdla_core_rstn)
  );
  assign _1017_[11:0] = _0769_;
  assign _1018_[12:0] = _0980_;
  assign _1020_[14:13] = { _1020_[15], _1020_[15] };
  assign _1021_[14] = 1'b0;
  assign _1022_[14] = 1'bx;
  assign _1023_[14] = 1'bx;
  assign _1024_[14] = 1'bx;
  assign _1025_[14] = 1'bx;
  assign _1168_[12:5] = { _1168_[13], _1168_[13], _1168_[13], _1168_[13], _1168_[13], _1168_[13], _1168_[13], _1168_[13] };
  assign _1169_[12:5] = { _1169_[13], _1169_[13], _1169_[13], _1169_[13], _1169_[13], _1169_[13], _1169_[13], _1169_[13] };
  assign _1173_[12] = 1'bx;
  assign _1234_[2] = 1'b0;
  assign _1237_[7:6] = 2'b0x;
  assign _1238_[7] = 1'b0;
  assign _1240_[5] = 1'bx;
  assign _1251_[16] = 1'bx;
  assign _1252_[16] = 1'bx;
  assign _1253_[16] = 1'bx;
  assign _1254_[16] = 1'bx;
  assign cbuf_reset = sc2cdma_dat_pending_req;
  assign dat_out_flag_l0 = dat_rsp_pd[26:18];
  assign dat_out_pvld_l0 = dat_rsp_pvld;
  assign dat_out_wg_16b = { dat_pra_dat_ch3[255:240], dat_pra_dat_ch2[255:240], dat_pra_dat_ch1[255:240], dat_pra_dat_ch0[255:240], dat_pra_dat_ch3[239:224], dat_pra_dat_ch2[239:224], dat_pra_dat_ch1[239:224], dat_pra_dat_ch0[239:224], dat_pra_dat_ch3[223:208], dat_pra_dat_ch2[223:208], dat_pra_dat_ch1[223:208], dat_pra_dat_ch0[223:208], dat_pra_dat_ch3[207:192], dat_pra_dat_ch2[207:192], dat_pra_dat_ch1[207:192], dat_pra_dat_ch0[207:192], dat_pra_dat_ch3[191:176], dat_pra_dat_ch2[191:176], dat_pra_dat_ch1[191:176], dat_pra_dat_ch0[191:176], dat_pra_dat_ch3[175:160], dat_pra_dat_ch2[175:160], dat_pra_dat_ch1[175:160], dat_pra_dat_ch0[175:160], dat_pra_dat_ch3[159:144], dat_pra_dat_ch2[159:144], dat_pra_dat_ch1[159:144], dat_pra_dat_ch0[159:144], dat_pra_dat_ch3[143:128], dat_pra_dat_ch2[143:128], dat_pra_dat_ch1[143:128], dat_pra_dat_ch0[143:128], dat_pra_dat_ch3[127:112], dat_pra_dat_ch2[127:112], dat_pra_dat_ch1[127:112], dat_pra_dat_ch0[127:112], dat_pra_dat_ch3[111:96], dat_pra_dat_ch2[111:96], dat_pra_dat_ch1[111:96], dat_pra_dat_ch0[111:96], dat_pra_dat_ch3[95:80], dat_pra_dat_ch2[95:80], dat_pra_dat_ch1[95:80], dat_pra_dat_ch0[95:80], dat_pra_dat_ch3[79:64], dat_pra_dat_ch2[79:64], dat_pra_dat_ch1[79:64], dat_pra_dat_ch0[79:64], dat_pra_dat_ch3[63:48], dat_pra_dat_ch2[63:48], dat_pra_dat_ch1[63:48], dat_pra_dat_ch0[63:48], dat_pra_dat_ch3[47:32], dat_pra_dat_ch2[47:32], dat_pra_dat_ch1[47:32], dat_pra_dat_ch0[47:32], dat_pra_dat_ch3[31:16], dat_pra_dat_ch2[31:16], dat_pra_dat_ch1[31:16], dat_pra_dat_ch0[31:16], dat_pra_dat_ch3[15:0], dat_pra_dat_ch2[15:0], dat_pra_dat_ch1[15:0], dat_pra_dat_ch0[15:0] };
  assign dat_out_wg_8b = { dat_pra_dat_ch3[247:240], dat_pra_dat_ch2[247:240], dat_pra_dat_ch1[247:240], dat_pra_dat_ch0[247:240], dat_pra_dat_ch3[231:224], dat_pra_dat_ch2[231:224], dat_pra_dat_ch1[231:224], dat_pra_dat_ch0[231:224], dat_pra_dat_ch3[215:208], dat_pra_dat_ch2[215:208], dat_pra_dat_ch1[215:208], dat_pra_dat_ch0[215:208], dat_pra_dat_ch3[199:192], dat_pra_dat_ch2[199:192], dat_pra_dat_ch1[199:192], dat_pra_dat_ch0[199:192], dat_pra_dat_ch3[183:176], dat_pra_dat_ch2[183:176], dat_pra_dat_ch1[183:176], dat_pra_dat_ch0[183:176], dat_pra_dat_ch3[167:160], dat_pra_dat_ch2[167:160], dat_pra_dat_ch1[167:160], dat_pra_dat_ch0[167:160], dat_pra_dat_ch3[151:144], dat_pra_dat_ch2[151:144], dat_pra_dat_ch1[151:144], dat_pra_dat_ch0[151:144], dat_pra_dat_ch3[135:128], dat_pra_dat_ch2[135:128], dat_pra_dat_ch1[135:128], dat_pra_dat_ch0[135:128], dat_pra_dat_ch3[119:112], dat_pra_dat_ch2[119:112], dat_pra_dat_ch1[119:112], dat_pra_dat_ch0[119:112], dat_pra_dat_ch3[103:96], dat_pra_dat_ch2[103:96], dat_pra_dat_ch1[103:96], dat_pra_dat_ch0[103:96], dat_pra_dat_ch3[87:80], dat_pra_dat_ch2[87:80], dat_pra_dat_ch1[87:80], dat_pra_dat_ch0[87:80], dat_pra_dat_ch3[71:64], dat_pra_dat_ch2[71:64], dat_pra_dat_ch1[71:64], dat_pra_dat_ch0[71:64], dat_pra_dat_ch3[55:48], dat_pra_dat_ch2[55:48], dat_pra_dat_ch1[55:48], dat_pra_dat_ch0[55:48], dat_pra_dat_ch3[39:32], dat_pra_dat_ch2[39:32], dat_pra_dat_ch1[39:32], dat_pra_dat_ch0[39:32], dat_pra_dat_ch3[23:16], dat_pra_dat_ch2[23:16], dat_pra_dat_ch1[23:16], dat_pra_dat_ch0[23:16], dat_pra_dat_ch3[7:0], dat_pra_dat_ch2[7:0], dat_pra_dat_ch1[7:0], dat_pra_dat_ch0[7:0] };
  assign { dat_out_wg_mask_fp16[126], dat_out_wg_mask_fp16[124], dat_out_wg_mask_fp16[122], dat_out_wg_mask_fp16[120], dat_out_wg_mask_fp16[118], dat_out_wg_mask_fp16[116], dat_out_wg_mask_fp16[114], dat_out_wg_mask_fp16[112], dat_out_wg_mask_fp16[110], dat_out_wg_mask_fp16[108], dat_out_wg_mask_fp16[106], dat_out_wg_mask_fp16[104], dat_out_wg_mask_fp16[102], dat_out_wg_mask_fp16[100], dat_out_wg_mask_fp16[98], dat_out_wg_mask_fp16[96], dat_out_wg_mask_fp16[94], dat_out_wg_mask_fp16[92], dat_out_wg_mask_fp16[90], dat_out_wg_mask_fp16[88], dat_out_wg_mask_fp16[86], dat_out_wg_mask_fp16[84], dat_out_wg_mask_fp16[82], dat_out_wg_mask_fp16[80], dat_out_wg_mask_fp16[78], dat_out_wg_mask_fp16[76], dat_out_wg_mask_fp16[74], dat_out_wg_mask_fp16[72], dat_out_wg_mask_fp16[70], dat_out_wg_mask_fp16[68], dat_out_wg_mask_fp16[66], dat_out_wg_mask_fp16[64], dat_out_wg_mask_fp16[62], dat_out_wg_mask_fp16[60], dat_out_wg_mask_fp16[58], dat_out_wg_mask_fp16[56], dat_out_wg_mask_fp16[54], dat_out_wg_mask_fp16[52], dat_out_wg_mask_fp16[50], dat_out_wg_mask_fp16[48], dat_out_wg_mask_fp16[46], dat_out_wg_mask_fp16[44], dat_out_wg_mask_fp16[42], dat_out_wg_mask_fp16[40], dat_out_wg_mask_fp16[38], dat_out_wg_mask_fp16[36], dat_out_wg_mask_fp16[34], dat_out_wg_mask_fp16[32], dat_out_wg_mask_fp16[30], dat_out_wg_mask_fp16[28], dat_out_wg_mask_fp16[26], dat_out_wg_mask_fp16[24], dat_out_wg_mask_fp16[22], dat_out_wg_mask_fp16[20], dat_out_wg_mask_fp16[18], dat_out_wg_mask_fp16[16], dat_out_wg_mask_fp16[14], dat_out_wg_mask_fp16[12], dat_out_wg_mask_fp16[10], dat_out_wg_mask_fp16[8], dat_out_wg_mask_fp16[6], dat_out_wg_mask_fp16[4], dat_out_wg_mask_fp16[2], dat_out_wg_mask_fp16[0] } = { dat_out_wg_mask_fp16[127], dat_out_wg_mask_fp16[125], dat_out_wg_mask_fp16[123], dat_out_wg_mask_fp16[121], dat_out_wg_mask_fp16[119], dat_out_wg_mask_fp16[117], dat_out_wg_mask_fp16[115], dat_out_wg_mask_fp16[113], dat_out_wg_mask_fp16[111], dat_out_wg_mask_fp16[109], dat_out_wg_mask_fp16[107], dat_out_wg_mask_fp16[105], dat_out_wg_mask_fp16[103], dat_out_wg_mask_fp16[101], dat_out_wg_mask_fp16[99], dat_out_wg_mask_fp16[97], dat_out_wg_mask_fp16[95], dat_out_wg_mask_fp16[93], dat_out_wg_mask_fp16[91], dat_out_wg_mask_fp16[89], dat_out_wg_mask_fp16[87], dat_out_wg_mask_fp16[85], dat_out_wg_mask_fp16[83], dat_out_wg_mask_fp16[81], dat_out_wg_mask_fp16[79], dat_out_wg_mask_fp16[77], dat_out_wg_mask_fp16[75], dat_out_wg_mask_fp16[73], dat_out_wg_mask_fp16[71], dat_out_wg_mask_fp16[69], dat_out_wg_mask_fp16[67], dat_out_wg_mask_fp16[65], dat_out_wg_mask_fp16[63], dat_out_wg_mask_fp16[61], dat_out_wg_mask_fp16[59], dat_out_wg_mask_fp16[57], dat_out_wg_mask_fp16[55], dat_out_wg_mask_fp16[53], dat_out_wg_mask_fp16[51], dat_out_wg_mask_fp16[49], dat_out_wg_mask_fp16[47], dat_out_wg_mask_fp16[45], dat_out_wg_mask_fp16[43], dat_out_wg_mask_fp16[41], dat_out_wg_mask_fp16[39], dat_out_wg_mask_fp16[37], dat_out_wg_mask_fp16[35], dat_out_wg_mask_fp16[33], dat_out_wg_mask_fp16[31], dat_out_wg_mask_fp16[29], dat_out_wg_mask_fp16[27], dat_out_wg_mask_fp16[25], dat_out_wg_mask_fp16[23], dat_out_wg_mask_fp16[21], dat_out_wg_mask_fp16[19], dat_out_wg_mask_fp16[17], dat_out_wg_mask_fp16[15], dat_out_wg_mask_fp16[13], dat_out_wg_mask_fp16[11], dat_out_wg_mask_fp16[9], dat_out_wg_mask_fp16[7], dat_out_wg_mask_fp16[5], dat_out_wg_mask_fp16[3], dat_out_wg_mask_fp16[1] };
  assign { dat_out_wg_mask_int16[126], dat_out_wg_mask_int16[124], dat_out_wg_mask_int16[122], dat_out_wg_mask_int16[120], dat_out_wg_mask_int16[118], dat_out_wg_mask_int16[116], dat_out_wg_mask_int16[114], dat_out_wg_mask_int16[112], dat_out_wg_mask_int16[110], dat_out_wg_mask_int16[108], dat_out_wg_mask_int16[106], dat_out_wg_mask_int16[104], dat_out_wg_mask_int16[102], dat_out_wg_mask_int16[100], dat_out_wg_mask_int16[98], dat_out_wg_mask_int16[96], dat_out_wg_mask_int16[94], dat_out_wg_mask_int16[92], dat_out_wg_mask_int16[90], dat_out_wg_mask_int16[88], dat_out_wg_mask_int16[86], dat_out_wg_mask_int16[84], dat_out_wg_mask_int16[82], dat_out_wg_mask_int16[80], dat_out_wg_mask_int16[78], dat_out_wg_mask_int16[76], dat_out_wg_mask_int16[74], dat_out_wg_mask_int16[72], dat_out_wg_mask_int16[70], dat_out_wg_mask_int16[68], dat_out_wg_mask_int16[66], dat_out_wg_mask_int16[64], dat_out_wg_mask_int16[62], dat_out_wg_mask_int16[60], dat_out_wg_mask_int16[58], dat_out_wg_mask_int16[56], dat_out_wg_mask_int16[54], dat_out_wg_mask_int16[52], dat_out_wg_mask_int16[50], dat_out_wg_mask_int16[48], dat_out_wg_mask_int16[46], dat_out_wg_mask_int16[44], dat_out_wg_mask_int16[42], dat_out_wg_mask_int16[40], dat_out_wg_mask_int16[38], dat_out_wg_mask_int16[36], dat_out_wg_mask_int16[34], dat_out_wg_mask_int16[32], dat_out_wg_mask_int16[30], dat_out_wg_mask_int16[28], dat_out_wg_mask_int16[26], dat_out_wg_mask_int16[24], dat_out_wg_mask_int16[22], dat_out_wg_mask_int16[20], dat_out_wg_mask_int16[18], dat_out_wg_mask_int16[16], dat_out_wg_mask_int16[14], dat_out_wg_mask_int16[12], dat_out_wg_mask_int16[10], dat_out_wg_mask_int16[8], dat_out_wg_mask_int16[6], dat_out_wg_mask_int16[4], dat_out_wg_mask_int16[2], dat_out_wg_mask_int16[0] } = { dat_out_wg_mask_int16[127], dat_out_wg_mask_int16[125], dat_out_wg_mask_int16[123], dat_out_wg_mask_int16[121], dat_out_wg_mask_int16[119], dat_out_wg_mask_int16[117], dat_out_wg_mask_int16[115], dat_out_wg_mask_int16[113], dat_out_wg_mask_int16[111], dat_out_wg_mask_int16[109], dat_out_wg_mask_int16[107], dat_out_wg_mask_int16[105], dat_out_wg_mask_int16[103], dat_out_wg_mask_int16[101], dat_out_wg_mask_int16[99], dat_out_wg_mask_int16[97], dat_out_wg_mask_int16[95], dat_out_wg_mask_int16[93], dat_out_wg_mask_int16[91], dat_out_wg_mask_int16[89], dat_out_wg_mask_int16[87], dat_out_wg_mask_int16[85], dat_out_wg_mask_int16[83], dat_out_wg_mask_int16[81], dat_out_wg_mask_int16[79], dat_out_wg_mask_int16[77], dat_out_wg_mask_int16[75], dat_out_wg_mask_int16[73], dat_out_wg_mask_int16[71], dat_out_wg_mask_int16[69], dat_out_wg_mask_int16[67], dat_out_wg_mask_int16[65], dat_out_wg_mask_int16[63], dat_out_wg_mask_int16[61], dat_out_wg_mask_int16[59], dat_out_wg_mask_int16[57], dat_out_wg_mask_int16[55], dat_out_wg_mask_int16[53], dat_out_wg_mask_int16[51], dat_out_wg_mask_int16[49], dat_out_wg_mask_int16[47], dat_out_wg_mask_int16[45], dat_out_wg_mask_int16[43], dat_out_wg_mask_int16[41], dat_out_wg_mask_int16[39], dat_out_wg_mask_int16[37], dat_out_wg_mask_int16[35], dat_out_wg_mask_int16[33], dat_out_wg_mask_int16[31], dat_out_wg_mask_int16[29], dat_out_wg_mask_int16[27], dat_out_wg_mask_int16[25], dat_out_wg_mask_int16[23], dat_out_wg_mask_int16[21], dat_out_wg_mask_int16[19], dat_out_wg_mask_int16[17], dat_out_wg_mask_int16[15], dat_out_wg_mask_int16[13], dat_out_wg_mask_int16[11], dat_out_wg_mask_int16[9], dat_out_wg_mask_int16[7], dat_out_wg_mask_int16[5], dat_out_wg_mask_int16[3], dat_out_wg_mask_int16[1] };
  assign dat_pra_dat = { dat_pra_dat_ch3, dat_pra_dat_ch2, dat_pra_dat_ch1, dat_pra_dat_ch0 };
  assign dat_req_base_d1 = dat_entry_st;
  assign dat_req_batch_index = batch_cnt;
  assign dat_req_channel_end = dl_pd[27];
  assign dat_req_exec_dummy = dat_req_dummy_d2;
  assign dat_req_exec_pvld = dat_exec_valid_d2;
  assign dat_req_exec_sub_h = dat_req_sub_h_d2;
  assign dat_req_flag_w = { dl_pd[29], dl_pd[27], dat_req_stripe_end, dat_req_stripe_st, batch_cnt };
  assign dat_req_layer_end = dl_pd[29];
  assign dat_req_pipe_bytes = dat_req_bytes_d2;
  assign dat_req_pipe_ch_end = dat_req_ch_end_d2;
  assign dat_req_pipe_ch_odd = dat_req_ch_odd_d2;
  assign dat_req_pipe_cur_sub_h = dat_req_cur_sub_h_d2;
  assign dat_req_pipe_dummy = dat_req_dummy_d2;
  assign dat_req_pipe_flag = dat_req_flag_d2;
  assign dat_req_pipe_pd = { dat_req_flag_d2, dat_req_rls_d2, dat_req_sub_w_st_d2, dat_req_dummy_d2, dat_req_cur_sub_h_d2, dat_req_bytes_d2, dat_req_ch_odd_d2, dat_req_ch_end_d2, dat_req_sub_c_d2, dat_req_sub_h_d2, dat_req_sub_w_d2 };
  assign dat_req_pipe_pvld = dat_pipe_valid_d2;
  assign dat_req_pipe_rls = dat_req_rls_d2;
  assign dat_req_pipe_sub_c = dat_req_sub_c_d2;
  assign dat_req_pipe_sub_h = dat_req_sub_h_d2;
  assign dat_req_pipe_sub_w = dat_req_sub_w_d2;
  assign dat_req_pipe_sub_w_st = dat_req_sub_w_st_d2;
  assign dat_rsp_batch_index = dat_rsp_pd[22:18];
  assign dat_rsp_bytes = dat_rsp_pd[14:7];
  assign dat_rsp_ch_end = dat_rsp_pd[5];
  assign dat_rsp_ch_odd = dat_rsp_pd[6];
  assign dat_rsp_channel_end = dat_rsp_pd[25];
  assign dat_rsp_cur_h_e2_mask_16b = { dat_rsp_cur_h_mask_p1, 64'b1111111111111111111111111111111111111111111111111111111111111111 };
  assign dat_rsp_cur_h_e2_mask_8b = { dat_rsp_cur_h_mask_p1[31:0], 32'b11111111111111111111111111111111 };
  assign dat_rsp_cur_h_e4_mask_16b = { dat_rsp_cur_h_mask_p3, dat_rsp_cur_h_mask_p2, dat_rsp_cur_h_mask_p1[31:0], 32'b11111111111111111111111111111111 };
  assign dat_rsp_cur_h_e4_mask_8b = { dat_rsp_cur_h_mask_p3[15:0], dat_rsp_cur_h_mask_p2[15:0], dat_rsp_cur_h_mask_p1[15:0], 16'b1111111111111111 };
  assign dat_rsp_cur_sub_h = dat_rsp_pd[16:15];
  assign dat_rsp_data_w = dat_out_bypass_data_w;
  assign dat_rsp_exec_dummy = dat_rsp_exec_dummy_d6;
  assign dat_rsp_exec_dummy_d0 = dat_req_dummy_d2;
  assign dat_rsp_exec_pvld = dat_rsp_exec_pvld_d6;
  assign dat_rsp_exec_pvld_d0 = dat_exec_valid_d2;
  assign dat_rsp_exec_sub_h = dat_rsp_exec_sub_h_d6;
  assign dat_rsp_exec_sub_h_d0 = dat_req_sub_h_d2;
  assign dat_rsp_flag = dat_rsp_pd[26:18];
  assign dat_rsp_l0_block_end = dat_rsp_pd_d1[4];
  assign dat_rsp_l0_ch_odd = dat_rsp_pd_d1[6];
  assign dat_rsp_l0_flag = dat_rsp_pd_d1[26:18];
  assign dat_rsp_l0_pvld = dat_rsp_pvld_d1;
  assign dat_rsp_l0_stripe_end = dat_rsp_pd_d1[24];
  assign dat_rsp_l0_sub_c = dat_rsp_pd_d1[4];
  assign dat_rsp_l1_block_end = dat_rsp_pd_d2[4];
  assign dat_rsp_l1_ch_odd = dat_rsp_pd_d2[6];
  assign dat_rsp_l1_flag = dat_rsp_pd_d2[26:18];
  assign dat_rsp_l1_pvld = dat_rsp_pvld_d2;
  assign dat_rsp_l1_stripe_end = dat_rsp_pd_d2[24];
  assign dat_rsp_l1_sub_c = dat_rsp_pd_d2[4];
  assign dat_rsp_l2_block_end = dat_rsp_pd_d3[4];
  assign dat_rsp_l2_ch_odd = dat_rsp_pd_d3[6];
  assign dat_rsp_l2_flag = dat_rsp_pd_d3[26:18];
  assign dat_rsp_l2_pvld = dat_rsp_pvld_d3;
  assign dat_rsp_l2_stripe_end = dat_rsp_pd_d3[24];
  assign dat_rsp_l2_sub_c = dat_rsp_pd_d3[4];
  assign dat_rsp_l3_block_end = dat_rsp_pd_d4[4];
  assign dat_rsp_l3_ch_odd = dat_rsp_pd_d4[6];
  assign dat_rsp_l3_flag = dat_rsp_pd_d4[26:18];
  assign dat_rsp_l3_pvld = dat_rsp_pvld_d4;
  assign dat_rsp_l3_stripe_end = dat_rsp_pd_d4[24];
  assign dat_rsp_l3_sub_c = dat_rsp_pd_d4[4];
  assign dat_rsp_layer_end = dat_rsp_pd[26];
  assign { dat_rsp_mask_val_fp16[126], dat_rsp_mask_val_fp16[124], dat_rsp_mask_val_fp16[122], dat_rsp_mask_val_fp16[120], dat_rsp_mask_val_fp16[118], dat_rsp_mask_val_fp16[116], dat_rsp_mask_val_fp16[114], dat_rsp_mask_val_fp16[112], dat_rsp_mask_val_fp16[110], dat_rsp_mask_val_fp16[108], dat_rsp_mask_val_fp16[106], dat_rsp_mask_val_fp16[104], dat_rsp_mask_val_fp16[102], dat_rsp_mask_val_fp16[100], dat_rsp_mask_val_fp16[98], dat_rsp_mask_val_fp16[96], dat_rsp_mask_val_fp16[94], dat_rsp_mask_val_fp16[92], dat_rsp_mask_val_fp16[90], dat_rsp_mask_val_fp16[88], dat_rsp_mask_val_fp16[86], dat_rsp_mask_val_fp16[84], dat_rsp_mask_val_fp16[82], dat_rsp_mask_val_fp16[80], dat_rsp_mask_val_fp16[78], dat_rsp_mask_val_fp16[76], dat_rsp_mask_val_fp16[74], dat_rsp_mask_val_fp16[72], dat_rsp_mask_val_fp16[70], dat_rsp_mask_val_fp16[68], dat_rsp_mask_val_fp16[66], dat_rsp_mask_val_fp16[64], dat_rsp_mask_val_fp16[62], dat_rsp_mask_val_fp16[60], dat_rsp_mask_val_fp16[58], dat_rsp_mask_val_fp16[56], dat_rsp_mask_val_fp16[54], dat_rsp_mask_val_fp16[52], dat_rsp_mask_val_fp16[50], dat_rsp_mask_val_fp16[48], dat_rsp_mask_val_fp16[46], dat_rsp_mask_val_fp16[44], dat_rsp_mask_val_fp16[42], dat_rsp_mask_val_fp16[40], dat_rsp_mask_val_fp16[38], dat_rsp_mask_val_fp16[36], dat_rsp_mask_val_fp16[34], dat_rsp_mask_val_fp16[32], dat_rsp_mask_val_fp16[30], dat_rsp_mask_val_fp16[28], dat_rsp_mask_val_fp16[26], dat_rsp_mask_val_fp16[24], dat_rsp_mask_val_fp16[22], dat_rsp_mask_val_fp16[20], dat_rsp_mask_val_fp16[18], dat_rsp_mask_val_fp16[16], dat_rsp_mask_val_fp16[14], dat_rsp_mask_val_fp16[12], dat_rsp_mask_val_fp16[10], dat_rsp_mask_val_fp16[8], dat_rsp_mask_val_fp16[6], dat_rsp_mask_val_fp16[4], dat_rsp_mask_val_fp16[2], dat_rsp_mask_val_fp16[0] } = { dat_rsp_mask_val_fp16[127], dat_rsp_mask_val_fp16[125], dat_rsp_mask_val_fp16[123], dat_rsp_mask_val_fp16[121], dat_rsp_mask_val_fp16[119], dat_rsp_mask_val_fp16[117], dat_rsp_mask_val_fp16[115], dat_rsp_mask_val_fp16[113], dat_rsp_mask_val_fp16[111], dat_rsp_mask_val_fp16[109], dat_rsp_mask_val_fp16[107], dat_rsp_mask_val_fp16[105], dat_rsp_mask_val_fp16[103], dat_rsp_mask_val_fp16[101], dat_rsp_mask_val_fp16[99], dat_rsp_mask_val_fp16[97], dat_rsp_mask_val_fp16[95], dat_rsp_mask_val_fp16[93], dat_rsp_mask_val_fp16[91], dat_rsp_mask_val_fp16[89], dat_rsp_mask_val_fp16[87], dat_rsp_mask_val_fp16[85], dat_rsp_mask_val_fp16[83], dat_rsp_mask_val_fp16[81], dat_rsp_mask_val_fp16[79], dat_rsp_mask_val_fp16[77], dat_rsp_mask_val_fp16[75], dat_rsp_mask_val_fp16[73], dat_rsp_mask_val_fp16[71], dat_rsp_mask_val_fp16[69], dat_rsp_mask_val_fp16[67], dat_rsp_mask_val_fp16[65], dat_rsp_mask_val_fp16[63], dat_rsp_mask_val_fp16[61], dat_rsp_mask_val_fp16[59], dat_rsp_mask_val_fp16[57], dat_rsp_mask_val_fp16[55], dat_rsp_mask_val_fp16[53], dat_rsp_mask_val_fp16[51], dat_rsp_mask_val_fp16[49], dat_rsp_mask_val_fp16[47], dat_rsp_mask_val_fp16[45], dat_rsp_mask_val_fp16[43], dat_rsp_mask_val_fp16[41], dat_rsp_mask_val_fp16[39], dat_rsp_mask_val_fp16[37], dat_rsp_mask_val_fp16[35], dat_rsp_mask_val_fp16[33], dat_rsp_mask_val_fp16[31], dat_rsp_mask_val_fp16[29], dat_rsp_mask_val_fp16[27], dat_rsp_mask_val_fp16[25], dat_rsp_mask_val_fp16[23], dat_rsp_mask_val_fp16[21], dat_rsp_mask_val_fp16[19], dat_rsp_mask_val_fp16[17], dat_rsp_mask_val_fp16[15], dat_rsp_mask_val_fp16[13], dat_rsp_mask_val_fp16[11], dat_rsp_mask_val_fp16[9], dat_rsp_mask_val_fp16[7], dat_rsp_mask_val_fp16[5], dat_rsp_mask_val_fp16[3], dat_rsp_mask_val_fp16[1] };
  assign { dat_rsp_mask_val_int16[126], dat_rsp_mask_val_int16[124], dat_rsp_mask_val_int16[122], dat_rsp_mask_val_int16[120], dat_rsp_mask_val_int16[118], dat_rsp_mask_val_int16[116], dat_rsp_mask_val_int16[114], dat_rsp_mask_val_int16[112], dat_rsp_mask_val_int16[110], dat_rsp_mask_val_int16[108], dat_rsp_mask_val_int16[106], dat_rsp_mask_val_int16[104], dat_rsp_mask_val_int16[102], dat_rsp_mask_val_int16[100], dat_rsp_mask_val_int16[98], dat_rsp_mask_val_int16[96], dat_rsp_mask_val_int16[94], dat_rsp_mask_val_int16[92], dat_rsp_mask_val_int16[90], dat_rsp_mask_val_int16[88], dat_rsp_mask_val_int16[86], dat_rsp_mask_val_int16[84], dat_rsp_mask_val_int16[82], dat_rsp_mask_val_int16[80], dat_rsp_mask_val_int16[78], dat_rsp_mask_val_int16[76], dat_rsp_mask_val_int16[74], dat_rsp_mask_val_int16[72], dat_rsp_mask_val_int16[70], dat_rsp_mask_val_int16[68], dat_rsp_mask_val_int16[66], dat_rsp_mask_val_int16[64], dat_rsp_mask_val_int16[62], dat_rsp_mask_val_int16[60], dat_rsp_mask_val_int16[58], dat_rsp_mask_val_int16[56], dat_rsp_mask_val_int16[54], dat_rsp_mask_val_int16[52], dat_rsp_mask_val_int16[50], dat_rsp_mask_val_int16[48], dat_rsp_mask_val_int16[46], dat_rsp_mask_val_int16[44], dat_rsp_mask_val_int16[42], dat_rsp_mask_val_int16[40], dat_rsp_mask_val_int16[38], dat_rsp_mask_val_int16[36], dat_rsp_mask_val_int16[34], dat_rsp_mask_val_int16[32], dat_rsp_mask_val_int16[30], dat_rsp_mask_val_int16[28], dat_rsp_mask_val_int16[26], dat_rsp_mask_val_int16[24], dat_rsp_mask_val_int16[22], dat_rsp_mask_val_int16[20], dat_rsp_mask_val_int16[18], dat_rsp_mask_val_int16[16], dat_rsp_mask_val_int16[14], dat_rsp_mask_val_int16[12], dat_rsp_mask_val_int16[10], dat_rsp_mask_val_int16[8], dat_rsp_mask_val_int16[6], dat_rsp_mask_val_int16[4], dat_rsp_mask_val_int16[2], dat_rsp_mask_val_int16[0] } = { dat_rsp_mask_val_int16[127], dat_rsp_mask_val_int16[125], dat_rsp_mask_val_int16[123], dat_rsp_mask_val_int16[121], dat_rsp_mask_val_int16[119], dat_rsp_mask_val_int16[117], dat_rsp_mask_val_int16[115], dat_rsp_mask_val_int16[113], dat_rsp_mask_val_int16[111], dat_rsp_mask_val_int16[109], dat_rsp_mask_val_int16[107], dat_rsp_mask_val_int16[105], dat_rsp_mask_val_int16[103], dat_rsp_mask_val_int16[101], dat_rsp_mask_val_int16[99], dat_rsp_mask_val_int16[97], dat_rsp_mask_val_int16[95], dat_rsp_mask_val_int16[93], dat_rsp_mask_val_int16[91], dat_rsp_mask_val_int16[89], dat_rsp_mask_val_int16[87], dat_rsp_mask_val_int16[85], dat_rsp_mask_val_int16[83], dat_rsp_mask_val_int16[81], dat_rsp_mask_val_int16[79], dat_rsp_mask_val_int16[77], dat_rsp_mask_val_int16[75], dat_rsp_mask_val_int16[73], dat_rsp_mask_val_int16[71], dat_rsp_mask_val_int16[69], dat_rsp_mask_val_int16[67], dat_rsp_mask_val_int16[65], dat_rsp_mask_val_int16[63], dat_rsp_mask_val_int16[61], dat_rsp_mask_val_int16[59], dat_rsp_mask_val_int16[57], dat_rsp_mask_val_int16[55], dat_rsp_mask_val_int16[53], dat_rsp_mask_val_int16[51], dat_rsp_mask_val_int16[49], dat_rsp_mask_val_int16[47], dat_rsp_mask_val_int16[45], dat_rsp_mask_val_int16[43], dat_rsp_mask_val_int16[41], dat_rsp_mask_val_int16[39], dat_rsp_mask_val_int16[37], dat_rsp_mask_val_int16[35], dat_rsp_mask_val_int16[33], dat_rsp_mask_val_int16[31], dat_rsp_mask_val_int16[29], dat_rsp_mask_val_int16[27], dat_rsp_mask_val_int16[25], dat_rsp_mask_val_int16[23], dat_rsp_mask_val_int16[21], dat_rsp_mask_val_int16[19], dat_rsp_mask_val_int16[17], dat_rsp_mask_val_int16[15], dat_rsp_mask_val_int16[13], dat_rsp_mask_val_int16[11], dat_rsp_mask_val_int16[9], dat_rsp_mask_val_int16[7], dat_rsp_mask_val_int16[5], dat_rsp_mask_val_int16[3], dat_rsp_mask_val_int16[1] };
  assign dat_rsp_mask_w = dat_out_bypass_mask_w;
  assign dat_rsp_p0_vld_w = dat_out_bypass_p0_vld_w;
  assign dat_rsp_p1_vld_w = dat_out_bypass_p1_vld_w;
  assign dat_rsp_pd_d0 = { dat_rsp_pipe_pd_d6[28:19], dat_rsp_pipe_pd_d6[16:0] };
  assign dat_rsp_pipe_bytes = dat_rsp_pipe_pd_d6[14:7];
  assign dat_rsp_pipe_ch_end = dat_rsp_pipe_pd_d6[5];
  assign dat_rsp_pipe_ch_odd = dat_rsp_pipe_pd_d6[6];
  assign dat_rsp_pipe_cur_sub_h = dat_rsp_pipe_pd_d6[16:15];
  assign dat_rsp_pipe_dummy = dat_rsp_pipe_pd_d6[17];
  assign dat_rsp_pipe_flag = dat_rsp_pipe_pd_d6[28:20];
  assign dat_rsp_pipe_pd = dat_rsp_pipe_pd_d6;
  assign dat_rsp_pipe_pd_d0 = { dat_req_flag_d2, dat_req_rls_d2, dat_req_sub_w_st_d2, dat_req_dummy_d2, dat_req_cur_sub_h_d2, dat_req_bytes_d2, dat_req_ch_odd_d2, dat_req_ch_end_d2, dat_req_sub_c_d2, dat_req_sub_h_d2, dat_req_sub_w_d2 };
  assign dat_rsp_pipe_pvld = dat_rsp_pipe_pvld_d6;
  assign dat_rsp_pipe_pvld_d0 = dat_pipe_valid_d2;
  assign dat_rsp_pipe_rls = dat_rsp_pipe_pd_d6[19];
  assign dat_rsp_pipe_sub_c = dat_rsp_pipe_pd_d6[4];
  assign dat_rsp_pipe_sub_h = dat_rsp_pipe_pd_d6[3:2];
  assign dat_rsp_pipe_sub_w = dat_rsp_pipe_pd_d6[1:0];
  assign dat_rsp_pipe_sub_w_st = dat_rsp_pipe_pd_d6[18];
  assign dat_rsp_pra_en_d1[3:1] = { dat_rsp_pra_en_d1[0], dat_rsp_pra_en_d1[0], dat_rsp_pra_en_d1[0] };
  assign dat_rsp_pvld_d0 = dat_rsp_pipe_pvld_d6;
  assign dat_rsp_rls = dat_rsp_pd[17];
  assign dat_rsp_stripe_end = dat_rsp_pd[24];
  assign dat_rsp_stripe_st = dat_rsp_pd[23];
  assign dat_rsp_sub_c = dat_rsp_pd[4];
  assign dat_rsp_sub_h = dat_rsp_pd[3:2];
  assign dat_rsp_sub_w = dat_rsp_pd[1:0];
  assign dat_rsp_wg_lb = { dat_wg[2303:2048], dat_wg[1919:1664], dat_wg[1535:1280], dat_wg[1151:896] };
  assign dat_rsp_wg_lt = { dat_wg[1535:1280], dat_wg[1151:896], dat_wg[767:512], dat_wg[383:128] };
  assign dat_rsp_wg_rb = { dat_wg[2175:1920], dat_wg[1791:1536], dat_wg[1407:1152], dat_wg[1023:768] };
  assign dat_rsp_wg_rt = { dat_wg[1407:1152], dat_wg[1023:768], dat_wg[639:384], dat_wg[255:0] };
  assign dat_wg_16b_ch0 = { dat_rsp_wg[975:960], dat_rsp_wg[911:896], dat_rsp_wg[847:832], dat_rsp_wg[783:768], dat_rsp_wg[719:704], dat_rsp_wg[655:640], dat_rsp_wg[591:576], dat_rsp_wg[527:512], dat_rsp_wg[463:448], dat_rsp_wg[399:384], dat_rsp_wg[335:320], dat_rsp_wg[271:256], dat_rsp_wg[207:192], dat_rsp_wg[143:128], dat_rsp_wg[79:64], dat_rsp_wg[15:0] };
  assign dat_wg_16b_ch1 = { dat_rsp_wg[991:976], dat_rsp_wg[927:912], dat_rsp_wg[863:848], dat_rsp_wg[799:784], dat_rsp_wg[735:720], dat_rsp_wg[671:656], dat_rsp_wg[607:592], dat_rsp_wg[543:528], dat_rsp_wg[479:464], dat_rsp_wg[415:400], dat_rsp_wg[351:336], dat_rsp_wg[287:272], dat_rsp_wg[223:208], dat_rsp_wg[159:144], dat_rsp_wg[95:80], dat_rsp_wg[31:16] };
  assign dat_wg_16b_ch2 = { dat_rsp_wg[1007:992], dat_rsp_wg[943:928], dat_rsp_wg[879:864], dat_rsp_wg[815:800], dat_rsp_wg[751:736], dat_rsp_wg[687:672], dat_rsp_wg[623:608], dat_rsp_wg[559:544], dat_rsp_wg[495:480], dat_rsp_wg[431:416], dat_rsp_wg[367:352], dat_rsp_wg[303:288], dat_rsp_wg[239:224], dat_rsp_wg[175:160], dat_rsp_wg[111:96], dat_rsp_wg[47:32] };
  assign dat_wg_16b_ch3 = { dat_rsp_wg[1023:1008], dat_rsp_wg[959:944], dat_rsp_wg[895:880], dat_rsp_wg[831:816], dat_rsp_wg[767:752], dat_rsp_wg[703:688], dat_rsp_wg[639:624], dat_rsp_wg[575:560], dat_rsp_wg[511:496], dat_rsp_wg[447:432], dat_rsp_wg[383:368], dat_rsp_wg[319:304], dat_rsp_wg[255:240], dat_rsp_wg[191:176], dat_rsp_wg[127:112], dat_rsp_wg[63:48] };
  assign dat_wg_8b_ch0 = { dat_rsp_wg[967], dat_rsp_wg[967], dat_rsp_wg[967], dat_rsp_wg[967], dat_rsp_wg[967], dat_rsp_wg[967], dat_rsp_wg[967], dat_rsp_wg[967], dat_rsp_wg[967:960], dat_rsp_wg[903], dat_rsp_wg[903], dat_rsp_wg[903], dat_rsp_wg[903], dat_rsp_wg[903], dat_rsp_wg[903], dat_rsp_wg[903], dat_rsp_wg[903], dat_rsp_wg[903:896], dat_rsp_wg[839], dat_rsp_wg[839], dat_rsp_wg[839], dat_rsp_wg[839], dat_rsp_wg[839], dat_rsp_wg[839], dat_rsp_wg[839], dat_rsp_wg[839], dat_rsp_wg[839:832], dat_rsp_wg[775], dat_rsp_wg[775], dat_rsp_wg[775], dat_rsp_wg[775], dat_rsp_wg[775], dat_rsp_wg[775], dat_rsp_wg[775], dat_rsp_wg[775], dat_rsp_wg[775:768], dat_rsp_wg[711], dat_rsp_wg[711], dat_rsp_wg[711], dat_rsp_wg[711], dat_rsp_wg[711], dat_rsp_wg[711], dat_rsp_wg[711], dat_rsp_wg[711], dat_rsp_wg[711:704], dat_rsp_wg[647], dat_rsp_wg[647], dat_rsp_wg[647], dat_rsp_wg[647], dat_rsp_wg[647], dat_rsp_wg[647], dat_rsp_wg[647], dat_rsp_wg[647], dat_rsp_wg[647:640], dat_rsp_wg[583], dat_rsp_wg[583], dat_rsp_wg[583], dat_rsp_wg[583], dat_rsp_wg[583], dat_rsp_wg[583], dat_rsp_wg[583], dat_rsp_wg[583], dat_rsp_wg[583:576], dat_rsp_wg[519], dat_rsp_wg[519], dat_rsp_wg[519], dat_rsp_wg[519], dat_rsp_wg[519], dat_rsp_wg[519], dat_rsp_wg[519], dat_rsp_wg[519], dat_rsp_wg[519:512], dat_rsp_wg[455], dat_rsp_wg[455], dat_rsp_wg[455], dat_rsp_wg[455], dat_rsp_wg[455], dat_rsp_wg[455], dat_rsp_wg[455], dat_rsp_wg[455], dat_rsp_wg[455:448], dat_rsp_wg[391], dat_rsp_wg[391], dat_rsp_wg[391], dat_rsp_wg[391], dat_rsp_wg[391], dat_rsp_wg[391], dat_rsp_wg[391], dat_rsp_wg[391], dat_rsp_wg[391:384], dat_rsp_wg[327], dat_rsp_wg[327], dat_rsp_wg[327], dat_rsp_wg[327], dat_rsp_wg[327], dat_rsp_wg[327], dat_rsp_wg[327], dat_rsp_wg[327], dat_rsp_wg[327:320], dat_rsp_wg[263], dat_rsp_wg[263], dat_rsp_wg[263], dat_rsp_wg[263], dat_rsp_wg[263], dat_rsp_wg[263], dat_rsp_wg[263], dat_rsp_wg[263], dat_rsp_wg[263:256], dat_rsp_wg[199], dat_rsp_wg[199], dat_rsp_wg[199], dat_rsp_wg[199], dat_rsp_wg[199], dat_rsp_wg[199], dat_rsp_wg[199], dat_rsp_wg[199], dat_rsp_wg[199:192], dat_rsp_wg[135], dat_rsp_wg[135], dat_rsp_wg[135], dat_rsp_wg[135], dat_rsp_wg[135], dat_rsp_wg[135], dat_rsp_wg[135], dat_rsp_wg[135], dat_rsp_wg[135:128], dat_rsp_wg[71], dat_rsp_wg[71], dat_rsp_wg[71], dat_rsp_wg[71], dat_rsp_wg[71], dat_rsp_wg[71], dat_rsp_wg[71], dat_rsp_wg[71], dat_rsp_wg[71:64], dat_rsp_wg[7], dat_rsp_wg[7], dat_rsp_wg[7], dat_rsp_wg[7], dat_rsp_wg[7], dat_rsp_wg[7], dat_rsp_wg[7], dat_rsp_wg[7], dat_rsp_wg[7:0] };
  assign dat_wg_8b_ch1 = { dat_rsp_wg[975], dat_rsp_wg[975], dat_rsp_wg[975], dat_rsp_wg[975], dat_rsp_wg[975], dat_rsp_wg[975], dat_rsp_wg[975], dat_rsp_wg[975], dat_rsp_wg[975:968], dat_rsp_wg[911], dat_rsp_wg[911], dat_rsp_wg[911], dat_rsp_wg[911], dat_rsp_wg[911], dat_rsp_wg[911], dat_rsp_wg[911], dat_rsp_wg[911], dat_rsp_wg[911:904], dat_rsp_wg[847], dat_rsp_wg[847], dat_rsp_wg[847], dat_rsp_wg[847], dat_rsp_wg[847], dat_rsp_wg[847], dat_rsp_wg[847], dat_rsp_wg[847], dat_rsp_wg[847:840], dat_rsp_wg[783], dat_rsp_wg[783], dat_rsp_wg[783], dat_rsp_wg[783], dat_rsp_wg[783], dat_rsp_wg[783], dat_rsp_wg[783], dat_rsp_wg[783], dat_rsp_wg[783:776], dat_rsp_wg[719], dat_rsp_wg[719], dat_rsp_wg[719], dat_rsp_wg[719], dat_rsp_wg[719], dat_rsp_wg[719], dat_rsp_wg[719], dat_rsp_wg[719], dat_rsp_wg[719:712], dat_rsp_wg[655], dat_rsp_wg[655], dat_rsp_wg[655], dat_rsp_wg[655], dat_rsp_wg[655], dat_rsp_wg[655], dat_rsp_wg[655], dat_rsp_wg[655], dat_rsp_wg[655:648], dat_rsp_wg[591], dat_rsp_wg[591], dat_rsp_wg[591], dat_rsp_wg[591], dat_rsp_wg[591], dat_rsp_wg[591], dat_rsp_wg[591], dat_rsp_wg[591], dat_rsp_wg[591:584], dat_rsp_wg[527], dat_rsp_wg[527], dat_rsp_wg[527], dat_rsp_wg[527], dat_rsp_wg[527], dat_rsp_wg[527], dat_rsp_wg[527], dat_rsp_wg[527], dat_rsp_wg[527:520], dat_rsp_wg[463], dat_rsp_wg[463], dat_rsp_wg[463], dat_rsp_wg[463], dat_rsp_wg[463], dat_rsp_wg[463], dat_rsp_wg[463], dat_rsp_wg[463], dat_rsp_wg[463:456], dat_rsp_wg[399], dat_rsp_wg[399], dat_rsp_wg[399], dat_rsp_wg[399], dat_rsp_wg[399], dat_rsp_wg[399], dat_rsp_wg[399], dat_rsp_wg[399], dat_rsp_wg[399:392], dat_rsp_wg[335], dat_rsp_wg[335], dat_rsp_wg[335], dat_rsp_wg[335], dat_rsp_wg[335], dat_rsp_wg[335], dat_rsp_wg[335], dat_rsp_wg[335], dat_rsp_wg[335:328], dat_rsp_wg[271], dat_rsp_wg[271], dat_rsp_wg[271], dat_rsp_wg[271], dat_rsp_wg[271], dat_rsp_wg[271], dat_rsp_wg[271], dat_rsp_wg[271], dat_rsp_wg[271:264], dat_rsp_wg[207], dat_rsp_wg[207], dat_rsp_wg[207], dat_rsp_wg[207], dat_rsp_wg[207], dat_rsp_wg[207], dat_rsp_wg[207], dat_rsp_wg[207], dat_rsp_wg[207:200], dat_rsp_wg[143], dat_rsp_wg[143], dat_rsp_wg[143], dat_rsp_wg[143], dat_rsp_wg[143], dat_rsp_wg[143], dat_rsp_wg[143], dat_rsp_wg[143], dat_rsp_wg[143:136], dat_rsp_wg[79], dat_rsp_wg[79], dat_rsp_wg[79], dat_rsp_wg[79], dat_rsp_wg[79], dat_rsp_wg[79], dat_rsp_wg[79], dat_rsp_wg[79], dat_rsp_wg[79:72], dat_rsp_wg[15], dat_rsp_wg[15], dat_rsp_wg[15], dat_rsp_wg[15], dat_rsp_wg[15], dat_rsp_wg[15], dat_rsp_wg[15], dat_rsp_wg[15], dat_rsp_wg[15:8] };
  assign dat_wg_8b_ch2 = { dat_rsp_wg[983], dat_rsp_wg[983], dat_rsp_wg[983], dat_rsp_wg[983], dat_rsp_wg[983], dat_rsp_wg[983], dat_rsp_wg[983], dat_rsp_wg[983], dat_rsp_wg[983:976], dat_rsp_wg[919], dat_rsp_wg[919], dat_rsp_wg[919], dat_rsp_wg[919], dat_rsp_wg[919], dat_rsp_wg[919], dat_rsp_wg[919], dat_rsp_wg[919], dat_rsp_wg[919:912], dat_rsp_wg[855], dat_rsp_wg[855], dat_rsp_wg[855], dat_rsp_wg[855], dat_rsp_wg[855], dat_rsp_wg[855], dat_rsp_wg[855], dat_rsp_wg[855], dat_rsp_wg[855:848], dat_rsp_wg[791], dat_rsp_wg[791], dat_rsp_wg[791], dat_rsp_wg[791], dat_rsp_wg[791], dat_rsp_wg[791], dat_rsp_wg[791], dat_rsp_wg[791], dat_rsp_wg[791:784], dat_rsp_wg[727], dat_rsp_wg[727], dat_rsp_wg[727], dat_rsp_wg[727], dat_rsp_wg[727], dat_rsp_wg[727], dat_rsp_wg[727], dat_rsp_wg[727], dat_rsp_wg[727:720], dat_rsp_wg[663], dat_rsp_wg[663], dat_rsp_wg[663], dat_rsp_wg[663], dat_rsp_wg[663], dat_rsp_wg[663], dat_rsp_wg[663], dat_rsp_wg[663], dat_rsp_wg[663:656], dat_rsp_wg[599], dat_rsp_wg[599], dat_rsp_wg[599], dat_rsp_wg[599], dat_rsp_wg[599], dat_rsp_wg[599], dat_rsp_wg[599], dat_rsp_wg[599], dat_rsp_wg[599:592], dat_rsp_wg[535], dat_rsp_wg[535], dat_rsp_wg[535], dat_rsp_wg[535], dat_rsp_wg[535], dat_rsp_wg[535], dat_rsp_wg[535], dat_rsp_wg[535], dat_rsp_wg[535:528], dat_rsp_wg[471], dat_rsp_wg[471], dat_rsp_wg[471], dat_rsp_wg[471], dat_rsp_wg[471], dat_rsp_wg[471], dat_rsp_wg[471], dat_rsp_wg[471], dat_rsp_wg[471:464], dat_rsp_wg[407], dat_rsp_wg[407], dat_rsp_wg[407], dat_rsp_wg[407], dat_rsp_wg[407], dat_rsp_wg[407], dat_rsp_wg[407], dat_rsp_wg[407], dat_rsp_wg[407:400], dat_rsp_wg[343], dat_rsp_wg[343], dat_rsp_wg[343], dat_rsp_wg[343], dat_rsp_wg[343], dat_rsp_wg[343], dat_rsp_wg[343], dat_rsp_wg[343], dat_rsp_wg[343:336], dat_rsp_wg[279], dat_rsp_wg[279], dat_rsp_wg[279], dat_rsp_wg[279], dat_rsp_wg[279], dat_rsp_wg[279], dat_rsp_wg[279], dat_rsp_wg[279], dat_rsp_wg[279:272], dat_rsp_wg[215], dat_rsp_wg[215], dat_rsp_wg[215], dat_rsp_wg[215], dat_rsp_wg[215], dat_rsp_wg[215], dat_rsp_wg[215], dat_rsp_wg[215], dat_rsp_wg[215:208], dat_rsp_wg[151], dat_rsp_wg[151], dat_rsp_wg[151], dat_rsp_wg[151], dat_rsp_wg[151], dat_rsp_wg[151], dat_rsp_wg[151], dat_rsp_wg[151], dat_rsp_wg[151:144], dat_rsp_wg[87], dat_rsp_wg[87], dat_rsp_wg[87], dat_rsp_wg[87], dat_rsp_wg[87], dat_rsp_wg[87], dat_rsp_wg[87], dat_rsp_wg[87], dat_rsp_wg[87:80], dat_rsp_wg[23], dat_rsp_wg[23], dat_rsp_wg[23], dat_rsp_wg[23], dat_rsp_wg[23], dat_rsp_wg[23], dat_rsp_wg[23], dat_rsp_wg[23], dat_rsp_wg[23:16] };
  assign dat_wg_8b_ch3 = { dat_rsp_wg[991], dat_rsp_wg[991], dat_rsp_wg[991], dat_rsp_wg[991], dat_rsp_wg[991], dat_rsp_wg[991], dat_rsp_wg[991], dat_rsp_wg[991], dat_rsp_wg[991:984], dat_rsp_wg[927], dat_rsp_wg[927], dat_rsp_wg[927], dat_rsp_wg[927], dat_rsp_wg[927], dat_rsp_wg[927], dat_rsp_wg[927], dat_rsp_wg[927], dat_rsp_wg[927:920], dat_rsp_wg[863], dat_rsp_wg[863], dat_rsp_wg[863], dat_rsp_wg[863], dat_rsp_wg[863], dat_rsp_wg[863], dat_rsp_wg[863], dat_rsp_wg[863], dat_rsp_wg[863:856], dat_rsp_wg[799], dat_rsp_wg[799], dat_rsp_wg[799], dat_rsp_wg[799], dat_rsp_wg[799], dat_rsp_wg[799], dat_rsp_wg[799], dat_rsp_wg[799], dat_rsp_wg[799:792], dat_rsp_wg[735], dat_rsp_wg[735], dat_rsp_wg[735], dat_rsp_wg[735], dat_rsp_wg[735], dat_rsp_wg[735], dat_rsp_wg[735], dat_rsp_wg[735], dat_rsp_wg[735:728], dat_rsp_wg[671], dat_rsp_wg[671], dat_rsp_wg[671], dat_rsp_wg[671], dat_rsp_wg[671], dat_rsp_wg[671], dat_rsp_wg[671], dat_rsp_wg[671], dat_rsp_wg[671:664], dat_rsp_wg[607], dat_rsp_wg[607], dat_rsp_wg[607], dat_rsp_wg[607], dat_rsp_wg[607], dat_rsp_wg[607], dat_rsp_wg[607], dat_rsp_wg[607], dat_rsp_wg[607:600], dat_rsp_wg[543], dat_rsp_wg[543], dat_rsp_wg[543], dat_rsp_wg[543], dat_rsp_wg[543], dat_rsp_wg[543], dat_rsp_wg[543], dat_rsp_wg[543], dat_rsp_wg[543:536], dat_rsp_wg[479], dat_rsp_wg[479], dat_rsp_wg[479], dat_rsp_wg[479], dat_rsp_wg[479], dat_rsp_wg[479], dat_rsp_wg[479], dat_rsp_wg[479], dat_rsp_wg[479:472], dat_rsp_wg[415], dat_rsp_wg[415], dat_rsp_wg[415], dat_rsp_wg[415], dat_rsp_wg[415], dat_rsp_wg[415], dat_rsp_wg[415], dat_rsp_wg[415], dat_rsp_wg[415:408], dat_rsp_wg[351], dat_rsp_wg[351], dat_rsp_wg[351], dat_rsp_wg[351], dat_rsp_wg[351], dat_rsp_wg[351], dat_rsp_wg[351], dat_rsp_wg[351], dat_rsp_wg[351:344], dat_rsp_wg[287], dat_rsp_wg[287], dat_rsp_wg[287], dat_rsp_wg[287], dat_rsp_wg[287], dat_rsp_wg[287], dat_rsp_wg[287], dat_rsp_wg[287], dat_rsp_wg[287:280], dat_rsp_wg[223], dat_rsp_wg[223], dat_rsp_wg[223], dat_rsp_wg[223], dat_rsp_wg[223], dat_rsp_wg[223], dat_rsp_wg[223], dat_rsp_wg[223], dat_rsp_wg[223:216], dat_rsp_wg[159], dat_rsp_wg[159], dat_rsp_wg[159], dat_rsp_wg[159], dat_rsp_wg[159], dat_rsp_wg[159], dat_rsp_wg[159], dat_rsp_wg[159], dat_rsp_wg[159:152], dat_rsp_wg[95], dat_rsp_wg[95], dat_rsp_wg[95], dat_rsp_wg[95], dat_rsp_wg[95], dat_rsp_wg[95], dat_rsp_wg[95], dat_rsp_wg[95], dat_rsp_wg[95:88], dat_rsp_wg[31], dat_rsp_wg[31], dat_rsp_wg[31], dat_rsp_wg[31], dat_rsp_wg[31], dat_rsp_wg[31], dat_rsp_wg[31], dat_rsp_wg[31], dat_rsp_wg[31:24] };
  assign dat_wg_8b_ch4 = { dat_rsp_wg[999], dat_rsp_wg[999], dat_rsp_wg[999], dat_rsp_wg[999], dat_rsp_wg[999], dat_rsp_wg[999], dat_rsp_wg[999], dat_rsp_wg[999], dat_rsp_wg[999:992], dat_rsp_wg[935], dat_rsp_wg[935], dat_rsp_wg[935], dat_rsp_wg[935], dat_rsp_wg[935], dat_rsp_wg[935], dat_rsp_wg[935], dat_rsp_wg[935], dat_rsp_wg[935:928], dat_rsp_wg[871], dat_rsp_wg[871], dat_rsp_wg[871], dat_rsp_wg[871], dat_rsp_wg[871], dat_rsp_wg[871], dat_rsp_wg[871], dat_rsp_wg[871], dat_rsp_wg[871:864], dat_rsp_wg[807], dat_rsp_wg[807], dat_rsp_wg[807], dat_rsp_wg[807], dat_rsp_wg[807], dat_rsp_wg[807], dat_rsp_wg[807], dat_rsp_wg[807], dat_rsp_wg[807:800], dat_rsp_wg[743], dat_rsp_wg[743], dat_rsp_wg[743], dat_rsp_wg[743], dat_rsp_wg[743], dat_rsp_wg[743], dat_rsp_wg[743], dat_rsp_wg[743], dat_rsp_wg[743:736], dat_rsp_wg[679], dat_rsp_wg[679], dat_rsp_wg[679], dat_rsp_wg[679], dat_rsp_wg[679], dat_rsp_wg[679], dat_rsp_wg[679], dat_rsp_wg[679], dat_rsp_wg[679:672], dat_rsp_wg[615], dat_rsp_wg[615], dat_rsp_wg[615], dat_rsp_wg[615], dat_rsp_wg[615], dat_rsp_wg[615], dat_rsp_wg[615], dat_rsp_wg[615], dat_rsp_wg[615:608], dat_rsp_wg[551], dat_rsp_wg[551], dat_rsp_wg[551], dat_rsp_wg[551], dat_rsp_wg[551], dat_rsp_wg[551], dat_rsp_wg[551], dat_rsp_wg[551], dat_rsp_wg[551:544], dat_rsp_wg[487], dat_rsp_wg[487], dat_rsp_wg[487], dat_rsp_wg[487], dat_rsp_wg[487], dat_rsp_wg[487], dat_rsp_wg[487], dat_rsp_wg[487], dat_rsp_wg[487:480], dat_rsp_wg[423], dat_rsp_wg[423], dat_rsp_wg[423], dat_rsp_wg[423], dat_rsp_wg[423], dat_rsp_wg[423], dat_rsp_wg[423], dat_rsp_wg[423], dat_rsp_wg[423:416], dat_rsp_wg[359], dat_rsp_wg[359], dat_rsp_wg[359], dat_rsp_wg[359], dat_rsp_wg[359], dat_rsp_wg[359], dat_rsp_wg[359], dat_rsp_wg[359], dat_rsp_wg[359:352], dat_rsp_wg[295], dat_rsp_wg[295], dat_rsp_wg[295], dat_rsp_wg[295], dat_rsp_wg[295], dat_rsp_wg[295], dat_rsp_wg[295], dat_rsp_wg[295], dat_rsp_wg[295:288], dat_rsp_wg[231], dat_rsp_wg[231], dat_rsp_wg[231], dat_rsp_wg[231], dat_rsp_wg[231], dat_rsp_wg[231], dat_rsp_wg[231], dat_rsp_wg[231], dat_rsp_wg[231:224], dat_rsp_wg[167], dat_rsp_wg[167], dat_rsp_wg[167], dat_rsp_wg[167], dat_rsp_wg[167], dat_rsp_wg[167], dat_rsp_wg[167], dat_rsp_wg[167], dat_rsp_wg[167:160], dat_rsp_wg[103], dat_rsp_wg[103], dat_rsp_wg[103], dat_rsp_wg[103], dat_rsp_wg[103], dat_rsp_wg[103], dat_rsp_wg[103], dat_rsp_wg[103], dat_rsp_wg[103:96], dat_rsp_wg[39], dat_rsp_wg[39], dat_rsp_wg[39], dat_rsp_wg[39], dat_rsp_wg[39], dat_rsp_wg[39], dat_rsp_wg[39], dat_rsp_wg[39], dat_rsp_wg[39:32] };
  assign dat_wg_8b_ch5 = { dat_rsp_wg[1007], dat_rsp_wg[1007], dat_rsp_wg[1007], dat_rsp_wg[1007], dat_rsp_wg[1007], dat_rsp_wg[1007], dat_rsp_wg[1007], dat_rsp_wg[1007], dat_rsp_wg[1007:1000], dat_rsp_wg[943], dat_rsp_wg[943], dat_rsp_wg[943], dat_rsp_wg[943], dat_rsp_wg[943], dat_rsp_wg[943], dat_rsp_wg[943], dat_rsp_wg[943], dat_rsp_wg[943:936], dat_rsp_wg[879], dat_rsp_wg[879], dat_rsp_wg[879], dat_rsp_wg[879], dat_rsp_wg[879], dat_rsp_wg[879], dat_rsp_wg[879], dat_rsp_wg[879], dat_rsp_wg[879:872], dat_rsp_wg[815], dat_rsp_wg[815], dat_rsp_wg[815], dat_rsp_wg[815], dat_rsp_wg[815], dat_rsp_wg[815], dat_rsp_wg[815], dat_rsp_wg[815], dat_rsp_wg[815:808], dat_rsp_wg[751], dat_rsp_wg[751], dat_rsp_wg[751], dat_rsp_wg[751], dat_rsp_wg[751], dat_rsp_wg[751], dat_rsp_wg[751], dat_rsp_wg[751], dat_rsp_wg[751:744], dat_rsp_wg[687], dat_rsp_wg[687], dat_rsp_wg[687], dat_rsp_wg[687], dat_rsp_wg[687], dat_rsp_wg[687], dat_rsp_wg[687], dat_rsp_wg[687], dat_rsp_wg[687:680], dat_rsp_wg[623], dat_rsp_wg[623], dat_rsp_wg[623], dat_rsp_wg[623], dat_rsp_wg[623], dat_rsp_wg[623], dat_rsp_wg[623], dat_rsp_wg[623], dat_rsp_wg[623:616], dat_rsp_wg[559], dat_rsp_wg[559], dat_rsp_wg[559], dat_rsp_wg[559], dat_rsp_wg[559], dat_rsp_wg[559], dat_rsp_wg[559], dat_rsp_wg[559], dat_rsp_wg[559:552], dat_rsp_wg[495], dat_rsp_wg[495], dat_rsp_wg[495], dat_rsp_wg[495], dat_rsp_wg[495], dat_rsp_wg[495], dat_rsp_wg[495], dat_rsp_wg[495], dat_rsp_wg[495:488], dat_rsp_wg[431], dat_rsp_wg[431], dat_rsp_wg[431], dat_rsp_wg[431], dat_rsp_wg[431], dat_rsp_wg[431], dat_rsp_wg[431], dat_rsp_wg[431], dat_rsp_wg[431:424], dat_rsp_wg[367], dat_rsp_wg[367], dat_rsp_wg[367], dat_rsp_wg[367], dat_rsp_wg[367], dat_rsp_wg[367], dat_rsp_wg[367], dat_rsp_wg[367], dat_rsp_wg[367:360], dat_rsp_wg[303], dat_rsp_wg[303], dat_rsp_wg[303], dat_rsp_wg[303], dat_rsp_wg[303], dat_rsp_wg[303], dat_rsp_wg[303], dat_rsp_wg[303], dat_rsp_wg[303:296], dat_rsp_wg[239], dat_rsp_wg[239], dat_rsp_wg[239], dat_rsp_wg[239], dat_rsp_wg[239], dat_rsp_wg[239], dat_rsp_wg[239], dat_rsp_wg[239], dat_rsp_wg[239:232], dat_rsp_wg[175], dat_rsp_wg[175], dat_rsp_wg[175], dat_rsp_wg[175], dat_rsp_wg[175], dat_rsp_wg[175], dat_rsp_wg[175], dat_rsp_wg[175], dat_rsp_wg[175:168], dat_rsp_wg[111], dat_rsp_wg[111], dat_rsp_wg[111], dat_rsp_wg[111], dat_rsp_wg[111], dat_rsp_wg[111], dat_rsp_wg[111], dat_rsp_wg[111], dat_rsp_wg[111:104], dat_rsp_wg[47], dat_rsp_wg[47], dat_rsp_wg[47], dat_rsp_wg[47], dat_rsp_wg[47], dat_rsp_wg[47], dat_rsp_wg[47], dat_rsp_wg[47], dat_rsp_wg[47:40] };
  assign dat_wg_8b_ch6 = { dat_rsp_wg[1015], dat_rsp_wg[1015], dat_rsp_wg[1015], dat_rsp_wg[1015], dat_rsp_wg[1015], dat_rsp_wg[1015], dat_rsp_wg[1015], dat_rsp_wg[1015], dat_rsp_wg[1015:1008], dat_rsp_wg[951], dat_rsp_wg[951], dat_rsp_wg[951], dat_rsp_wg[951], dat_rsp_wg[951], dat_rsp_wg[951], dat_rsp_wg[951], dat_rsp_wg[951], dat_rsp_wg[951:944], dat_rsp_wg[887], dat_rsp_wg[887], dat_rsp_wg[887], dat_rsp_wg[887], dat_rsp_wg[887], dat_rsp_wg[887], dat_rsp_wg[887], dat_rsp_wg[887], dat_rsp_wg[887:880], dat_rsp_wg[823], dat_rsp_wg[823], dat_rsp_wg[823], dat_rsp_wg[823], dat_rsp_wg[823], dat_rsp_wg[823], dat_rsp_wg[823], dat_rsp_wg[823], dat_rsp_wg[823:816], dat_rsp_wg[759], dat_rsp_wg[759], dat_rsp_wg[759], dat_rsp_wg[759], dat_rsp_wg[759], dat_rsp_wg[759], dat_rsp_wg[759], dat_rsp_wg[759], dat_rsp_wg[759:752], dat_rsp_wg[695], dat_rsp_wg[695], dat_rsp_wg[695], dat_rsp_wg[695], dat_rsp_wg[695], dat_rsp_wg[695], dat_rsp_wg[695], dat_rsp_wg[695], dat_rsp_wg[695:688], dat_rsp_wg[631], dat_rsp_wg[631], dat_rsp_wg[631], dat_rsp_wg[631], dat_rsp_wg[631], dat_rsp_wg[631], dat_rsp_wg[631], dat_rsp_wg[631], dat_rsp_wg[631:624], dat_rsp_wg[567], dat_rsp_wg[567], dat_rsp_wg[567], dat_rsp_wg[567], dat_rsp_wg[567], dat_rsp_wg[567], dat_rsp_wg[567], dat_rsp_wg[567], dat_rsp_wg[567:560], dat_rsp_wg[503], dat_rsp_wg[503], dat_rsp_wg[503], dat_rsp_wg[503], dat_rsp_wg[503], dat_rsp_wg[503], dat_rsp_wg[503], dat_rsp_wg[503], dat_rsp_wg[503:496], dat_rsp_wg[439], dat_rsp_wg[439], dat_rsp_wg[439], dat_rsp_wg[439], dat_rsp_wg[439], dat_rsp_wg[439], dat_rsp_wg[439], dat_rsp_wg[439], dat_rsp_wg[439:432], dat_rsp_wg[375], dat_rsp_wg[375], dat_rsp_wg[375], dat_rsp_wg[375], dat_rsp_wg[375], dat_rsp_wg[375], dat_rsp_wg[375], dat_rsp_wg[375], dat_rsp_wg[375:368], dat_rsp_wg[311], dat_rsp_wg[311], dat_rsp_wg[311], dat_rsp_wg[311], dat_rsp_wg[311], dat_rsp_wg[311], dat_rsp_wg[311], dat_rsp_wg[311], dat_rsp_wg[311:304], dat_rsp_wg[247], dat_rsp_wg[247], dat_rsp_wg[247], dat_rsp_wg[247], dat_rsp_wg[247], dat_rsp_wg[247], dat_rsp_wg[247], dat_rsp_wg[247], dat_rsp_wg[247:240], dat_rsp_wg[183], dat_rsp_wg[183], dat_rsp_wg[183], dat_rsp_wg[183], dat_rsp_wg[183], dat_rsp_wg[183], dat_rsp_wg[183], dat_rsp_wg[183], dat_rsp_wg[183:176], dat_rsp_wg[119], dat_rsp_wg[119], dat_rsp_wg[119], dat_rsp_wg[119], dat_rsp_wg[119], dat_rsp_wg[119], dat_rsp_wg[119], dat_rsp_wg[119], dat_rsp_wg[119:112], dat_rsp_wg[55], dat_rsp_wg[55], dat_rsp_wg[55], dat_rsp_wg[55], dat_rsp_wg[55], dat_rsp_wg[55], dat_rsp_wg[55], dat_rsp_wg[55], dat_rsp_wg[55:48] };
  assign dat_wg_8b_ch7 = { dat_rsp_wg[1023], dat_rsp_wg[1023], dat_rsp_wg[1023], dat_rsp_wg[1023], dat_rsp_wg[1023], dat_rsp_wg[1023], dat_rsp_wg[1023], dat_rsp_wg[1023], dat_rsp_wg[1023:1016], dat_rsp_wg[959], dat_rsp_wg[959], dat_rsp_wg[959], dat_rsp_wg[959], dat_rsp_wg[959], dat_rsp_wg[959], dat_rsp_wg[959], dat_rsp_wg[959], dat_rsp_wg[959:952], dat_rsp_wg[895], dat_rsp_wg[895], dat_rsp_wg[895], dat_rsp_wg[895], dat_rsp_wg[895], dat_rsp_wg[895], dat_rsp_wg[895], dat_rsp_wg[895], dat_rsp_wg[895:888], dat_rsp_wg[831], dat_rsp_wg[831], dat_rsp_wg[831], dat_rsp_wg[831], dat_rsp_wg[831], dat_rsp_wg[831], dat_rsp_wg[831], dat_rsp_wg[831], dat_rsp_wg[831:824], dat_rsp_wg[767], dat_rsp_wg[767], dat_rsp_wg[767], dat_rsp_wg[767], dat_rsp_wg[767], dat_rsp_wg[767], dat_rsp_wg[767], dat_rsp_wg[767], dat_rsp_wg[767:760], dat_rsp_wg[703], dat_rsp_wg[703], dat_rsp_wg[703], dat_rsp_wg[703], dat_rsp_wg[703], dat_rsp_wg[703], dat_rsp_wg[703], dat_rsp_wg[703], dat_rsp_wg[703:696], dat_rsp_wg[639], dat_rsp_wg[639], dat_rsp_wg[639], dat_rsp_wg[639], dat_rsp_wg[639], dat_rsp_wg[639], dat_rsp_wg[639], dat_rsp_wg[639], dat_rsp_wg[639:632], dat_rsp_wg[575], dat_rsp_wg[575], dat_rsp_wg[575], dat_rsp_wg[575], dat_rsp_wg[575], dat_rsp_wg[575], dat_rsp_wg[575], dat_rsp_wg[575], dat_rsp_wg[575:568], dat_rsp_wg[511], dat_rsp_wg[511], dat_rsp_wg[511], dat_rsp_wg[511], dat_rsp_wg[511], dat_rsp_wg[511], dat_rsp_wg[511], dat_rsp_wg[511], dat_rsp_wg[511:504], dat_rsp_wg[447], dat_rsp_wg[447], dat_rsp_wg[447], dat_rsp_wg[447], dat_rsp_wg[447], dat_rsp_wg[447], dat_rsp_wg[447], dat_rsp_wg[447], dat_rsp_wg[447:440], dat_rsp_wg[383], dat_rsp_wg[383], dat_rsp_wg[383], dat_rsp_wg[383], dat_rsp_wg[383], dat_rsp_wg[383], dat_rsp_wg[383], dat_rsp_wg[383], dat_rsp_wg[383:376], dat_rsp_wg[319], dat_rsp_wg[319], dat_rsp_wg[319], dat_rsp_wg[319], dat_rsp_wg[319], dat_rsp_wg[319], dat_rsp_wg[319], dat_rsp_wg[319], dat_rsp_wg[319:312], dat_rsp_wg[255], dat_rsp_wg[255], dat_rsp_wg[255], dat_rsp_wg[255], dat_rsp_wg[255], dat_rsp_wg[255], dat_rsp_wg[255], dat_rsp_wg[255], dat_rsp_wg[255:248], dat_rsp_wg[191], dat_rsp_wg[191], dat_rsp_wg[191], dat_rsp_wg[191], dat_rsp_wg[191], dat_rsp_wg[191], dat_rsp_wg[191], dat_rsp_wg[191], dat_rsp_wg[191:184], dat_rsp_wg[127], dat_rsp_wg[127], dat_rsp_wg[127], dat_rsp_wg[127], dat_rsp_wg[127], dat_rsp_wg[127], dat_rsp_wg[127], dat_rsp_wg[127], dat_rsp_wg[127:120], dat_rsp_wg[63], dat_rsp_wg[63], dat_rsp_wg[63], dat_rsp_wg[63], dat_rsp_wg[63], dat_rsp_wg[63], dat_rsp_wg[63], dat_rsp_wg[63], dat_rsp_wg[63:56] };
  assign dat_wg_req_dummy = 1'b0;
  assign datain_c_cnt_reg_en = c_bias_reg_en;
  assign datain_height_cmp_w = reg2dp_datain_height_ext;
  assign datain_width_cmp_w = reg2dp_datain_width_ext;
  assign dataout_w_add = sub_h_cmp_g1;
  assign dataout_w_init[11:3] = { dataout_w_init[12], dataout_w_init[12], dataout_w_init[12], dataout_w_init[12], dataout_w_init[12], dataout_w_init[12], dataout_w_init[12], dataout_w_init[12], dataout_w_init[12] };
  assign dataout_w_ori_reg_en = datain_h_ori_reg_en;
  assign dataout_width_cmp_w = reg2dp_dataout_width;
  assign dl_block_end = dl_pd[26];
  assign dl_channel_end = dl_pd[27];
  assign dl_channel_size = dl_pd[16:10];
  assign dl_cur_sub_h = dl_pd[25:24];
  assign dl_dat_release = dl_pd[30];
  assign dl_group_end = dl_pd[28];
  assign dl_h_offset = dl_pd[9:5];
  assign dl_in_pd = dl_pd_d0;
  assign dl_in_pd_d0 = sg2dl_pd;
  assign dl_in_pvld_d0 = sg2dl_pvld;
  assign dl_layer_end = dl_pd[29];
  assign dl_out_pvld_d1 = sc2mac_dat_b_pvld;
  assign dl_pvld = dat_req_stripe_st;
  assign dl_pvld_d0 = dl_in_pvld;
  assign dl_stripe_length = dl_pd[23:17];
  assign dl_w_offset = dl_pd[4:0];
  assign h_bias_reg_en[0] = dat_exec_valid;
  assign is_pixel = reg2dp_datain_format;
  assign is_winograd = reg2dp_conv_mode;
  assign mon_batch_cnt_w = 1'bx;
  assign mon_c_bias_w = 1'bx;
  assign mon_datain_w_cnt_inc = 1'bx;
  assign mon_entries_w = 1'bx;
  assign mon_h_bias_3_w = 2'bxx;
  assign mon_pixel_w_cnt_w = 1'bx;
  assign mon_pixel_x_init_w = 2'bxx;
  assign mon_slice_left_w = 2'bxx;
  assign pixel_ch_stride_w = { pixel_x_stride_w, 6'b000000 };
  assign pixel_req_ch_odd_ori_en = pixel_ch_ori_reg_en;
  assign pixel_w_cur = pixel_w_cnt[15:6];
  assign pixel_w_ori_reg_en = pixel_req_ch_odd_en;
  assign pra_precision_0 = pra_precision[1:0];
  assign pra_precision_1 = pra_precision[3:2];
  assign pra_precision_2 = pra_precision[5:4];
  assign pra_precision_3 = pra_precision[7:6];
  assign pra_truncate_0 = pra_truncate[1:0];
  assign pra_truncate_1 = pra_truncate[3:2];
  assign pra_truncate_2 = pra_truncate[5:4];
  assign pra_truncate_3 = pra_truncate[7:6];
  assign reuse_rls = sg2dl_reuse_rls;
  assign sc2mac_dat_a_pvld = sc2mac_dat_b_pvld;
  assign slcg_wg_en = slcg_wg_en_d3;
  assign w_bias_reg_en = dat_exec_valid;
endmodule
