module exp(clk, rst, in, out);
  reg out;
  input clk;
  input rst;
  input in;
  output out;
endmodule
