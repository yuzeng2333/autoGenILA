module SDP_X_leading_sign_23_0(mantissa, rtn);
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:287" *)
  wire _000_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:295" *)
  wire _001_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:298" *)
  wire _002_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:299" *)
  wire _003_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:299" *)
  wire _004_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:300" *)
  wire _005_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:301" *)
  wire _006_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:301" *)
  wire _007_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:304" *)
  wire _008_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:304" *)
  wire _009_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:305" *)
  wire _010_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:305" *)
  wire _011_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:305" *)
  wire _012_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:306" *)
  wire _013_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:307" *)
  wire _014_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:307" *)
  wire _015_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:307" *)
  wire _016_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:307" *)
  wire _017_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:308" *)
  wire _018_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:308" *)
  wire _019_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:308" *)
  wire _020_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:279" *)
  wire _021_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:286" *)
  wire _022_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:306" *)
  wire _023_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:275" *)
  wire _024_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:276" *)
  wire _025_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:277" *)
  wire _026_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:281" *)
  wire _027_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:282" *)
  wire _028_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:283" *)
  wire _029_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:288" *)
  wire _030_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:289" *)
  wire _031_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:290" *)
  wire _032_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:303" *)
  wire _033_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:304" *)
  wire _034_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:304" *)
  wire _035_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:305" *)
  wire _036_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:306" *)
  wire _037_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:293" *)
  wire _038_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:295" *)
  wire _039_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:295" *)
  wire _040_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:299" *)
  wire _041_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:299" *)
  wire _042_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:301" *)
  wire _043_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:301" *)
  wire _044_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:303" *)
  wire _045_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:303" *)
  wire _046_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:304" *)
  wire _047_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:304" *)
  wire _048_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:304" *)
  wire _049_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:304" *)
  wire _050_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:305" *)
  wire _051_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:305" *)
  wire _052_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:305" *)
  wire _053_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:305" *)
  wire _054_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:306" *)
  wire _055_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:306" *)
  wire _056_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:306" *)
  wire _057_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:307" *)
  wire _058_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:307" *)
  wire _059_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:307" *)
  wire _060_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:307" *)
  wire _061_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:295" *)
  wire _062_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:295" *)
  wire _063_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:297" *)
  wire _064_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:299" *)
  wire _065_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:301" *)
  wire _066_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:303" *)
  wire _067_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:304" *)
  wire _068_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:304" *)
  wire _069_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:305" *)
  wire _070_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:306" *)
  wire _071_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:273" *)
  wire IntLeadZero_23U_leading_sign_23_0_rtn_IntLeadZero_23U_leading_sign_23_0_rtn_or_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:271" *)
  wire IntLeadZero_23U_leading_sign_23_0_rtn_and_83_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:270" *)
  wire IntLeadZero_23U_leading_sign_23_0_rtn_and_85_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:272" *)
  wire IntLeadZero_23U_leading_sign_23_0_rtn_and_90_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:260" *)
  wire IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_14_2_sdt_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:255" *)
  wire IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_18_3_sdt_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:261" *)
  wire IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_26_2_sdt_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:256" *)
  wire IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_26_2_sdt_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:262" *)
  wire IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_34_2_sdt_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:257" *)
  wire IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_42_4_sdt_4;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:263" *)
  wire IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_50_2_sdt_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:258" *)
  wire IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_50_2_sdt_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:264" *)
  wire IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_56_2_sdt_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:259" *)
  wire IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_6_2_sdt_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:254" *)
  wire IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_6_2_sdt_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:269" *)
  wire c_h_1_10;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:265" *)
  wire c_h_1_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:266" *)
  wire c_h_1_5;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:267" *)
  wire c_h_1_6;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:268" *)
  wire c_h_1_9;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:251" *)
  input [22:0] mantissa;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:252" *)
  output [4:0] rtn;
  assign c_h_1_2 = IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_6_2_sdt_1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:278" *) IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_6_2_sdt_2;
  assign IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_18_3_sdt_3 = _021_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:280" *) IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_14_2_sdt_1;
  assign c_h_1_5 = IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_26_2_sdt_1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:284" *) IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_26_2_sdt_2;
  assign c_h_1_6 = c_h_1_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:285" *) IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_18_3_sdt_3;
  assign _000_ = _022_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:287" *) IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_34_2_sdt_1;
  assign IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_42_4_sdt_4 = _000_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:287" *) c_h_1_5;
  assign c_h_1_9 = IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_50_2_sdt_1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:291" *) IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_50_2_sdt_2;
  assign c_h_1_10 = c_h_1_6 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:292" *) IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_42_4_sdt_4;
  assign IntLeadZero_23U_leading_sign_23_0_rtn_and_85_nl = c_h_1_6 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:293" *) _038_;
  assign _001_ = c_h_1_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:295" *) _062_;
  assign IntLeadZero_23U_leading_sign_23_0_rtn_and_83_nl = _001_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:295" *) _063_;
  assign _002_ = IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_6_2_sdt_1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:298" *) _064_;
  assign _003_ = IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_26_2_sdt_1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:299" *) _065_;
  assign _004_ = _041_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:299" *) c_h_1_6;
  assign _005_ = _002_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:300" *) _042_;
  assign _006_ = IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_50_2_sdt_1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:301" *) _066_;
  assign _007_ = _043_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:301" *) c_h_1_10;
  assign IntLeadZero_23U_leading_sign_23_0_rtn_and_90_nl = _005_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:301" *) _044_;
  assign _008_ = _068_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:304" *) c_h_1_2;
  assign _009_ = _046_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:304" *) _048_;
  assign _010_ = _070_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:305" *) c_h_1_5;
  assign _011_ = _050_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:305" *) _052_;
  assign _012_ = _053_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:305" *) c_h_1_6;
  assign _013_ = _009_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:306" *) _054_;
  assign _014_ = _057_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:307" *) c_h_1_9;
  assign _015_ = _056_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:307" *) _058_;
  assign _016_ = _059_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:307" *) c_h_1_10;
  assign _017_ = _013_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:307" *) _060_;
  assign _018_ = _061_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:308" *) IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_56_2_sdt_1;
  assign _019_ = _018_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:308" *) c_h_1_9;
  assign _020_ = _019_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:308" *) c_h_1_10;
  assign _021_ = ! (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:279" *) mantissa[16:15];
  assign _022_ = ! (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:286" *) mantissa[8:7];
  assign _023_ = mantissa[2:1] == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:306" *) 1'b1;
  assign _024_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:275" *) mantissa[20:19];
  assign _025_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:276" *) mantissa[22:21];
  assign _026_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:277" *) mantissa[18:17];
  assign _027_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:281" *) mantissa[12:11];
  assign _028_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:282" *) mantissa[14:13];
  assign _029_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:283" *) mantissa[10:9];
  assign _030_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:288" *) mantissa[4:3];
  assign _031_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:289" *) mantissa[6:5];
  assign _032_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:290" *) mantissa[2:1];
  assign _033_ = mantissa[21:20] != (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:303" *) 1'b1;
  assign _034_ = mantissa[17:16] != (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:304" *) 1'b1;
  assign _035_ = mantissa[13:12] != (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:304" *) 1'b1;
  assign _036_ = mantissa[9:8] != (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:305" *) 1'b1;
  assign _037_ = mantissa[5:4] != (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:306" *) 1'b1;
  assign IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_6_2_sdt_2 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:275" *) _024_;
  assign IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_6_2_sdt_1 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:276" *) _025_;
  assign IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_14_2_sdt_1 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:277" *) _026_;
  assign IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_26_2_sdt_2 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:281" *) _027_;
  assign IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_26_2_sdt_1 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:282" *) _028_;
  assign IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_34_2_sdt_1 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:283" *) _029_;
  assign IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_50_2_sdt_2 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:288" *) _030_;
  assign IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_50_2_sdt_1 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:289" *) _031_;
  assign IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_56_2_sdt_1 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:290" *) _032_;
  assign _038_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:293" *) IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_42_4_sdt_4;
  assign _039_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:295" *) IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_18_3_sdt_3;
  assign _040_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:295" *) c_h_1_10;
  assign _041_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:299" *) _003_;
  assign _042_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:299" *) _004_;
  assign _043_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:301" *) _006_;
  assign _044_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:301" *) _007_;
  assign _045_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:303" *) _033_;
  assign _046_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:303" *) _067_;
  assign _047_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:304" *) _034_;
  assign _048_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:304" *) _008_;
  assign _049_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:304" *) _035_;
  assign _050_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:304" *) _069_;
  assign _051_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:305" *) _036_;
  assign _052_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:305" *) _010_;
  assign _053_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:305" *) _011_;
  assign _054_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:305" *) _012_;
  assign _055_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:306" *) _037_;
  assign _056_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:306" *) _071_;
  assign _057_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:306" *) _023_;
  assign _058_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:307" *) _014_;
  assign _059_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:307" *) _015_;
  assign _060_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:307" *) _016_;
  assign _061_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:307" *) mantissa[0];
  assign _062_ = c_h_1_5 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:295" *) _039_;
  assign _063_ = c_h_1_9 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:295" *) _040_;
  assign _064_ = IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_14_2_sdt_1 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:297" *) _024_;
  assign _065_ = IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_34_2_sdt_1 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:299" *) _027_;
  assign _066_ = IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_56_2_sdt_1 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:301" *) _030_;
  assign _067_ = mantissa[22] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:303" *) _045_;
  assign _068_ = mantissa[18] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:304" *) _047_;
  assign _069_ = mantissa[14] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:304" *) _049_;
  assign _070_ = mantissa[10] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:305" *) _051_;
  assign _071_ = mantissa[6] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:306" *) _055_;
  assign IntLeadZero_23U_leading_sign_23_0_rtn_IntLeadZero_23U_leading_sign_23_0_rtn_or_2_nl = _017_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:308" *) _020_;
  assign rtn = { c_h_1_10, IntLeadZero_23U_leading_sign_23_0_rtn_and_85_nl, IntLeadZero_23U_leading_sign_23_0_rtn_and_83_nl, IntLeadZero_23U_leading_sign_23_0_rtn_and_90_nl, IntLeadZero_23U_leading_sign_23_0_rtn_IntLeadZero_23U_leading_sign_23_0_rtn_or_2_nl };
endmodule
