module expand_key_128(clk, in, out_1, out_2, rcon);
  (* src = "expand_key_128.v:28|S4.v:26|S.v:11" *)
  wire [7:0] _0000_;
  wire _0001_;
  wire _0002_;
  wire _0003_;
  wire _0004_;
  wire _0005_;
  wire _0006_;
  wire _0007_;
  wire _0008_;
  wire _0009_;
  wire _0010_;
  wire _0011_;
  wire _0012_;
  wire _0013_;
  wire _0014_;
  wire _0015_;
  wire _0016_;
  wire _0017_;
  wire _0018_;
  wire _0019_;
  wire _0020_;
  wire _0021_;
  wire _0022_;
  wire _0023_;
  wire _0024_;
  wire _0025_;
  wire _0026_;
  wire _0027_;
  wire _0028_;
  wire _0029_;
  wire _0030_;
  wire _0031_;
  wire _0032_;
  wire _0033_;
  wire _0034_;
  wire _0035_;
  wire _0036_;
  wire _0037_;
  wire _0038_;
  wire _0039_;
  wire _0040_;
  wire _0041_;
  wire _0042_;
  wire _0043_;
  wire _0044_;
  wire _0045_;
  wire _0046_;
  wire _0047_;
  wire _0048_;
  wire _0049_;
  wire _0050_;
  wire _0051_;
  wire _0052_;
  wire _0053_;
  wire _0054_;
  wire _0055_;
  wire _0056_;
  wire _0057_;
  wire _0058_;
  wire _0059_;
  wire _0060_;
  wire _0061_;
  wire _0062_;
  wire _0063_;
  wire _0064_;
  wire _0065_;
  wire _0066_;
  wire _0067_;
  wire _0068_;
  wire _0069_;
  wire _0070_;
  wire _0071_;
  wire _0072_;
  wire _0073_;
  wire _0074_;
  wire _0075_;
  wire _0076_;
  wire _0077_;
  wire _0078_;
  wire _0079_;
  wire _0080_;
  wire _0081_;
  wire _0082_;
  wire _0083_;
  wire _0084_;
  wire _0085_;
  wire _0086_;
  wire _0087_;
  wire _0088_;
  wire _0089_;
  wire _0090_;
  wire _0091_;
  wire _0092_;
  wire _0093_;
  wire _0094_;
  wire _0095_;
  wire _0096_;
  wire _0097_;
  wire _0098_;
  wire _0099_;
  wire _0100_;
  wire _0101_;
  wire _0102_;
  wire _0103_;
  wire _0104_;
  wire _0105_;
  wire _0106_;
  wire _0107_;
  wire _0108_;
  wire _0109_;
  wire _0110_;
  wire _0111_;
  wire _0112_;
  wire _0113_;
  wire _0114_;
  wire _0115_;
  wire _0116_;
  wire _0117_;
  wire _0118_;
  wire _0119_;
  wire _0120_;
  wire _0121_;
  wire _0122_;
  wire _0123_;
  wire _0124_;
  wire _0125_;
  wire _0126_;
  wire _0127_;
  wire _0128_;
  wire _0129_;
  wire _0130_;
  wire _0131_;
  wire _0132_;
  wire _0133_;
  wire _0134_;
  wire _0135_;
  wire _0136_;
  wire _0137_;
  wire _0138_;
  wire _0139_;
  wire _0140_;
  wire _0141_;
  wire _0142_;
  wire _0143_;
  wire _0144_;
  wire _0145_;
  wire _0146_;
  wire _0147_;
  wire _0148_;
  wire _0149_;
  wire _0150_;
  wire _0151_;
  wire _0152_;
  wire _0153_;
  wire _0154_;
  wire _0155_;
  wire _0156_;
  wire _0157_;
  wire _0158_;
  wire _0159_;
  wire _0160_;
  wire _0161_;
  wire _0162_;
  wire _0163_;
  wire _0164_;
  wire _0165_;
  wire _0166_;
  wire _0167_;
  wire _0168_;
  wire _0169_;
  wire _0170_;
  wire _0171_;
  wire _0172_;
  wire _0173_;
  wire _0174_;
  wire _0175_;
  wire _0176_;
  wire _0177_;
  wire _0178_;
  wire _0179_;
  wire _0180_;
  wire _0181_;
  wire _0182_;
  wire _0183_;
  wire _0184_;
  wire _0185_;
  wire _0186_;
  wire _0187_;
  wire _0188_;
  wire _0189_;
  wire _0190_;
  wire _0191_;
  wire _0192_;
  wire _0193_;
  wire _0194_;
  wire _0195_;
  wire _0196_;
  wire _0197_;
  wire _0198_;
  wire _0199_;
  wire _0200_;
  wire _0201_;
  wire _0202_;
  wire _0203_;
  wire _0204_;
  wire _0205_;
  wire _0206_;
  wire _0207_;
  wire _0208_;
  wire _0209_;
  wire _0210_;
  wire _0211_;
  wire _0212_;
  wire _0213_;
  wire _0214_;
  wire _0215_;
  wire _0216_;
  wire _0217_;
  wire _0218_;
  wire _0219_;
  wire _0220_;
  wire _0221_;
  wire _0222_;
  wire _0223_;
  wire _0224_;
  wire _0225_;
  wire _0226_;
  wire _0227_;
  wire _0228_;
  wire _0229_;
  wire _0230_;
  wire _0231_;
  wire _0232_;
  wire _0233_;
  wire _0234_;
  wire _0235_;
  wire _0236_;
  wire _0237_;
  wire _0238_;
  wire _0239_;
  wire _0240_;
  wire _0241_;
  wire _0242_;
  wire _0243_;
  wire _0244_;
  wire _0245_;
  wire _0246_;
  wire _0247_;
  wire _0248_;
  wire _0249_;
  wire _0250_;
  wire _0251_;
  wire _0252_;
  wire _0253_;
  wire _0254_;
  wire _0255_;
  wire _0256_;
  (* src = "expand_key_128.v:28|S4.v:26|S.v:11" *)
  wire [7:0] _0257_;
  wire _0258_;
  wire _0259_;
  wire _0260_;
  wire _0261_;
  wire _0262_;
  wire _0263_;
  wire _0264_;
  wire _0265_;
  wire _0266_;
  wire _0267_;
  wire _0268_;
  wire _0269_;
  wire _0270_;
  wire _0271_;
  wire _0272_;
  wire _0273_;
  wire _0274_;
  wire _0275_;
  wire _0276_;
  wire _0277_;
  wire _0278_;
  wire _0279_;
  wire _0280_;
  wire _0281_;
  wire _0282_;
  wire _0283_;
  wire _0284_;
  wire _0285_;
  wire _0286_;
  wire _0287_;
  wire _0288_;
  wire _0289_;
  wire _0290_;
  wire _0291_;
  wire _0292_;
  wire _0293_;
  wire _0294_;
  wire _0295_;
  wire _0296_;
  wire _0297_;
  wire _0298_;
  wire _0299_;
  wire _0300_;
  wire _0301_;
  wire _0302_;
  wire _0303_;
  wire _0304_;
  wire _0305_;
  wire _0306_;
  wire _0307_;
  wire _0308_;
  wire _0309_;
  wire _0310_;
  wire _0311_;
  wire _0312_;
  wire _0313_;
  wire _0314_;
  wire _0315_;
  wire _0316_;
  wire _0317_;
  wire _0318_;
  wire _0319_;
  wire _0320_;
  wire _0321_;
  wire _0322_;
  wire _0323_;
  wire _0324_;
  wire _0325_;
  wire _0326_;
  wire _0327_;
  wire _0328_;
  wire _0329_;
  wire _0330_;
  wire _0331_;
  wire _0332_;
  wire _0333_;
  wire _0334_;
  wire _0335_;
  wire _0336_;
  wire _0337_;
  wire _0338_;
  wire _0339_;
  wire _0340_;
  wire _0341_;
  wire _0342_;
  wire _0343_;
  wire _0344_;
  wire _0345_;
  wire _0346_;
  wire _0347_;
  wire _0348_;
  wire _0349_;
  wire _0350_;
  wire _0351_;
  wire _0352_;
  wire _0353_;
  wire _0354_;
  wire _0355_;
  wire _0356_;
  wire _0357_;
  wire _0358_;
  wire _0359_;
  wire _0360_;
  wire _0361_;
  wire _0362_;
  wire _0363_;
  wire _0364_;
  wire _0365_;
  wire _0366_;
  wire _0367_;
  wire _0368_;
  wire _0369_;
  wire _0370_;
  wire _0371_;
  wire _0372_;
  wire _0373_;
  wire _0374_;
  wire _0375_;
  wire _0376_;
  wire _0377_;
  wire _0378_;
  wire _0379_;
  wire _0380_;
  wire _0381_;
  wire _0382_;
  wire _0383_;
  wire _0384_;
  wire _0385_;
  wire _0386_;
  wire _0387_;
  wire _0388_;
  wire _0389_;
  wire _0390_;
  wire _0391_;
  wire _0392_;
  wire _0393_;
  wire _0394_;
  wire _0395_;
  wire _0396_;
  wire _0397_;
  wire _0398_;
  wire _0399_;
  wire _0400_;
  wire _0401_;
  wire _0402_;
  wire _0403_;
  wire _0404_;
  wire _0405_;
  wire _0406_;
  wire _0407_;
  wire _0408_;
  wire _0409_;
  wire _0410_;
  wire _0411_;
  wire _0412_;
  wire _0413_;
  wire _0414_;
  wire _0415_;
  wire _0416_;
  wire _0417_;
  wire _0418_;
  wire _0419_;
  wire _0420_;
  wire _0421_;
  wire _0422_;
  wire _0423_;
  wire _0424_;
  wire _0425_;
  wire _0426_;
  wire _0427_;
  wire _0428_;
  wire _0429_;
  wire _0430_;
  wire _0431_;
  wire _0432_;
  wire _0433_;
  wire _0434_;
  wire _0435_;
  wire _0436_;
  wire _0437_;
  wire _0438_;
  wire _0439_;
  wire _0440_;
  wire _0441_;
  wire _0442_;
  wire _0443_;
  wire _0444_;
  wire _0445_;
  wire _0446_;
  wire _0447_;
  wire _0448_;
  wire _0449_;
  wire _0450_;
  wire _0451_;
  wire _0452_;
  wire _0453_;
  wire _0454_;
  wire _0455_;
  wire _0456_;
  wire _0457_;
  wire _0458_;
  wire _0459_;
  wire _0460_;
  wire _0461_;
  wire _0462_;
  wire _0463_;
  wire _0464_;
  wire _0465_;
  wire _0466_;
  wire _0467_;
  wire _0468_;
  wire _0469_;
  wire _0470_;
  wire _0471_;
  wire _0472_;
  wire _0473_;
  wire _0474_;
  wire _0475_;
  wire _0476_;
  wire _0477_;
  wire _0478_;
  wire _0479_;
  wire _0480_;
  wire _0481_;
  wire _0482_;
  wire _0483_;
  wire _0484_;
  wire _0485_;
  wire _0486_;
  wire _0487_;
  wire _0488_;
  wire _0489_;
  wire _0490_;
  wire _0491_;
  wire _0492_;
  wire _0493_;
  wire _0494_;
  wire _0495_;
  wire _0496_;
  wire _0497_;
  wire _0498_;
  wire _0499_;
  wire _0500_;
  wire _0501_;
  wire _0502_;
  wire _0503_;
  wire _0504_;
  wire _0505_;
  wire _0506_;
  wire _0507_;
  wire _0508_;
  wire _0509_;
  wire _0510_;
  wire _0511_;
  wire _0512_;
  wire _0513_;
  (* src = "expand_key_128.v:28|S4.v:26|S.v:11" *)
  wire [7:0] _0514_;
  wire _0515_;
  wire _0516_;
  wire _0517_;
  wire _0518_;
  wire _0519_;
  wire _0520_;
  wire _0521_;
  wire _0522_;
  wire _0523_;
  wire _0524_;
  wire _0525_;
  wire _0526_;
  wire _0527_;
  wire _0528_;
  wire _0529_;
  wire _0530_;
  wire _0531_;
  wire _0532_;
  wire _0533_;
  wire _0534_;
  wire _0535_;
  wire _0536_;
  wire _0537_;
  wire _0538_;
  wire _0539_;
  wire _0540_;
  wire _0541_;
  wire _0542_;
  wire _0543_;
  wire _0544_;
  wire _0545_;
  wire _0546_;
  wire _0547_;
  wire _0548_;
  wire _0549_;
  wire _0550_;
  wire _0551_;
  wire _0552_;
  wire _0553_;
  wire _0554_;
  wire _0555_;
  wire _0556_;
  wire _0557_;
  wire _0558_;
  wire _0559_;
  wire _0560_;
  wire _0561_;
  wire _0562_;
  wire _0563_;
  wire _0564_;
  wire _0565_;
  wire _0566_;
  wire _0567_;
  wire _0568_;
  wire _0569_;
  wire _0570_;
  wire _0571_;
  wire _0572_;
  wire _0573_;
  wire _0574_;
  wire _0575_;
  wire _0576_;
  wire _0577_;
  wire _0578_;
  wire _0579_;
  wire _0580_;
  wire _0581_;
  wire _0582_;
  wire _0583_;
  wire _0584_;
  wire _0585_;
  wire _0586_;
  wire _0587_;
  wire _0588_;
  wire _0589_;
  wire _0590_;
  wire _0591_;
  wire _0592_;
  wire _0593_;
  wire _0594_;
  wire _0595_;
  wire _0596_;
  wire _0597_;
  wire _0598_;
  wire _0599_;
  wire _0600_;
  wire _0601_;
  wire _0602_;
  wire _0603_;
  wire _0604_;
  wire _0605_;
  wire _0606_;
  wire _0607_;
  wire _0608_;
  wire _0609_;
  wire _0610_;
  wire _0611_;
  wire _0612_;
  wire _0613_;
  wire _0614_;
  wire _0615_;
  wire _0616_;
  wire _0617_;
  wire _0618_;
  wire _0619_;
  wire _0620_;
  wire _0621_;
  wire _0622_;
  wire _0623_;
  wire _0624_;
  wire _0625_;
  wire _0626_;
  wire _0627_;
  wire _0628_;
  wire _0629_;
  wire _0630_;
  wire _0631_;
  wire _0632_;
  wire _0633_;
  wire _0634_;
  wire _0635_;
  wire _0636_;
  wire _0637_;
  wire _0638_;
  wire _0639_;
  wire _0640_;
  wire _0641_;
  wire _0642_;
  wire _0643_;
  wire _0644_;
  wire _0645_;
  wire _0646_;
  wire _0647_;
  wire _0648_;
  wire _0649_;
  wire _0650_;
  wire _0651_;
  wire _0652_;
  wire _0653_;
  wire _0654_;
  wire _0655_;
  wire _0656_;
  wire _0657_;
  wire _0658_;
  wire _0659_;
  wire _0660_;
  wire _0661_;
  wire _0662_;
  wire _0663_;
  wire _0664_;
  wire _0665_;
  wire _0666_;
  wire _0667_;
  wire _0668_;
  wire _0669_;
  wire _0670_;
  wire _0671_;
  wire _0672_;
  wire _0673_;
  wire _0674_;
  wire _0675_;
  wire _0676_;
  wire _0677_;
  wire _0678_;
  wire _0679_;
  wire _0680_;
  wire _0681_;
  wire _0682_;
  wire _0683_;
  wire _0684_;
  wire _0685_;
  wire _0686_;
  wire _0687_;
  wire _0688_;
  wire _0689_;
  wire _0690_;
  wire _0691_;
  wire _0692_;
  wire _0693_;
  wire _0694_;
  wire _0695_;
  wire _0696_;
  wire _0697_;
  wire _0698_;
  wire _0699_;
  wire _0700_;
  wire _0701_;
  wire _0702_;
  wire _0703_;
  wire _0704_;
  wire _0705_;
  wire _0706_;
  wire _0707_;
  wire _0708_;
  wire _0709_;
  wire _0710_;
  wire _0711_;
  wire _0712_;
  wire _0713_;
  wire _0714_;
  wire _0715_;
  wire _0716_;
  wire _0717_;
  wire _0718_;
  wire _0719_;
  wire _0720_;
  wire _0721_;
  wire _0722_;
  wire _0723_;
  wire _0724_;
  wire _0725_;
  wire _0726_;
  wire _0727_;
  wire _0728_;
  wire _0729_;
  wire _0730_;
  wire _0731_;
  wire _0732_;
  wire _0733_;
  wire _0734_;
  wire _0735_;
  wire _0736_;
  wire _0737_;
  wire _0738_;
  wire _0739_;
  wire _0740_;
  wire _0741_;
  wire _0742_;
  wire _0743_;
  wire _0744_;
  wire _0745_;
  wire _0746_;
  wire _0747_;
  wire _0748_;
  wire _0749_;
  wire _0750_;
  wire _0751_;
  wire _0752_;
  wire _0753_;
  wire _0754_;
  wire _0755_;
  wire _0756_;
  wire _0757_;
  wire _0758_;
  wire _0759_;
  wire _0760_;
  wire _0761_;
  wire _0762_;
  wire _0763_;
  wire _0764_;
  wire _0765_;
  wire _0766_;
  wire _0767_;
  wire _0768_;
  wire _0769_;
  wire _0770_;
  (* src = "expand_key_128.v:28|S4.v:26|S.v:11" *)
  wire [7:0] _0771_;
  wire _0772_;
  wire _0773_;
  wire _0774_;
  wire _0775_;
  wire _0776_;
  wire _0777_;
  wire _0778_;
  wire _0779_;
  wire _0780_;
  wire _0781_;
  wire _0782_;
  wire _0783_;
  wire _0784_;
  wire _0785_;
  wire _0786_;
  wire _0787_;
  wire _0788_;
  wire _0789_;
  wire _0790_;
  wire _0791_;
  wire _0792_;
  wire _0793_;
  wire _0794_;
  wire _0795_;
  wire _0796_;
  wire _0797_;
  wire _0798_;
  wire _0799_;
  wire _0800_;
  wire _0801_;
  wire _0802_;
  wire _0803_;
  wire _0804_;
  wire _0805_;
  wire _0806_;
  wire _0807_;
  wire _0808_;
  wire _0809_;
  wire _0810_;
  wire _0811_;
  wire _0812_;
  wire _0813_;
  wire _0814_;
  wire _0815_;
  wire _0816_;
  wire _0817_;
  wire _0818_;
  wire _0819_;
  wire _0820_;
  wire _0821_;
  wire _0822_;
  wire _0823_;
  wire _0824_;
  wire _0825_;
  wire _0826_;
  wire _0827_;
  wire _0828_;
  wire _0829_;
  wire _0830_;
  wire _0831_;
  wire _0832_;
  wire _0833_;
  wire _0834_;
  wire _0835_;
  wire _0836_;
  wire _0837_;
  wire _0838_;
  wire _0839_;
  wire _0840_;
  wire _0841_;
  wire _0842_;
  wire _0843_;
  wire _0844_;
  wire _0845_;
  wire _0846_;
  wire _0847_;
  wire _0848_;
  wire _0849_;
  wire _0850_;
  wire _0851_;
  wire _0852_;
  wire _0853_;
  wire _0854_;
  wire _0855_;
  wire _0856_;
  wire _0857_;
  wire _0858_;
  wire _0859_;
  wire _0860_;
  wire _0861_;
  wire _0862_;
  wire _0863_;
  wire _0864_;
  wire _0865_;
  wire _0866_;
  wire _0867_;
  wire _0868_;
  wire _0869_;
  wire _0870_;
  wire _0871_;
  wire _0872_;
  wire _0873_;
  wire _0874_;
  wire _0875_;
  wire _0876_;
  wire _0877_;
  wire _0878_;
  wire _0879_;
  wire _0880_;
  wire _0881_;
  wire _0882_;
  wire _0883_;
  wire _0884_;
  wire _0885_;
  wire _0886_;
  wire _0887_;
  wire _0888_;
  wire _0889_;
  wire _0890_;
  wire _0891_;
  wire _0892_;
  wire _0893_;
  wire _0894_;
  wire _0895_;
  wire _0896_;
  wire _0897_;
  wire _0898_;
  wire _0899_;
  wire _0900_;
  wire _0901_;
  wire _0902_;
  wire _0903_;
  wire _0904_;
  wire _0905_;
  wire _0906_;
  wire _0907_;
  wire _0908_;
  wire _0909_;
  wire _0910_;
  wire _0911_;
  wire _0912_;
  wire _0913_;
  wire _0914_;
  wire _0915_;
  wire _0916_;
  wire _0917_;
  wire _0918_;
  wire _0919_;
  wire _0920_;
  wire _0921_;
  wire _0922_;
  wire _0923_;
  wire _0924_;
  wire _0925_;
  wire _0926_;
  wire _0927_;
  wire _0928_;
  wire _0929_;
  wire _0930_;
  wire _0931_;
  wire _0932_;
  wire _0933_;
  wire _0934_;
  wire _0935_;
  wire _0936_;
  wire _0937_;
  wire _0938_;
  wire _0939_;
  wire _0940_;
  wire _0941_;
  wire _0942_;
  wire _0943_;
  wire _0944_;
  wire _0945_;
  wire _0946_;
  wire _0947_;
  wire _0948_;
  wire _0949_;
  wire _0950_;
  wire _0951_;
  wire _0952_;
  wire _0953_;
  wire _0954_;
  wire _0955_;
  wire _0956_;
  wire _0957_;
  wire _0958_;
  wire _0959_;
  wire _0960_;
  wire _0961_;
  wire _0962_;
  wire _0963_;
  wire _0964_;
  wire _0965_;
  wire _0966_;
  wire _0967_;
  wire _0968_;
  wire _0969_;
  wire _0970_;
  wire _0971_;
  wire _0972_;
  wire _0973_;
  wire _0974_;
  wire _0975_;
  wire _0976_;
  wire _0977_;
  wire _0978_;
  wire _0979_;
  wire _0980_;
  wire _0981_;
  wire _0982_;
  wire _0983_;
  wire _0984_;
  wire _0985_;
  wire _0986_;
  wire _0987_;
  wire _0988_;
  wire _0989_;
  wire _0990_;
  wire _0991_;
  wire _0992_;
  wire _0993_;
  wire _0994_;
  wire _0995_;
  wire _0996_;
  wire _0997_;
  wire _0998_;
  wire _0999_;
  wire _1000_;
  wire _1001_;
  wire _1002_;
  wire _1003_;
  wire _1004_;
  wire _1005_;
  wire _1006_;
  wire _1007_;
  wire _1008_;
  wire _1009_;
  wire _1010_;
  wire _1011_;
  wire _1012_;
  wire _1013_;
  wire _1014_;
  wire _1015_;
  wire _1016_;
  wire _1017_;
  wire _1018_;
  wire _1019_;
  wire _1020_;
  wire _1021_;
  wire _1022_;
  wire _1023_;
  wire _1024_;
  wire _1025_;
  wire _1026_;
  wire _1027_;
  (* src = "expand_key_128.v:28|S4.v:26|S.v:5" *)
  wire \S4_0.S_0.clk ;
  (* src = "expand_key_128.v:28|S4.v:26|S.v:6" *)
  wire [7:0] \S4_0.S_0.in ;
  (* src = "expand_key_128.v:28|S4.v:26|S.v:7" *)
  reg [7:0] \S4_0.S_0.out ;
  (* src = "expand_key_128.v:28|S4.v:26|S.v:5" *)
  wire \S4_0.S_1.clk ;
  (* src = "expand_key_128.v:28|S4.v:26|S.v:6" *)
  wire [7:0] \S4_0.S_1.in ;
  (* src = "expand_key_128.v:28|S4.v:26|S.v:7" *)
  reg [7:0] \S4_0.S_1.out ;
  (* src = "expand_key_128.v:28|S4.v:26|S.v:5" *)
  wire \S4_0.S_2.clk ;
  (* src = "expand_key_128.v:28|S4.v:26|S.v:6" *)
  wire [7:0] \S4_0.S_2.in ;
  (* src = "expand_key_128.v:28|S4.v:26|S.v:7" *)
  reg [7:0] \S4_0.S_2.out ;
  (* src = "expand_key_128.v:28|S4.v:26|S.v:5" *)
  wire \S4_0.S_3.clk ;
  (* src = "expand_key_128.v:28|S4.v:26|S.v:6" *)
  wire [7:0] \S4_0.S_3.in ;
  (* src = "expand_key_128.v:28|S4.v:26|S.v:7" *)
  reg [7:0] \S4_0.S_3.out ;
  (* src = "expand_key_128.v:28|S4.v:22" *)
  wire \S4_0.clk ;
  (* src = "expand_key_128.v:28|S4.v:23" *)
  wire [31:0] \S4_0.in ;
  (* src = "expand_key_128.v:28|S4.v:24" *)
  wire [31:0] \S4_0.out ;
  (* src = "expand_key_128.v:6" *)
  input clk;
  (* src = "expand_key_128.v:7" *)
  input [127:0] in;
  (* src = "expand_key_128.v:12" *)
  wire [31:0] k0;
  (* src = "expand_key_128.v:15" *)
  reg [31:0] k0a;
  (* src = "expand_key_128.v:16" *)
  wire [31:0] k0b;
  (* src = "expand_key_128.v:12" *)
  wire [31:0] k1;
  (* src = "expand_key_128.v:15" *)
  reg [31:0] k1a;
  (* src = "expand_key_128.v:16" *)
  wire [31:0] k1b;
  (* src = "expand_key_128.v:12" *)
  wire [31:0] k2;
  (* src = "expand_key_128.v:15" *)
  reg [31:0] k2a;
  (* src = "expand_key_128.v:16" *)
  wire [31:0] k2b;
  (* src = "expand_key_128.v:12" *)
  wire [31:0] k3;
  (* src = "expand_key_128.v:15" *)
  reg [31:0] k3a;
  (* src = "expand_key_128.v:16" *)
  wire [31:0] k3b;
  (* src = "expand_key_128.v:16" *)
  wire [31:0] k4a;
  (* src = "expand_key_128.v:9" *)
  output [127:0] out_1;
  reg [127:0] out_1;
  (* src = "expand_key_128.v:10" *)
  output [127:0] out_2;
  (* src = "expand_key_128.v:8" *)
  input [7:0] rcon;
  (* src = "expand_key_128.v:12" *)
  wire [31:0] v0;
  (* src = "expand_key_128.v:12" *)
  wire [31:0] v1;
  (* src = "expand_key_128.v:12" *)
  wire [31:0] v2;
  (* src = "expand_key_128.v:12" *)
  wire [31:0] v3;
  always @(posedge clk)
      out_1 <= { k0b, k1b, k2b, k3b };
  always @(posedge clk)
      k0a <= { v0[31:24], in[119:96] };
  always @(posedge clk)
      k1a <= v1;
  always @(posedge clk)
      k2a <= v2;
  always @(posedge clk)
      k3a <= v3;
  always @(posedge clk)
      \S4_0.S_0.out  <= _0000_;
  assign _0001_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'ha8;
  assign _0002_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'ha7;
  assign _0003_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'ha6;
  assign _0004_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'ha5;
  assign _0005_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'ha4;
  assign _0006_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'ha3;
  assign _0007_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'ha2;
  assign _0008_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'ha1;
  assign _0009_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'ha0;
  assign _0010_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'h9f;
  assign _0011_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'h9e;
  assign _0012_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'h9d;
  assign _0013_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'h9c;
  assign _0014_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'h9b;
  assign _0015_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'h9a;
  assign _0016_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'h99;
  assign _0017_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'h98;
  assign _0018_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'h97;
  assign _0019_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'h96;
  assign _0020_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'h95;
  function [7:0] _1054_;
    input [7:0] a;
    input [2047:0] b;
    input [255:0] s;
    (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *)
    (* parallel_case *)
    casez (s)
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1:
        _1054_ = b[7:0];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?:
        _1054_ = b[15:8];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??:
        _1054_ = b[23:16];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???:
        _1054_ = b[31:24];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????:
        _1054_ = b[39:32];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????:
        _1054_ = b[47:40];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????:
        _1054_ = b[55:48];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????:
        _1054_ = b[63:56];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????:
        _1054_ = b[71:64];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????:
        _1054_ = b[79:72];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????:
        _1054_ = b[87:80];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????:
        _1054_ = b[95:88];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????:
        _1054_ = b[103:96];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????:
        _1054_ = b[111:104];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????:
        _1054_ = b[119:112];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????:
        _1054_ = b[127:120];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????:
        _1054_ = b[135:128];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????:
        _1054_ = b[143:136];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????:
        _1054_ = b[151:144];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????:
        _1054_ = b[159:152];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????:
        _1054_ = b[167:160];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????:
        _1054_ = b[175:168];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????:
        _1054_ = b[183:176];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????:
        _1054_ = b[191:184];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????:
        _1054_ = b[199:192];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????:
        _1054_ = b[207:200];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????:
        _1054_ = b[215:208];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????:
        _1054_ = b[223:216];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????:
        _1054_ = b[231:224];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????:
        _1054_ = b[239:232];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????:
        _1054_ = b[247:240];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????:
        _1054_ = b[255:248];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????:
        _1054_ = b[263:256];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????:
        _1054_ = b[271:264];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????:
        _1054_ = b[279:272];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????:
        _1054_ = b[287:280];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????:
        _1054_ = b[295:288];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????:
        _1054_ = b[303:296];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????:
        _1054_ = b[311:304];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????:
        _1054_ = b[319:312];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????:
        _1054_ = b[327:320];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????:
        _1054_ = b[335:328];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????:
        _1054_ = b[343:336];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????:
        _1054_ = b[351:344];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????:
        _1054_ = b[359:352];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????:
        _1054_ = b[367:360];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????:
        _1054_ = b[375:368];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????:
        _1054_ = b[383:376];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????:
        _1054_ = b[391:384];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????:
        _1054_ = b[399:392];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????:
        _1054_ = b[407:400];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????:
        _1054_ = b[415:408];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????:
        _1054_ = b[423:416];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????:
        _1054_ = b[431:424];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????:
        _1054_ = b[439:432];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????:
        _1054_ = b[447:440];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????:
        _1054_ = b[455:448];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????:
        _1054_ = b[463:456];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????:
        _1054_ = b[471:464];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????:
        _1054_ = b[479:472];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????:
        _1054_ = b[487:480];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????:
        _1054_ = b[495:488];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????:
        _1054_ = b[503:496];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????:
        _1054_ = b[511:504];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????:
        _1054_ = b[519:512];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????:
        _1054_ = b[527:520];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????:
        _1054_ = b[535:528];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????:
        _1054_ = b[543:536];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????:
        _1054_ = b[551:544];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????:
        _1054_ = b[559:552];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????:
        _1054_ = b[567:560];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????:
        _1054_ = b[575:568];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????:
        _1054_ = b[583:576];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????:
        _1054_ = b[591:584];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????:
        _1054_ = b[599:592];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????:
        _1054_ = b[607:600];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????:
        _1054_ = b[615:608];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????:
        _1054_ = b[623:616];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????:
        _1054_ = b[631:624];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????:
        _1054_ = b[639:632];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????:
        _1054_ = b[647:640];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????:
        _1054_ = b[655:648];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????:
        _1054_ = b[663:656];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????:
        _1054_ = b[671:664];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????:
        _1054_ = b[679:672];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????:
        _1054_ = b[687:680];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????:
        _1054_ = b[695:688];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????:
        _1054_ = b[703:696];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????:
        _1054_ = b[711:704];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????:
        _1054_ = b[719:712];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????:
        _1054_ = b[727:720];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????:
        _1054_ = b[735:728];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????:
        _1054_ = b[743:736];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????:
        _1054_ = b[751:744];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????:
        _1054_ = b[759:752];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????:
        _1054_ = b[767:760];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????:
        _1054_ = b[775:768];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????:
        _1054_ = b[783:776];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????:
        _1054_ = b[791:784];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????:
        _1054_ = b[799:792];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1054_ = b[807:800];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1054_ = b[815:808];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1054_ = b[823:816];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1054_ = b[831:824];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1054_ = b[839:832];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1054_ = b[847:840];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1054_ = b[855:848];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1054_ = b[863:856];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1054_ = b[871:864];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1054_ = b[879:872];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1054_ = b[887:880];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1054_ = b[895:888];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1054_ = b[903:896];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1054_ = b[911:904];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1054_ = b[919:912];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1054_ = b[927:920];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1054_ = b[935:928];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1054_ = b[943:936];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1054_ = b[951:944];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1054_ = b[959:952];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1054_ = b[967:960];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1054_ = b[975:968];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1054_ = b[983:976];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1054_ = b[991:984];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1054_ = b[999:992];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1054_ = b[1007:1000];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1054_ = b[1015:1008];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1054_ = b[1023:1016];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1054_ = b[1031:1024];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1054_ = b[1039:1032];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1054_ = b[1047:1040];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1054_ = b[1055:1048];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1054_ = b[1063:1056];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1054_ = b[1071:1064];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1054_ = b[1079:1072];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1054_ = b[1087:1080];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1054_ = b[1095:1088];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1054_ = b[1103:1096];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1054_ = b[1111:1104];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1054_ = b[1119:1112];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1054_ = b[1127:1120];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1054_ = b[1135:1128];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1054_ = b[1143:1136];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1054_ = b[1151:1144];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1054_ = b[1159:1152];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1054_ = b[1167:1160];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1054_ = b[1175:1168];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1054_ = b[1183:1176];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1054_ = b[1191:1184];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1054_ = b[1199:1192];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1054_ = b[1207:1200];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1054_ = b[1215:1208];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1054_ = b[1223:1216];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1054_ = b[1231:1224];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1054_ = b[1239:1232];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1054_ = b[1247:1240];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1054_ = b[1255:1248];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1054_ = b[1263:1256];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1054_ = b[1271:1264];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1054_ = b[1279:1272];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1054_ = b[1287:1280];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1054_ = b[1295:1288];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1054_ = b[1303:1296];
      256'b????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1054_ = b[1311:1304];
      256'b???????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1054_ = b[1319:1312];
      256'b??????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1054_ = b[1327:1320];
      256'b?????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1054_ = b[1335:1328];
      256'b????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1054_ = b[1343:1336];
      256'b???????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1054_ = b[1351:1344];
      256'b??????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1054_ = b[1359:1352];
      256'b?????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1054_ = b[1367:1360];
      256'b????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1054_ = b[1375:1368];
      256'b???????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1054_ = b[1383:1376];
      256'b??????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1054_ = b[1391:1384];
      256'b?????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1054_ = b[1399:1392];
      256'b????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1054_ = b[1407:1400];
      256'b???????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1054_ = b[1415:1408];
      256'b??????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1054_ = b[1423:1416];
      256'b?????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1054_ = b[1431:1424];
      256'b????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1054_ = b[1439:1432];
      256'b???????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1054_ = b[1447:1440];
      256'b??????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1054_ = b[1455:1448];
      256'b?????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1054_ = b[1463:1456];
      256'b????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1054_ = b[1471:1464];
      256'b???????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1054_ = b[1479:1472];
      256'b??????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1054_ = b[1487:1480];
      256'b?????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1054_ = b[1495:1488];
      256'b????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1054_ = b[1503:1496];
      256'b???????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1054_ = b[1511:1504];
      256'b??????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1054_ = b[1519:1512];
      256'b?????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1054_ = b[1527:1520];
      256'b????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1054_ = b[1535:1528];
      256'b???????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1054_ = b[1543:1536];
      256'b??????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1054_ = b[1551:1544];
      256'b?????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1054_ = b[1559:1552];
      256'b????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1054_ = b[1567:1560];
      256'b???????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1054_ = b[1575:1568];
      256'b??????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1054_ = b[1583:1576];
      256'b?????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1054_ = b[1591:1584];
      256'b????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1054_ = b[1599:1592];
      256'b???????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1054_ = b[1607:1600];
      256'b??????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1054_ = b[1615:1608];
      256'b?????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1054_ = b[1623:1616];
      256'b????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1054_ = b[1631:1624];
      256'b???????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1054_ = b[1639:1632];
      256'b??????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1054_ = b[1647:1640];
      256'b?????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1054_ = b[1655:1648];
      256'b????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1054_ = b[1663:1656];
      256'b???????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1054_ = b[1671:1664];
      256'b??????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1054_ = b[1679:1672];
      256'b?????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1054_ = b[1687:1680];
      256'b????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1054_ = b[1695:1688];
      256'b???????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1054_ = b[1703:1696];
      256'b??????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1054_ = b[1711:1704];
      256'b?????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1054_ = b[1719:1712];
      256'b????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1054_ = b[1727:1720];
      256'b???????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1054_ = b[1735:1728];
      256'b??????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1054_ = b[1743:1736];
      256'b?????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1054_ = b[1751:1744];
      256'b????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1054_ = b[1759:1752];
      256'b???????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1054_ = b[1767:1760];
      256'b??????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1054_ = b[1775:1768];
      256'b?????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1054_ = b[1783:1776];
      256'b????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1054_ = b[1791:1784];
      256'b???????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1054_ = b[1799:1792];
      256'b??????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1054_ = b[1807:1800];
      256'b?????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1054_ = b[1815:1808];
      256'b????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1054_ = b[1823:1816];
      256'b???????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1054_ = b[1831:1824];
      256'b??????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1054_ = b[1839:1832];
      256'b?????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1054_ = b[1847:1840];
      256'b????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1054_ = b[1855:1848];
      256'b???????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1054_ = b[1863:1856];
      256'b??????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1054_ = b[1871:1864];
      256'b?????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1054_ = b[1879:1872];
      256'b????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1054_ = b[1887:1880];
      256'b???????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1054_ = b[1895:1888];
      256'b??????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1054_ = b[1903:1896];
      256'b?????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1054_ = b[1911:1904];
      256'b????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1054_ = b[1919:1912];
      256'b???????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1054_ = b[1927:1920];
      256'b??????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1054_ = b[1935:1928];
      256'b?????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1054_ = b[1943:1936];
      256'b????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1054_ = b[1951:1944];
      256'b???????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1054_ = b[1959:1952];
      256'b??????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1054_ = b[1967:1960];
      256'b?????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1054_ = b[1975:1968];
      256'b????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1054_ = b[1983:1976];
      256'b???????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1054_ = b[1991:1984];
      256'b??????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1054_ = b[1999:1992];
      256'b?????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1054_ = b[2007:2000];
      256'b????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1054_ = b[2015:2008];
      256'b???1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1054_ = b[2023:2016];
      256'b??1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1054_ = b[2031:2024];
      256'b?1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1054_ = b[2039:2032];
      256'b1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1054_ = b[2047:2040];
      default:
        _1054_ = a;
    endcase
  endfunction
  assign _0000_ = _1054_(\S4_0.S_0.out , 2048'h637c777bf26b6fc53001672bfed7ab76ca82c97dfa5947f0add4a2af9ca472c0b7fd9326363ff7cc34a5e5f171d8311504c723c31896059a071280e2eb27b27509832c1a1b6e5aa0523bd6b329e32f8453d100ed20fcb15b6acbbe394a4c58cfd0efaafb434d338545f9027f503c9fa851a3408f929d38f5bcb6da2110fff3d2cd0c13ec5f974417c4a77e3d645d197360814fdc222a908846eeb814de5e0bdbe0323a0a4906245cc2d3ac629195e479e7c8376d8dd54ea96c56f4ea657aae08ba78252e1ca6b4c6e8dd741f4bbd8b8a703eb5664803f60e613557b986c11d9ee1f8981169d98e949b1e87e9ce5528df8ca1890dbfe6426841992d0fb054bb16, { _0182_, _0181_, _0180_, _0179_, _0178_, _0177_, _0176_, _0175_, _0174_, _0172_, _0171_, _0170_, _0169_, _0168_, _0167_, _0166_, _0165_, _0164_, _0163_, _0161_, _0160_, _0159_, _0158_, _0157_, _0156_, _0155_, _0154_, _0153_, _0152_, _0150_, _0149_, _0148_, _0147_, _0146_, _0145_, _0144_, _0143_, _0142_, _0141_, _0139_, _0138_, _0137_, _0136_, _0135_, _0134_, _0133_, _0132_, _0131_, _0130_, _0128_, _0127_, _0126_, _0125_, _0124_, _0123_, _0122_, _0121_, _0120_, _0119_, _0117_, _0116_, _0115_, _0114_, _0113_, _0112_, _0111_, _0110_, _0109_, _0108_, _0106_, _0105_, _0104_, _0103_, _0102_, _0101_, _0100_, _0099_, _0098_, _0097_, _0095_, _0094_, _0093_, _0092_, _0091_, _0090_, _0089_, _0088_, _0087_, _0086_, _0084_, _0083_, _0082_, _0081_, _0080_, _0079_, _0078_, _0077_, _0076_, _0075_, _0073_, _0072_, _0071_, _0070_, _0069_, _0068_, _0067_, _0066_, _0065_, _0064_, _0062_, _0061_, _0060_, _0059_, _0058_, _0057_, _0056_, _0055_, _0054_, _0053_, _0051_, _0050_, _0049_, _0048_, _0047_, _0046_, _0045_, _0044_, _0043_, _0042_, _0040_, _0039_, _0038_, _0037_, _0036_, _0035_, _0034_, _0033_, _0032_, _0031_, _0030_, _0029_, _0028_, _0027_, _0026_, _0025_, _0024_, _0023_, _0022_, _0021_, _0020_, _0019_, _0018_, _0017_, _0016_, _0015_, _0014_, _0013_, _0012_, _0011_, _0010_, _0009_, _0008_, _0007_, _0006_, _0005_, _0004_, _0003_, _0002_, _0001_, _0256_, _0255_, _0254_, _0253_, _0252_, _0251_, _0250_, _0249_, _0248_, _0247_, _0246_, _0245_, _0244_, _0243_, _0242_, _0241_, _0240_, _0239_, _0238_, _0237_, _0236_, _0235_, _0234_, _0233_, _0232_, _0231_, _0230_, _0229_, _0228_, _0227_, _0226_, _0225_, _0224_, _0223_, _0222_, _0221_, _0220_, _0219_, _0218_, _0217_, _0216_, _0215_, _0214_, _0213_, _0212_, _0211_, _0210_, _0209_, _0208_, _0207_, _0206_, _0205_, _0204_, _0203_, _0202_, _0201_, _0200_, _0199_, _0198_, _0197_, _0196_, _0195_, _0194_, _0193_, _0192_, _0191_, _0190_, _0189_, _0188_, _0187_, _0186_, _0185_, _0184_, _0183_, _0173_, _0162_, _0151_, _0140_, _0129_, _0118_, _0107_, _0096_, _0085_, _0074_, _0063_, _0052_, _0041_ });
  assign _0021_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'h94;
  assign _0022_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'h93;
  assign _0023_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'h92;
  assign _0024_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'h91;
  assign _0025_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'h90;
  assign _0026_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'h8f;
  assign _0027_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'h8e;
  assign _0028_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'h8d;
  assign _0029_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'h8c;
  assign _0030_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'h8b;
  assign _0031_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'h8a;
  assign _0032_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'h89;
  assign _0033_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'h88;
  assign _0034_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'h87;
  assign _0035_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'h86;
  assign _0036_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'h85;
  assign _0037_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'h84;
  assign _0038_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'h83;
  assign _0039_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'h82;
  assign _0040_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'h81;
  assign _0041_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hff;
  assign _0042_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'h80;
  assign _0043_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h7f;
  assign _0044_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h7e;
  assign _0045_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h7d;
  assign _0046_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h7c;
  assign _0047_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h7b;
  assign _0048_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h7a;
  assign _0049_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h79;
  assign _0050_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h78;
  assign _0051_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h77;
  assign _0052_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hfe;
  assign _0053_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h76;
  assign _0054_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h75;
  assign _0055_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h74;
  assign _0056_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h73;
  assign _0057_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h72;
  assign _0058_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h71;
  assign _0059_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h70;
  assign _0060_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h6f;
  assign _0061_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h6e;
  assign _0062_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h6d;
  assign _0063_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hfd;
  assign _0064_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h6c;
  assign _0065_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h6b;
  assign _0066_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h6a;
  assign _0067_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h69;
  assign _0068_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h68;
  assign _0069_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h67;
  assign _0070_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h66;
  assign _0071_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h65;
  assign _0072_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h64;
  assign _0073_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h63;
  assign _0074_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hfc;
  assign _0075_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h62;
  assign _0076_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h61;
  assign _0077_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h60;
  assign _0078_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h5f;
  assign _0079_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h5e;
  assign _0080_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h5d;
  assign _0081_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h5c;
  assign _0082_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h5b;
  assign _0083_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h5a;
  assign _0084_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h59;
  assign _0085_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hfb;
  assign _0086_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h58;
  assign _0087_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h57;
  assign _0088_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h56;
  assign _0089_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h55;
  assign _0090_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h54;
  assign _0091_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h53;
  assign _0092_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h52;
  assign _0093_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h51;
  assign _0094_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h50;
  assign _0095_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h4f;
  assign _0096_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hfa;
  assign _0097_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h4e;
  assign _0098_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h4d;
  assign _0099_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h4c;
  assign _0100_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h4b;
  assign _0101_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h4a;
  assign _0102_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h49;
  assign _0103_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h48;
  assign _0104_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h47;
  assign _0105_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h46;
  assign _0106_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h45;
  assign _0107_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hf9;
  assign _0108_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h44;
  assign _0109_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h43;
  assign _0110_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h42;
  assign _0111_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h41;
  assign _0112_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h40;
  assign _0113_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 6'h3f;
  assign _0114_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 6'h3e;
  assign _0115_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 6'h3d;
  assign _0116_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 6'h3c;
  assign _0117_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 6'h3b;
  assign _0118_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hf8;
  assign _0119_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 6'h3a;
  assign _0120_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 6'h39;
  assign _0121_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 6'h38;
  assign _0122_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 6'h37;
  assign _0123_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 6'h36;
  assign _0124_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 6'h35;
  assign _0125_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 6'h34;
  assign _0126_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 6'h33;
  assign _0127_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 6'h32;
  assign _0128_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 6'h31;
  assign _0129_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hf7;
  assign _0130_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 6'h30;
  assign _0131_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 6'h2f;
  assign _0132_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 6'h2e;
  assign _0133_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 6'h2d;
  assign _0134_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 6'h2c;
  assign _0135_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 6'h2b;
  assign _0136_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 6'h2a;
  assign _0137_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 6'h29;
  assign _0138_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 6'h28;
  assign _0139_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 6'h27;
  assign _0140_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hf6;
  assign _0141_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 6'h26;
  assign _0142_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 6'h25;
  assign _0143_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 6'h24;
  assign _0144_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 6'h23;
  assign _0145_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 6'h22;
  assign _0146_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 6'h21;
  assign _0147_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 6'h20;
  assign _0148_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 5'h1f;
  assign _0149_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 5'h1e;
  assign _0150_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 5'h1d;
  assign _0151_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hf5;
  assign _0152_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 5'h1c;
  assign _0153_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 5'h1b;
  assign _0154_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 5'h1a;
  assign _0155_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 5'h19;
  assign _0156_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 5'h18;
  assign _0157_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 5'h17;
  assign _0158_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 5'h16;
  assign _0159_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 5'h15;
  assign _0160_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 5'h14;
  assign _0161_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 5'h13;
  assign _0162_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hf4;
  assign _0163_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 5'h12;
  assign _0164_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 5'h11;
  assign _0165_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 5'h10;
  assign _0166_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 4'hf;
  assign _0167_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 4'he;
  assign _0168_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 4'hd;
  assign _0169_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 4'hc;
  assign _0170_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 4'hb;
  assign _0171_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 4'ha;
  assign _0172_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 4'h9;
  assign _0173_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hf3;
  assign _0174_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 4'h8;
  assign _0175_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 3'h7;
  assign _0176_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 3'h6;
  assign _0177_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 3'h5;
  assign _0178_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 3'h4;
  assign _0179_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 2'h3;
  assign _0180_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 2'h2;
  assign _0181_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 1'h1;
  assign _0182_ = ! (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) in[23:16];
  assign _0183_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hf2;
  assign _0184_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hf1;
  assign _0185_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hf0;
  assign _0186_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hef;
  assign _0187_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hee;
  assign _0188_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hed;
  assign _0189_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hec;
  assign _0190_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'heb;
  assign _0191_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hea;
  assign _0192_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'he9;
  assign _0193_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'he8;
  assign _0194_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'he7;
  assign _0195_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'he6;
  assign _0196_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'he5;
  assign _0197_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'he4;
  assign _0198_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'he3;
  assign _0199_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'he2;
  assign _0200_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'he1;
  assign _0201_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'he0;
  assign _0202_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hdf;
  assign _0203_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hde;
  assign _0204_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hdd;
  assign _0205_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hdc;
  assign _0206_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hdb;
  assign _0207_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hda;
  assign _0208_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hd9;
  assign _0209_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hd8;
  assign _0210_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hd7;
  assign _0211_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hd6;
  assign _0212_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hd5;
  assign _0213_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hd4;
  assign _0214_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hd3;
  assign _0215_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hd2;
  assign _0216_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hd1;
  assign _0217_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hd0;
  assign _0218_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hcf;
  assign _0219_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hce;
  assign _0220_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hcd;
  assign _0221_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hcc;
  assign _0222_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hcb;
  assign _0223_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hca;
  assign _0224_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hc9;
  assign _0225_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hc8;
  assign _0226_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hc7;
  assign _0227_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hc6;
  assign _0228_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hc5;
  assign _0229_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hc4;
  assign _0230_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hc3;
  assign _0231_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hc2;
  assign _0232_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hc1;
  assign _0233_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hc0;
  assign _0234_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hbf;
  assign _0235_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hbe;
  assign _0236_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hbd;
  assign _0237_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hbc;
  assign _0238_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hbb;
  assign _0239_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hba;
  assign _0240_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hb9;
  assign _0241_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hb8;
  assign _0242_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hb7;
  assign _0243_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hb6;
  assign _0244_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hb5;
  assign _0245_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hb4;
  assign _0246_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hb3;
  assign _0247_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hb2;
  assign _0248_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hb1;
  assign _0249_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hb0;
  assign _0250_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'haf;
  assign _0251_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hae;
  assign _0252_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'had;
  assign _0253_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hac;
  assign _0254_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hab;
  assign _0255_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'haa;
  assign _0256_ = in[23:16] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'ha9;
  always @(posedge clk)
      \S4_0.S_1.out  <= _0257_;
  assign _0258_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'ha8;
  assign _0259_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'ha7;
  assign _0260_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'ha6;
  assign _0261_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'ha5;
  assign _0262_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'ha4;
  assign _0263_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'ha3;
  assign _0264_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'ha2;
  assign _0265_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'ha1;
  assign _0266_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'ha0;
  assign _0267_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'h9f;
  assign _0268_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'h9e;
  assign _0269_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'h9d;
  assign _0270_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'h9c;
  assign _0271_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'h9b;
  assign _0272_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'h9a;
  assign _0273_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'h99;
  assign _0274_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'h98;
  assign _0275_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'h97;
  assign _0276_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'h96;
  assign _0277_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'h95;
  function [7:0] _1312_;
    input [7:0] a;
    input [2047:0] b;
    input [255:0] s;
    (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *)
    (* parallel_case *)
    casez (s)
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1:
        _1312_ = b[7:0];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?:
        _1312_ = b[15:8];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??:
        _1312_ = b[23:16];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???:
        _1312_ = b[31:24];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????:
        _1312_ = b[39:32];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????:
        _1312_ = b[47:40];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????:
        _1312_ = b[55:48];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????:
        _1312_ = b[63:56];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????:
        _1312_ = b[71:64];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????:
        _1312_ = b[79:72];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????:
        _1312_ = b[87:80];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????:
        _1312_ = b[95:88];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????:
        _1312_ = b[103:96];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????:
        _1312_ = b[111:104];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????:
        _1312_ = b[119:112];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????:
        _1312_ = b[127:120];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????:
        _1312_ = b[135:128];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????:
        _1312_ = b[143:136];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????:
        _1312_ = b[151:144];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????:
        _1312_ = b[159:152];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????:
        _1312_ = b[167:160];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????:
        _1312_ = b[175:168];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????:
        _1312_ = b[183:176];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????:
        _1312_ = b[191:184];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????:
        _1312_ = b[199:192];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????:
        _1312_ = b[207:200];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????:
        _1312_ = b[215:208];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????:
        _1312_ = b[223:216];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????:
        _1312_ = b[231:224];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????:
        _1312_ = b[239:232];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????:
        _1312_ = b[247:240];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????:
        _1312_ = b[255:248];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????:
        _1312_ = b[263:256];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????:
        _1312_ = b[271:264];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????:
        _1312_ = b[279:272];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????:
        _1312_ = b[287:280];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????:
        _1312_ = b[295:288];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????:
        _1312_ = b[303:296];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????:
        _1312_ = b[311:304];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????:
        _1312_ = b[319:312];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????:
        _1312_ = b[327:320];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????:
        _1312_ = b[335:328];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????:
        _1312_ = b[343:336];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????:
        _1312_ = b[351:344];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????:
        _1312_ = b[359:352];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????:
        _1312_ = b[367:360];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????:
        _1312_ = b[375:368];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????:
        _1312_ = b[383:376];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????:
        _1312_ = b[391:384];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????:
        _1312_ = b[399:392];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????:
        _1312_ = b[407:400];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????:
        _1312_ = b[415:408];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????:
        _1312_ = b[423:416];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????:
        _1312_ = b[431:424];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????:
        _1312_ = b[439:432];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????:
        _1312_ = b[447:440];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????:
        _1312_ = b[455:448];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????:
        _1312_ = b[463:456];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????:
        _1312_ = b[471:464];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????:
        _1312_ = b[479:472];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????:
        _1312_ = b[487:480];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????:
        _1312_ = b[495:488];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????:
        _1312_ = b[503:496];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????:
        _1312_ = b[511:504];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????:
        _1312_ = b[519:512];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????:
        _1312_ = b[527:520];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????:
        _1312_ = b[535:528];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????:
        _1312_ = b[543:536];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????:
        _1312_ = b[551:544];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????:
        _1312_ = b[559:552];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????:
        _1312_ = b[567:560];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????:
        _1312_ = b[575:568];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????:
        _1312_ = b[583:576];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????:
        _1312_ = b[591:584];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????:
        _1312_ = b[599:592];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????:
        _1312_ = b[607:600];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????:
        _1312_ = b[615:608];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????:
        _1312_ = b[623:616];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????:
        _1312_ = b[631:624];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????:
        _1312_ = b[639:632];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????:
        _1312_ = b[647:640];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????:
        _1312_ = b[655:648];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????:
        _1312_ = b[663:656];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????:
        _1312_ = b[671:664];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????:
        _1312_ = b[679:672];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????:
        _1312_ = b[687:680];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????:
        _1312_ = b[695:688];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????:
        _1312_ = b[703:696];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????:
        _1312_ = b[711:704];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????:
        _1312_ = b[719:712];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????:
        _1312_ = b[727:720];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????:
        _1312_ = b[735:728];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????:
        _1312_ = b[743:736];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????:
        _1312_ = b[751:744];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????:
        _1312_ = b[759:752];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????:
        _1312_ = b[767:760];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????:
        _1312_ = b[775:768];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????:
        _1312_ = b[783:776];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????:
        _1312_ = b[791:784];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????:
        _1312_ = b[799:792];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1312_ = b[807:800];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1312_ = b[815:808];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1312_ = b[823:816];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1312_ = b[831:824];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1312_ = b[839:832];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1312_ = b[847:840];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1312_ = b[855:848];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1312_ = b[863:856];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1312_ = b[871:864];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1312_ = b[879:872];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1312_ = b[887:880];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1312_ = b[895:888];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1312_ = b[903:896];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1312_ = b[911:904];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1312_ = b[919:912];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1312_ = b[927:920];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1312_ = b[935:928];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1312_ = b[943:936];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1312_ = b[951:944];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1312_ = b[959:952];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1312_ = b[967:960];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1312_ = b[975:968];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1312_ = b[983:976];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1312_ = b[991:984];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1312_ = b[999:992];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1312_ = b[1007:1000];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1312_ = b[1015:1008];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1312_ = b[1023:1016];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1312_ = b[1031:1024];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1312_ = b[1039:1032];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1312_ = b[1047:1040];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1312_ = b[1055:1048];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1312_ = b[1063:1056];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1312_ = b[1071:1064];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1312_ = b[1079:1072];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1312_ = b[1087:1080];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1312_ = b[1095:1088];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1312_ = b[1103:1096];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1312_ = b[1111:1104];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1312_ = b[1119:1112];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1312_ = b[1127:1120];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1312_ = b[1135:1128];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1312_ = b[1143:1136];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1312_ = b[1151:1144];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1312_ = b[1159:1152];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1312_ = b[1167:1160];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1312_ = b[1175:1168];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1312_ = b[1183:1176];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1312_ = b[1191:1184];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1312_ = b[1199:1192];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1312_ = b[1207:1200];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1312_ = b[1215:1208];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1312_ = b[1223:1216];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1312_ = b[1231:1224];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1312_ = b[1239:1232];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1312_ = b[1247:1240];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1312_ = b[1255:1248];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1312_ = b[1263:1256];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1312_ = b[1271:1264];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1312_ = b[1279:1272];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1312_ = b[1287:1280];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1312_ = b[1295:1288];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1312_ = b[1303:1296];
      256'b????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1312_ = b[1311:1304];
      256'b???????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1312_ = b[1319:1312];
      256'b??????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1312_ = b[1327:1320];
      256'b?????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1312_ = b[1335:1328];
      256'b????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1312_ = b[1343:1336];
      256'b???????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1312_ = b[1351:1344];
      256'b??????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1312_ = b[1359:1352];
      256'b?????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1312_ = b[1367:1360];
      256'b????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1312_ = b[1375:1368];
      256'b???????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1312_ = b[1383:1376];
      256'b??????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1312_ = b[1391:1384];
      256'b?????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1312_ = b[1399:1392];
      256'b????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1312_ = b[1407:1400];
      256'b???????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1312_ = b[1415:1408];
      256'b??????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1312_ = b[1423:1416];
      256'b?????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1312_ = b[1431:1424];
      256'b????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1312_ = b[1439:1432];
      256'b???????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1312_ = b[1447:1440];
      256'b??????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1312_ = b[1455:1448];
      256'b?????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1312_ = b[1463:1456];
      256'b????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1312_ = b[1471:1464];
      256'b???????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1312_ = b[1479:1472];
      256'b??????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1312_ = b[1487:1480];
      256'b?????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1312_ = b[1495:1488];
      256'b????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1312_ = b[1503:1496];
      256'b???????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1312_ = b[1511:1504];
      256'b??????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1312_ = b[1519:1512];
      256'b?????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1312_ = b[1527:1520];
      256'b????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1312_ = b[1535:1528];
      256'b???????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1312_ = b[1543:1536];
      256'b??????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1312_ = b[1551:1544];
      256'b?????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1312_ = b[1559:1552];
      256'b????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1312_ = b[1567:1560];
      256'b???????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1312_ = b[1575:1568];
      256'b??????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1312_ = b[1583:1576];
      256'b?????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1312_ = b[1591:1584];
      256'b????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1312_ = b[1599:1592];
      256'b???????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1312_ = b[1607:1600];
      256'b??????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1312_ = b[1615:1608];
      256'b?????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1312_ = b[1623:1616];
      256'b????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1312_ = b[1631:1624];
      256'b???????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1312_ = b[1639:1632];
      256'b??????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1312_ = b[1647:1640];
      256'b?????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1312_ = b[1655:1648];
      256'b????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1312_ = b[1663:1656];
      256'b???????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1312_ = b[1671:1664];
      256'b??????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1312_ = b[1679:1672];
      256'b?????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1312_ = b[1687:1680];
      256'b????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1312_ = b[1695:1688];
      256'b???????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1312_ = b[1703:1696];
      256'b??????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1312_ = b[1711:1704];
      256'b?????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1312_ = b[1719:1712];
      256'b????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1312_ = b[1727:1720];
      256'b???????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1312_ = b[1735:1728];
      256'b??????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1312_ = b[1743:1736];
      256'b?????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1312_ = b[1751:1744];
      256'b????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1312_ = b[1759:1752];
      256'b???????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1312_ = b[1767:1760];
      256'b??????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1312_ = b[1775:1768];
      256'b?????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1312_ = b[1783:1776];
      256'b????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1312_ = b[1791:1784];
      256'b???????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1312_ = b[1799:1792];
      256'b??????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1312_ = b[1807:1800];
      256'b?????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1312_ = b[1815:1808];
      256'b????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1312_ = b[1823:1816];
      256'b???????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1312_ = b[1831:1824];
      256'b??????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1312_ = b[1839:1832];
      256'b?????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1312_ = b[1847:1840];
      256'b????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1312_ = b[1855:1848];
      256'b???????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1312_ = b[1863:1856];
      256'b??????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1312_ = b[1871:1864];
      256'b?????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1312_ = b[1879:1872];
      256'b????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1312_ = b[1887:1880];
      256'b???????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1312_ = b[1895:1888];
      256'b??????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1312_ = b[1903:1896];
      256'b?????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1312_ = b[1911:1904];
      256'b????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1312_ = b[1919:1912];
      256'b???????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1312_ = b[1927:1920];
      256'b??????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1312_ = b[1935:1928];
      256'b?????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1312_ = b[1943:1936];
      256'b????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1312_ = b[1951:1944];
      256'b???????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1312_ = b[1959:1952];
      256'b??????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1312_ = b[1967:1960];
      256'b?????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1312_ = b[1975:1968];
      256'b????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1312_ = b[1983:1976];
      256'b???????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1312_ = b[1991:1984];
      256'b??????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1312_ = b[1999:1992];
      256'b?????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1312_ = b[2007:2000];
      256'b????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1312_ = b[2015:2008];
      256'b???1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1312_ = b[2023:2016];
      256'b??1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1312_ = b[2031:2024];
      256'b?1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1312_ = b[2039:2032];
      256'b1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1312_ = b[2047:2040];
      default:
        _1312_ = a;
    endcase
  endfunction
  assign _0257_ = _1312_(\S4_0.S_1.out , 2048'h637c777bf26b6fc53001672bfed7ab76ca82c97dfa5947f0add4a2af9ca472c0b7fd9326363ff7cc34a5e5f171d8311504c723c31896059a071280e2eb27b27509832c1a1b6e5aa0523bd6b329e32f8453d100ed20fcb15b6acbbe394a4c58cfd0efaafb434d338545f9027f503c9fa851a3408f929d38f5bcb6da2110fff3d2cd0c13ec5f974417c4a77e3d645d197360814fdc222a908846eeb814de5e0bdbe0323a0a4906245cc2d3ac629195e479e7c8376d8dd54ea96c56f4ea657aae08ba78252e1ca6b4c6e8dd741f4bbd8b8a703eb5664803f60e613557b986c11d9ee1f8981169d98e949b1e87e9ce5528df8ca1890dbfe6426841992d0fb054bb16, { _0439_, _0438_, _0437_, _0436_, _0435_, _0434_, _0433_, _0432_, _0431_, _0429_, _0428_, _0427_, _0426_, _0425_, _0424_, _0423_, _0422_, _0421_, _0420_, _0418_, _0417_, _0416_, _0415_, _0414_, _0413_, _0412_, _0411_, _0410_, _0409_, _0407_, _0406_, _0405_, _0404_, _0403_, _0402_, _0401_, _0400_, _0399_, _0398_, _0396_, _0395_, _0394_, _0393_, _0392_, _0391_, _0390_, _0389_, _0388_, _0387_, _0385_, _0384_, _0383_, _0382_, _0381_, _0380_, _0379_, _0378_, _0377_, _0376_, _0374_, _0373_, _0372_, _0371_, _0370_, _0369_, _0368_, _0367_, _0366_, _0365_, _0363_, _0362_, _0361_, _0360_, _0359_, _0358_, _0357_, _0356_, _0355_, _0354_, _0352_, _0351_, _0350_, _0349_, _0348_, _0347_, _0346_, _0345_, _0344_, _0343_, _0341_, _0340_, _0339_, _0338_, _0337_, _0336_, _0335_, _0334_, _0333_, _0332_, _0330_, _0329_, _0328_, _0327_, _0326_, _0325_, _0324_, _0323_, _0322_, _0321_, _0319_, _0318_, _0317_, _0316_, _0315_, _0314_, _0313_, _0312_, _0311_, _0310_, _0308_, _0307_, _0306_, _0305_, _0304_, _0303_, _0302_, _0301_, _0300_, _0299_, _0297_, _0296_, _0295_, _0294_, _0293_, _0292_, _0291_, _0290_, _0289_, _0288_, _0287_, _0286_, _0285_, _0284_, _0283_, _0282_, _0281_, _0280_, _0279_, _0278_, _0277_, _0276_, _0275_, _0274_, _0273_, _0272_, _0271_, _0270_, _0269_, _0268_, _0267_, _0266_, _0265_, _0264_, _0263_, _0262_, _0261_, _0260_, _0259_, _0258_, _0513_, _0512_, _0511_, _0510_, _0509_, _0508_, _0507_, _0506_, _0505_, _0504_, _0503_, _0502_, _0501_, _0500_, _0499_, _0498_, _0497_, _0496_, _0495_, _0494_, _0493_, _0492_, _0491_, _0490_, _0489_, _0488_, _0487_, _0486_, _0485_, _0484_, _0483_, _0482_, _0481_, _0480_, _0479_, _0478_, _0477_, _0476_, _0475_, _0474_, _0473_, _0472_, _0471_, _0470_, _0469_, _0468_, _0467_, _0466_, _0465_, _0464_, _0463_, _0462_, _0461_, _0460_, _0459_, _0458_, _0457_, _0456_, _0455_, _0454_, _0453_, _0452_, _0451_, _0450_, _0449_, _0448_, _0447_, _0446_, _0445_, _0444_, _0443_, _0442_, _0441_, _0440_, _0430_, _0419_, _0408_, _0397_, _0386_, _0375_, _0364_, _0353_, _0342_, _0331_, _0320_, _0309_, _0298_ });
  assign _0278_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'h94;
  assign _0279_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'h93;
  assign _0280_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'h92;
  assign _0281_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'h91;
  assign _0282_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'h90;
  assign _0283_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'h8f;
  assign _0284_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'h8e;
  assign _0285_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'h8d;
  assign _0286_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'h8c;
  assign _0287_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'h8b;
  assign _0288_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'h8a;
  assign _0289_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'h89;
  assign _0290_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'h88;
  assign _0291_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'h87;
  assign _0292_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'h86;
  assign _0293_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'h85;
  assign _0294_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'h84;
  assign _0295_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'h83;
  assign _0296_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'h82;
  assign _0297_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'h81;
  assign _0298_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hff;
  assign _0299_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'h80;
  assign _0300_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h7f;
  assign _0301_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h7e;
  assign _0302_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h7d;
  assign _0303_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h7c;
  assign _0304_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h7b;
  assign _0305_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h7a;
  assign _0306_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h79;
  assign _0307_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h78;
  assign _0308_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h77;
  assign _0309_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hfe;
  assign _0310_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h76;
  assign _0311_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h75;
  assign _0312_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h74;
  assign _0313_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h73;
  assign _0314_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h72;
  assign _0315_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h71;
  assign _0316_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h70;
  assign _0317_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h6f;
  assign _0318_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h6e;
  assign _0319_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h6d;
  assign _0320_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hfd;
  assign _0321_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h6c;
  assign _0322_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h6b;
  assign _0323_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h6a;
  assign _0324_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h69;
  assign _0325_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h68;
  assign _0326_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h67;
  assign _0327_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h66;
  assign _0328_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h65;
  assign _0329_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h64;
  assign _0330_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h63;
  assign _0331_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hfc;
  assign _0332_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h62;
  assign _0333_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h61;
  assign _0334_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h60;
  assign _0335_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h5f;
  assign _0336_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h5e;
  assign _0337_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h5d;
  assign _0338_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h5c;
  assign _0339_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h5b;
  assign _0340_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h5a;
  assign _0341_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h59;
  assign _0342_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hfb;
  assign _0343_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h58;
  assign _0344_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h57;
  assign _0345_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h56;
  assign _0346_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h55;
  assign _0347_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h54;
  assign _0348_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h53;
  assign _0349_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h52;
  assign _0350_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h51;
  assign _0351_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h50;
  assign _0352_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h4f;
  assign _0353_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hfa;
  assign _0354_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h4e;
  assign _0355_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h4d;
  assign _0356_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h4c;
  assign _0357_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h4b;
  assign _0358_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h4a;
  assign _0359_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h49;
  assign _0360_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h48;
  assign _0361_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h47;
  assign _0362_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h46;
  assign _0363_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h45;
  assign _0364_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hf9;
  assign _0365_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h44;
  assign _0366_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h43;
  assign _0367_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h42;
  assign _0368_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h41;
  assign _0369_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h40;
  assign _0370_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 6'h3f;
  assign _0371_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 6'h3e;
  assign _0372_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 6'h3d;
  assign _0373_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 6'h3c;
  assign _0374_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 6'h3b;
  assign _0375_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hf8;
  assign _0376_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 6'h3a;
  assign _0377_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 6'h39;
  assign _0378_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 6'h38;
  assign _0379_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 6'h37;
  assign _0380_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 6'h36;
  assign _0381_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 6'h35;
  assign _0382_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 6'h34;
  assign _0383_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 6'h33;
  assign _0384_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 6'h32;
  assign _0385_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 6'h31;
  assign _0386_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hf7;
  assign _0387_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 6'h30;
  assign _0388_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 6'h2f;
  assign _0389_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 6'h2e;
  assign _0390_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 6'h2d;
  assign _0391_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 6'h2c;
  assign _0392_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 6'h2b;
  assign _0393_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 6'h2a;
  assign _0394_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 6'h29;
  assign _0395_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 6'h28;
  assign _0396_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 6'h27;
  assign _0397_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hf6;
  assign _0398_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 6'h26;
  assign _0399_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 6'h25;
  assign _0400_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 6'h24;
  assign _0401_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 6'h23;
  assign _0402_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 6'h22;
  assign _0403_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 6'h21;
  assign _0404_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 6'h20;
  assign _0405_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 5'h1f;
  assign _0406_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 5'h1e;
  assign _0407_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 5'h1d;
  assign _0408_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hf5;
  assign _0409_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 5'h1c;
  assign _0410_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 5'h1b;
  assign _0411_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 5'h1a;
  assign _0412_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 5'h19;
  assign _0413_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 5'h18;
  assign _0414_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 5'h17;
  assign _0415_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 5'h16;
  assign _0416_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 5'h15;
  assign _0417_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 5'h14;
  assign _0418_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 5'h13;
  assign _0419_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hf4;
  assign _0420_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 5'h12;
  assign _0421_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 5'h11;
  assign _0422_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 5'h10;
  assign _0423_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 4'hf;
  assign _0424_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 4'he;
  assign _0425_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 4'hd;
  assign _0426_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 4'hc;
  assign _0427_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 4'hb;
  assign _0428_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 4'ha;
  assign _0429_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 4'h9;
  assign _0430_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hf3;
  assign _0431_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 4'h8;
  assign _0432_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 3'h7;
  assign _0433_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 3'h6;
  assign _0434_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 3'h5;
  assign _0435_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 3'h4;
  assign _0436_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 2'h3;
  assign _0437_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 2'h2;
  assign _0438_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 1'h1;
  assign _0439_ = ! (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) in[15:8];
  assign _0440_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hf2;
  assign _0441_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hf1;
  assign _0442_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hf0;
  assign _0443_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hef;
  assign _0444_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hee;
  assign _0445_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hed;
  assign _0446_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hec;
  assign _0447_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'heb;
  assign _0448_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hea;
  assign _0449_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'he9;
  assign _0450_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'he8;
  assign _0451_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'he7;
  assign _0452_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'he6;
  assign _0453_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'he5;
  assign _0454_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'he4;
  assign _0455_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'he3;
  assign _0456_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'he2;
  assign _0457_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'he1;
  assign _0458_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'he0;
  assign _0459_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hdf;
  assign _0460_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hde;
  assign _0461_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hdd;
  assign _0462_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hdc;
  assign _0463_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hdb;
  assign _0464_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hda;
  assign _0465_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hd9;
  assign _0466_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hd8;
  assign _0467_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hd7;
  assign _0468_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hd6;
  assign _0469_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hd5;
  assign _0470_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hd4;
  assign _0471_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hd3;
  assign _0472_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hd2;
  assign _0473_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hd1;
  assign _0474_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hd0;
  assign _0475_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hcf;
  assign _0476_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hce;
  assign _0477_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hcd;
  assign _0478_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hcc;
  assign _0479_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hcb;
  assign _0480_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hca;
  assign _0481_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hc9;
  assign _0482_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hc8;
  assign _0483_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hc7;
  assign _0484_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hc6;
  assign _0485_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hc5;
  assign _0486_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hc4;
  assign _0487_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hc3;
  assign _0488_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hc2;
  assign _0489_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hc1;
  assign _0490_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hc0;
  assign _0491_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hbf;
  assign _0492_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hbe;
  assign _0493_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hbd;
  assign _0494_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hbc;
  assign _0495_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hbb;
  assign _0496_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hba;
  assign _0497_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hb9;
  assign _0498_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hb8;
  assign _0499_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hb7;
  assign _0500_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hb6;
  assign _0501_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hb5;
  assign _0502_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hb4;
  assign _0503_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hb3;
  assign _0504_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hb2;
  assign _0505_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hb1;
  assign _0506_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hb0;
  assign _0507_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'haf;
  assign _0508_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hae;
  assign _0509_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'had;
  assign _0510_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hac;
  assign _0511_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hab;
  assign _0512_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'haa;
  assign _0513_ = in[15:8] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'ha9;
  always @(posedge clk)
      \S4_0.S_2.out  <= _0514_;
  assign _0515_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'ha8;
  assign _0516_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'ha7;
  assign _0517_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'ha6;
  assign _0518_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'ha5;
  assign _0519_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'ha4;
  assign _0520_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'ha3;
  assign _0521_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'ha2;
  assign _0522_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'ha1;
  assign _0523_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'ha0;
  assign _0524_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'h9f;
  assign _0525_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'h9e;
  assign _0526_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'h9d;
  assign _0527_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'h9c;
  assign _0528_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'h9b;
  assign _0529_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'h9a;
  assign _0530_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'h99;
  assign _0531_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'h98;
  assign _0532_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'h97;
  assign _0533_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'h96;
  assign _0534_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'h95;
  function [7:0] _1570_;
    input [7:0] a;
    input [2047:0] b;
    input [255:0] s;
    (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *)
    (* parallel_case *)
    casez (s)
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1:
        _1570_ = b[7:0];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?:
        _1570_ = b[15:8];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??:
        _1570_ = b[23:16];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???:
        _1570_ = b[31:24];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????:
        _1570_ = b[39:32];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????:
        _1570_ = b[47:40];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????:
        _1570_ = b[55:48];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????:
        _1570_ = b[63:56];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????:
        _1570_ = b[71:64];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????:
        _1570_ = b[79:72];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????:
        _1570_ = b[87:80];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????:
        _1570_ = b[95:88];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????:
        _1570_ = b[103:96];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????:
        _1570_ = b[111:104];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????:
        _1570_ = b[119:112];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????:
        _1570_ = b[127:120];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????:
        _1570_ = b[135:128];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????:
        _1570_ = b[143:136];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????:
        _1570_ = b[151:144];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????:
        _1570_ = b[159:152];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????:
        _1570_ = b[167:160];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????:
        _1570_ = b[175:168];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????:
        _1570_ = b[183:176];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????:
        _1570_ = b[191:184];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????:
        _1570_ = b[199:192];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????:
        _1570_ = b[207:200];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????:
        _1570_ = b[215:208];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????:
        _1570_ = b[223:216];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????:
        _1570_ = b[231:224];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????:
        _1570_ = b[239:232];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????:
        _1570_ = b[247:240];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????:
        _1570_ = b[255:248];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????:
        _1570_ = b[263:256];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????:
        _1570_ = b[271:264];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????:
        _1570_ = b[279:272];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????:
        _1570_ = b[287:280];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????:
        _1570_ = b[295:288];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????:
        _1570_ = b[303:296];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????:
        _1570_ = b[311:304];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????:
        _1570_ = b[319:312];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????:
        _1570_ = b[327:320];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????:
        _1570_ = b[335:328];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????:
        _1570_ = b[343:336];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????:
        _1570_ = b[351:344];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????:
        _1570_ = b[359:352];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????:
        _1570_ = b[367:360];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????:
        _1570_ = b[375:368];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????:
        _1570_ = b[383:376];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????:
        _1570_ = b[391:384];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????:
        _1570_ = b[399:392];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????:
        _1570_ = b[407:400];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????:
        _1570_ = b[415:408];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????:
        _1570_ = b[423:416];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????:
        _1570_ = b[431:424];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????:
        _1570_ = b[439:432];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????:
        _1570_ = b[447:440];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????:
        _1570_ = b[455:448];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????:
        _1570_ = b[463:456];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????:
        _1570_ = b[471:464];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????:
        _1570_ = b[479:472];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????:
        _1570_ = b[487:480];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????:
        _1570_ = b[495:488];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????:
        _1570_ = b[503:496];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????:
        _1570_ = b[511:504];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????:
        _1570_ = b[519:512];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????:
        _1570_ = b[527:520];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????:
        _1570_ = b[535:528];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????:
        _1570_ = b[543:536];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????:
        _1570_ = b[551:544];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????:
        _1570_ = b[559:552];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????:
        _1570_ = b[567:560];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????:
        _1570_ = b[575:568];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????:
        _1570_ = b[583:576];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????:
        _1570_ = b[591:584];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????:
        _1570_ = b[599:592];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????:
        _1570_ = b[607:600];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????:
        _1570_ = b[615:608];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????:
        _1570_ = b[623:616];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????:
        _1570_ = b[631:624];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????:
        _1570_ = b[639:632];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????:
        _1570_ = b[647:640];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????:
        _1570_ = b[655:648];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????:
        _1570_ = b[663:656];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????:
        _1570_ = b[671:664];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????:
        _1570_ = b[679:672];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????:
        _1570_ = b[687:680];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????:
        _1570_ = b[695:688];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????:
        _1570_ = b[703:696];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????:
        _1570_ = b[711:704];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????:
        _1570_ = b[719:712];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????:
        _1570_ = b[727:720];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????:
        _1570_ = b[735:728];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????:
        _1570_ = b[743:736];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????:
        _1570_ = b[751:744];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????:
        _1570_ = b[759:752];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????:
        _1570_ = b[767:760];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????:
        _1570_ = b[775:768];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????:
        _1570_ = b[783:776];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????:
        _1570_ = b[791:784];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????:
        _1570_ = b[799:792];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1570_ = b[807:800];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1570_ = b[815:808];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1570_ = b[823:816];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1570_ = b[831:824];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1570_ = b[839:832];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1570_ = b[847:840];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1570_ = b[855:848];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1570_ = b[863:856];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1570_ = b[871:864];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1570_ = b[879:872];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1570_ = b[887:880];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1570_ = b[895:888];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1570_ = b[903:896];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1570_ = b[911:904];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1570_ = b[919:912];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1570_ = b[927:920];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1570_ = b[935:928];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1570_ = b[943:936];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1570_ = b[951:944];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1570_ = b[959:952];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1570_ = b[967:960];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1570_ = b[975:968];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1570_ = b[983:976];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1570_ = b[991:984];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1570_ = b[999:992];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1570_ = b[1007:1000];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1570_ = b[1015:1008];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1570_ = b[1023:1016];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1570_ = b[1031:1024];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1570_ = b[1039:1032];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1570_ = b[1047:1040];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1570_ = b[1055:1048];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1570_ = b[1063:1056];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1570_ = b[1071:1064];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1570_ = b[1079:1072];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1570_ = b[1087:1080];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1570_ = b[1095:1088];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1570_ = b[1103:1096];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1570_ = b[1111:1104];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1570_ = b[1119:1112];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1570_ = b[1127:1120];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1570_ = b[1135:1128];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1570_ = b[1143:1136];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1570_ = b[1151:1144];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1570_ = b[1159:1152];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1570_ = b[1167:1160];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1570_ = b[1175:1168];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1570_ = b[1183:1176];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1570_ = b[1191:1184];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1570_ = b[1199:1192];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1570_ = b[1207:1200];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1570_ = b[1215:1208];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1570_ = b[1223:1216];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1570_ = b[1231:1224];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1570_ = b[1239:1232];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1570_ = b[1247:1240];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1570_ = b[1255:1248];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1570_ = b[1263:1256];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1570_ = b[1271:1264];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1570_ = b[1279:1272];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1570_ = b[1287:1280];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1570_ = b[1295:1288];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1570_ = b[1303:1296];
      256'b????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1570_ = b[1311:1304];
      256'b???????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1570_ = b[1319:1312];
      256'b??????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1570_ = b[1327:1320];
      256'b?????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1570_ = b[1335:1328];
      256'b????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1570_ = b[1343:1336];
      256'b???????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1570_ = b[1351:1344];
      256'b??????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1570_ = b[1359:1352];
      256'b?????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1570_ = b[1367:1360];
      256'b????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1570_ = b[1375:1368];
      256'b???????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1570_ = b[1383:1376];
      256'b??????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1570_ = b[1391:1384];
      256'b?????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1570_ = b[1399:1392];
      256'b????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1570_ = b[1407:1400];
      256'b???????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1570_ = b[1415:1408];
      256'b??????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1570_ = b[1423:1416];
      256'b?????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1570_ = b[1431:1424];
      256'b????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1570_ = b[1439:1432];
      256'b???????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1570_ = b[1447:1440];
      256'b??????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1570_ = b[1455:1448];
      256'b?????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1570_ = b[1463:1456];
      256'b????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1570_ = b[1471:1464];
      256'b???????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1570_ = b[1479:1472];
      256'b??????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1570_ = b[1487:1480];
      256'b?????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1570_ = b[1495:1488];
      256'b????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1570_ = b[1503:1496];
      256'b???????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1570_ = b[1511:1504];
      256'b??????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1570_ = b[1519:1512];
      256'b?????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1570_ = b[1527:1520];
      256'b????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1570_ = b[1535:1528];
      256'b???????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1570_ = b[1543:1536];
      256'b??????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1570_ = b[1551:1544];
      256'b?????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1570_ = b[1559:1552];
      256'b????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1570_ = b[1567:1560];
      256'b???????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1570_ = b[1575:1568];
      256'b??????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1570_ = b[1583:1576];
      256'b?????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1570_ = b[1591:1584];
      256'b????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1570_ = b[1599:1592];
      256'b???????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1570_ = b[1607:1600];
      256'b??????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1570_ = b[1615:1608];
      256'b?????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1570_ = b[1623:1616];
      256'b????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1570_ = b[1631:1624];
      256'b???????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1570_ = b[1639:1632];
      256'b??????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1570_ = b[1647:1640];
      256'b?????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1570_ = b[1655:1648];
      256'b????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1570_ = b[1663:1656];
      256'b???????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1570_ = b[1671:1664];
      256'b??????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1570_ = b[1679:1672];
      256'b?????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1570_ = b[1687:1680];
      256'b????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1570_ = b[1695:1688];
      256'b???????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1570_ = b[1703:1696];
      256'b??????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1570_ = b[1711:1704];
      256'b?????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1570_ = b[1719:1712];
      256'b????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1570_ = b[1727:1720];
      256'b???????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1570_ = b[1735:1728];
      256'b??????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1570_ = b[1743:1736];
      256'b?????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1570_ = b[1751:1744];
      256'b????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1570_ = b[1759:1752];
      256'b???????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1570_ = b[1767:1760];
      256'b??????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1570_ = b[1775:1768];
      256'b?????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1570_ = b[1783:1776];
      256'b????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1570_ = b[1791:1784];
      256'b???????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1570_ = b[1799:1792];
      256'b??????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1570_ = b[1807:1800];
      256'b?????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1570_ = b[1815:1808];
      256'b????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1570_ = b[1823:1816];
      256'b???????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1570_ = b[1831:1824];
      256'b??????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1570_ = b[1839:1832];
      256'b?????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1570_ = b[1847:1840];
      256'b????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1570_ = b[1855:1848];
      256'b???????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1570_ = b[1863:1856];
      256'b??????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1570_ = b[1871:1864];
      256'b?????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1570_ = b[1879:1872];
      256'b????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1570_ = b[1887:1880];
      256'b???????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1570_ = b[1895:1888];
      256'b??????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1570_ = b[1903:1896];
      256'b?????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1570_ = b[1911:1904];
      256'b????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1570_ = b[1919:1912];
      256'b???????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1570_ = b[1927:1920];
      256'b??????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1570_ = b[1935:1928];
      256'b?????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1570_ = b[1943:1936];
      256'b????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1570_ = b[1951:1944];
      256'b???????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1570_ = b[1959:1952];
      256'b??????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1570_ = b[1967:1960];
      256'b?????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1570_ = b[1975:1968];
      256'b????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1570_ = b[1983:1976];
      256'b???????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1570_ = b[1991:1984];
      256'b??????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1570_ = b[1999:1992];
      256'b?????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1570_ = b[2007:2000];
      256'b????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1570_ = b[2015:2008];
      256'b???1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1570_ = b[2023:2016];
      256'b??1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1570_ = b[2031:2024];
      256'b?1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1570_ = b[2039:2032];
      256'b1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1570_ = b[2047:2040];
      default:
        _1570_ = a;
    endcase
  endfunction
  assign _0514_ = _1570_(\S4_0.S_2.out , 2048'h637c777bf26b6fc53001672bfed7ab76ca82c97dfa5947f0add4a2af9ca472c0b7fd9326363ff7cc34a5e5f171d8311504c723c31896059a071280e2eb27b27509832c1a1b6e5aa0523bd6b329e32f8453d100ed20fcb15b6acbbe394a4c58cfd0efaafb434d338545f9027f503c9fa851a3408f929d38f5bcb6da2110fff3d2cd0c13ec5f974417c4a77e3d645d197360814fdc222a908846eeb814de5e0bdbe0323a0a4906245cc2d3ac629195e479e7c8376d8dd54ea96c56f4ea657aae08ba78252e1ca6b4c6e8dd741f4bbd8b8a703eb5664803f60e613557b986c11d9ee1f8981169d98e949b1e87e9ce5528df8ca1890dbfe6426841992d0fb054bb16, { _0696_, _0695_, _0694_, _0693_, _0692_, _0691_, _0690_, _0689_, _0688_, _0686_, _0685_, _0684_, _0683_, _0682_, _0681_, _0680_, _0679_, _0678_, _0677_, _0675_, _0674_, _0673_, _0672_, _0671_, _0670_, _0669_, _0668_, _0667_, _0666_, _0664_, _0663_, _0662_, _0661_, _0660_, _0659_, _0658_, _0657_, _0656_, _0655_, _0653_, _0652_, _0651_, _0650_, _0649_, _0648_, _0647_, _0646_, _0645_, _0644_, _0642_, _0641_, _0640_, _0639_, _0638_, _0637_, _0636_, _0635_, _0634_, _0633_, _0631_, _0630_, _0629_, _0628_, _0627_, _0626_, _0625_, _0624_, _0623_, _0622_, _0620_, _0619_, _0618_, _0617_, _0616_, _0615_, _0614_, _0613_, _0612_, _0611_, _0609_, _0608_, _0607_, _0606_, _0605_, _0604_, _0603_, _0602_, _0601_, _0600_, _0598_, _0597_, _0596_, _0595_, _0594_, _0593_, _0592_, _0591_, _0590_, _0589_, _0587_, _0586_, _0585_, _0584_, _0583_, _0582_, _0581_, _0580_, _0579_, _0578_, _0576_, _0575_, _0574_, _0573_, _0572_, _0571_, _0570_, _0569_, _0568_, _0567_, _0565_, _0564_, _0563_, _0562_, _0561_, _0560_, _0559_, _0558_, _0557_, _0556_, _0554_, _0553_, _0552_, _0551_, _0550_, _0549_, _0548_, _0547_, _0546_, _0545_, _0544_, _0543_, _0542_, _0541_, _0540_, _0539_, _0538_, _0537_, _0536_, _0535_, _0534_, _0533_, _0532_, _0531_, _0530_, _0529_, _0528_, _0527_, _0526_, _0525_, _0524_, _0523_, _0522_, _0521_, _0520_, _0519_, _0518_, _0517_, _0516_, _0515_, _0770_, _0769_, _0768_, _0767_, _0766_, _0765_, _0764_, _0763_, _0762_, _0761_, _0760_, _0759_, _0758_, _0757_, _0756_, _0755_, _0754_, _0753_, _0752_, _0751_, _0750_, _0749_, _0748_, _0747_, _0746_, _0745_, _0744_, _0743_, _0742_, _0741_, _0740_, _0739_, _0738_, _0737_, _0736_, _0735_, _0734_, _0733_, _0732_, _0731_, _0730_, _0729_, _0728_, _0727_, _0726_, _0725_, _0724_, _0723_, _0722_, _0721_, _0720_, _0719_, _0718_, _0717_, _0716_, _0715_, _0714_, _0713_, _0712_, _0711_, _0710_, _0709_, _0708_, _0707_, _0706_, _0705_, _0704_, _0703_, _0702_, _0701_, _0700_, _0699_, _0698_, _0697_, _0687_, _0676_, _0665_, _0654_, _0643_, _0632_, _0621_, _0610_, _0599_, _0588_, _0577_, _0566_, _0555_ });
  assign _0535_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'h94;
  assign _0536_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'h93;
  assign _0537_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'h92;
  assign _0538_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'h91;
  assign _0539_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'h90;
  assign _0540_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'h8f;
  assign _0541_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'h8e;
  assign _0542_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'h8d;
  assign _0543_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'h8c;
  assign _0544_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'h8b;
  assign _0545_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'h8a;
  assign _0546_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'h89;
  assign _0547_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'h88;
  assign _0548_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'h87;
  assign _0549_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'h86;
  assign _0550_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'h85;
  assign _0551_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'h84;
  assign _0552_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'h83;
  assign _0553_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'h82;
  assign _0554_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'h81;
  assign _0555_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hff;
  assign _0556_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'h80;
  assign _0557_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h7f;
  assign _0558_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h7e;
  assign _0559_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h7d;
  assign _0560_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h7c;
  assign _0561_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h7b;
  assign _0562_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h7a;
  assign _0563_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h79;
  assign _0564_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h78;
  assign _0565_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h77;
  assign _0566_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hfe;
  assign _0567_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h76;
  assign _0568_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h75;
  assign _0569_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h74;
  assign _0570_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h73;
  assign _0571_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h72;
  assign _0572_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h71;
  assign _0573_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h70;
  assign _0574_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h6f;
  assign _0575_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h6e;
  assign _0576_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h6d;
  assign _0577_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hfd;
  assign _0578_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h6c;
  assign _0579_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h6b;
  assign _0580_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h6a;
  assign _0581_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h69;
  assign _0582_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h68;
  assign _0583_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h67;
  assign _0584_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h66;
  assign _0585_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h65;
  assign _0586_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h64;
  assign _0587_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h63;
  assign _0588_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hfc;
  assign _0589_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h62;
  assign _0590_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h61;
  assign _0591_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h60;
  assign _0592_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h5f;
  assign _0593_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h5e;
  assign _0594_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h5d;
  assign _0595_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h5c;
  assign _0596_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h5b;
  assign _0597_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h5a;
  assign _0598_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h59;
  assign _0599_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hfb;
  assign _0600_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h58;
  assign _0601_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h57;
  assign _0602_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h56;
  assign _0603_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h55;
  assign _0604_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h54;
  assign _0605_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h53;
  assign _0606_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h52;
  assign _0607_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h51;
  assign _0608_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h50;
  assign _0609_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h4f;
  assign _0610_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hfa;
  assign _0611_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h4e;
  assign _0612_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h4d;
  assign _0613_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h4c;
  assign _0614_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h4b;
  assign _0615_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h4a;
  assign _0616_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h49;
  assign _0617_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h48;
  assign _0618_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h47;
  assign _0619_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h46;
  assign _0620_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h45;
  assign _0621_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hf9;
  assign _0622_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h44;
  assign _0623_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h43;
  assign _0624_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h42;
  assign _0625_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h41;
  assign _0626_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h40;
  assign _0627_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 6'h3f;
  assign _0628_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 6'h3e;
  assign _0629_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 6'h3d;
  assign _0630_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 6'h3c;
  assign _0631_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 6'h3b;
  assign _0632_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hf8;
  assign _0633_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 6'h3a;
  assign _0634_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 6'h39;
  assign _0635_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 6'h38;
  assign _0636_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 6'h37;
  assign _0637_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 6'h36;
  assign _0638_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 6'h35;
  assign _0639_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 6'h34;
  assign _0640_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 6'h33;
  assign _0641_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 6'h32;
  assign _0642_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 6'h31;
  assign _0643_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hf7;
  assign _0644_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 6'h30;
  assign _0645_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 6'h2f;
  assign _0646_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 6'h2e;
  assign _0647_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 6'h2d;
  assign _0648_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 6'h2c;
  assign _0649_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 6'h2b;
  assign _0650_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 6'h2a;
  assign _0651_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 6'h29;
  assign _0652_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 6'h28;
  assign _0653_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 6'h27;
  assign _0654_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hf6;
  assign _0655_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 6'h26;
  assign _0656_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 6'h25;
  assign _0657_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 6'h24;
  assign _0658_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 6'h23;
  assign _0659_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 6'h22;
  assign _0660_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 6'h21;
  assign _0661_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 6'h20;
  assign _0662_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 5'h1f;
  assign _0663_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 5'h1e;
  assign _0664_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 5'h1d;
  assign _0665_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hf5;
  assign _0666_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 5'h1c;
  assign _0667_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 5'h1b;
  assign _0668_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 5'h1a;
  assign _0669_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 5'h19;
  assign _0670_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 5'h18;
  assign _0671_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 5'h17;
  assign _0672_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 5'h16;
  assign _0673_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 5'h15;
  assign _0674_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 5'h14;
  assign _0675_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 5'h13;
  assign _0676_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hf4;
  assign _0677_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 5'h12;
  assign _0678_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 5'h11;
  assign _0679_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 5'h10;
  assign _0680_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 4'hf;
  assign _0681_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 4'he;
  assign _0682_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 4'hd;
  assign _0683_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 4'hc;
  assign _0684_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 4'hb;
  assign _0685_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 4'ha;
  assign _0686_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 4'h9;
  assign _0687_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hf3;
  assign _0688_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 4'h8;
  assign _0689_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 3'h7;
  assign _0690_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 3'h6;
  assign _0691_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 3'h5;
  assign _0692_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 3'h4;
  assign _0693_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 2'h3;
  assign _0694_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 2'h2;
  assign _0695_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 1'h1;
  assign _0696_ = ! (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) in[7:0];
  assign _0697_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hf2;
  assign _0698_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hf1;
  assign _0699_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hf0;
  assign _0700_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hef;
  assign _0701_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hee;
  assign _0702_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hed;
  assign _0703_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hec;
  assign _0704_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'heb;
  assign _0705_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hea;
  assign _0706_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'he9;
  assign _0707_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'he8;
  assign _0708_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'he7;
  assign _0709_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'he6;
  assign _0710_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'he5;
  assign _0711_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'he4;
  assign _0712_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'he3;
  assign _0713_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'he2;
  assign _0714_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'he1;
  assign _0715_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'he0;
  assign _0716_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hdf;
  assign _0717_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hde;
  assign _0718_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hdd;
  assign _0719_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hdc;
  assign _0720_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hdb;
  assign _0721_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hda;
  assign _0722_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hd9;
  assign _0723_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hd8;
  assign _0724_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hd7;
  assign _0725_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hd6;
  assign _0726_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hd5;
  assign _0727_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hd4;
  assign _0728_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hd3;
  assign _0729_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hd2;
  assign _0730_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hd1;
  assign _0731_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hd0;
  assign _0732_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hcf;
  assign _0733_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hce;
  assign _0734_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hcd;
  assign _0735_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hcc;
  assign _0736_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hcb;
  assign _0737_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hca;
  assign _0738_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hc9;
  assign _0739_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hc8;
  assign _0740_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hc7;
  assign _0741_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hc6;
  assign _0742_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hc5;
  assign _0743_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hc4;
  assign _0744_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hc3;
  assign _0745_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hc2;
  assign _0746_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hc1;
  assign _0747_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hc0;
  assign _0748_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hbf;
  assign _0749_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hbe;
  assign _0750_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hbd;
  assign _0751_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hbc;
  assign _0752_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hbb;
  assign _0753_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hba;
  assign _0754_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hb9;
  assign _0755_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hb8;
  assign _0756_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hb7;
  assign _0757_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hb6;
  assign _0758_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hb5;
  assign _0759_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hb4;
  assign _0760_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hb3;
  assign _0761_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hb2;
  assign _0762_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hb1;
  assign _0763_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hb0;
  assign _0764_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'haf;
  assign _0765_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hae;
  assign _0766_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'had;
  assign _0767_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hac;
  assign _0768_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hab;
  assign _0769_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'haa;
  assign _0770_ = in[7:0] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'ha9;
  always @(posedge clk)
      \S4_0.S_3.out  <= _0771_;
  assign _0772_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'ha8;
  assign _0773_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'ha7;
  assign _0774_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'ha6;
  assign _0775_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'ha5;
  assign _0776_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'ha4;
  assign _0777_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'ha3;
  assign _0778_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'ha2;
  assign _0779_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'ha1;
  assign _0780_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'ha0;
  assign _0781_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'h9f;
  assign _0782_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'h9e;
  assign _0783_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'h9d;
  assign _0784_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'h9c;
  assign _0785_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'h9b;
  assign _0786_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'h9a;
  assign _0787_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'h99;
  assign _0788_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'h98;
  assign _0789_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'h97;
  assign _0790_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'h96;
  assign _0791_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'h95;
  function [7:0] _1828_;
    input [7:0] a;
    input [2047:0] b;
    input [255:0] s;
    (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *)
    (* parallel_case *)
    casez (s)
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1:
        _1828_ = b[7:0];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?:
        _1828_ = b[15:8];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??:
        _1828_ = b[23:16];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???:
        _1828_ = b[31:24];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????:
        _1828_ = b[39:32];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????:
        _1828_ = b[47:40];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????:
        _1828_ = b[55:48];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????:
        _1828_ = b[63:56];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????:
        _1828_ = b[71:64];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????:
        _1828_ = b[79:72];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????:
        _1828_ = b[87:80];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????:
        _1828_ = b[95:88];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????:
        _1828_ = b[103:96];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????:
        _1828_ = b[111:104];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????:
        _1828_ = b[119:112];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????:
        _1828_ = b[127:120];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????:
        _1828_ = b[135:128];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????:
        _1828_ = b[143:136];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????:
        _1828_ = b[151:144];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????:
        _1828_ = b[159:152];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????:
        _1828_ = b[167:160];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????:
        _1828_ = b[175:168];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????:
        _1828_ = b[183:176];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????:
        _1828_ = b[191:184];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????:
        _1828_ = b[199:192];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????:
        _1828_ = b[207:200];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????:
        _1828_ = b[215:208];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????:
        _1828_ = b[223:216];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????:
        _1828_ = b[231:224];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????:
        _1828_ = b[239:232];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????:
        _1828_ = b[247:240];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????:
        _1828_ = b[255:248];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????:
        _1828_ = b[263:256];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????:
        _1828_ = b[271:264];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????:
        _1828_ = b[279:272];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????:
        _1828_ = b[287:280];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????:
        _1828_ = b[295:288];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????:
        _1828_ = b[303:296];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????:
        _1828_ = b[311:304];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????:
        _1828_ = b[319:312];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????:
        _1828_ = b[327:320];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????:
        _1828_ = b[335:328];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????:
        _1828_ = b[343:336];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????:
        _1828_ = b[351:344];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????:
        _1828_ = b[359:352];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????:
        _1828_ = b[367:360];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????:
        _1828_ = b[375:368];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????:
        _1828_ = b[383:376];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????:
        _1828_ = b[391:384];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????:
        _1828_ = b[399:392];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????:
        _1828_ = b[407:400];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????:
        _1828_ = b[415:408];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????:
        _1828_ = b[423:416];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????:
        _1828_ = b[431:424];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????:
        _1828_ = b[439:432];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????:
        _1828_ = b[447:440];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????:
        _1828_ = b[455:448];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????:
        _1828_ = b[463:456];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????:
        _1828_ = b[471:464];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????:
        _1828_ = b[479:472];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????:
        _1828_ = b[487:480];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????:
        _1828_ = b[495:488];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????:
        _1828_ = b[503:496];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????:
        _1828_ = b[511:504];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????:
        _1828_ = b[519:512];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????:
        _1828_ = b[527:520];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????:
        _1828_ = b[535:528];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????:
        _1828_ = b[543:536];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????:
        _1828_ = b[551:544];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????:
        _1828_ = b[559:552];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????:
        _1828_ = b[567:560];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????:
        _1828_ = b[575:568];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????:
        _1828_ = b[583:576];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????:
        _1828_ = b[591:584];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????:
        _1828_ = b[599:592];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????:
        _1828_ = b[607:600];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????:
        _1828_ = b[615:608];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????:
        _1828_ = b[623:616];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????:
        _1828_ = b[631:624];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????:
        _1828_ = b[639:632];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????:
        _1828_ = b[647:640];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????:
        _1828_ = b[655:648];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????:
        _1828_ = b[663:656];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????:
        _1828_ = b[671:664];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????:
        _1828_ = b[679:672];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????:
        _1828_ = b[687:680];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????:
        _1828_ = b[695:688];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????:
        _1828_ = b[703:696];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????:
        _1828_ = b[711:704];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????:
        _1828_ = b[719:712];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????:
        _1828_ = b[727:720];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????:
        _1828_ = b[735:728];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????:
        _1828_ = b[743:736];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????:
        _1828_ = b[751:744];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????:
        _1828_ = b[759:752];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????:
        _1828_ = b[767:760];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????:
        _1828_ = b[775:768];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????:
        _1828_ = b[783:776];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????:
        _1828_ = b[791:784];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????:
        _1828_ = b[799:792];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1828_ = b[807:800];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1828_ = b[815:808];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1828_ = b[823:816];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1828_ = b[831:824];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1828_ = b[839:832];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1828_ = b[847:840];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1828_ = b[855:848];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1828_ = b[863:856];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1828_ = b[871:864];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1828_ = b[879:872];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1828_ = b[887:880];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1828_ = b[895:888];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1828_ = b[903:896];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1828_ = b[911:904];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1828_ = b[919:912];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1828_ = b[927:920];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1828_ = b[935:928];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1828_ = b[943:936];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1828_ = b[951:944];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1828_ = b[959:952];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1828_ = b[967:960];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1828_ = b[975:968];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1828_ = b[983:976];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1828_ = b[991:984];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1828_ = b[999:992];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1828_ = b[1007:1000];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1828_ = b[1015:1008];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1828_ = b[1023:1016];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1828_ = b[1031:1024];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1828_ = b[1039:1032];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1828_ = b[1047:1040];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1828_ = b[1055:1048];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1828_ = b[1063:1056];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1828_ = b[1071:1064];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1828_ = b[1079:1072];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1828_ = b[1087:1080];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1828_ = b[1095:1088];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1828_ = b[1103:1096];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1828_ = b[1111:1104];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1828_ = b[1119:1112];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1828_ = b[1127:1120];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1828_ = b[1135:1128];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1828_ = b[1143:1136];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1828_ = b[1151:1144];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1828_ = b[1159:1152];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1828_ = b[1167:1160];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1828_ = b[1175:1168];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1828_ = b[1183:1176];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1828_ = b[1191:1184];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1828_ = b[1199:1192];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1828_ = b[1207:1200];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1828_ = b[1215:1208];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1828_ = b[1223:1216];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1828_ = b[1231:1224];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1828_ = b[1239:1232];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1828_ = b[1247:1240];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1828_ = b[1255:1248];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1828_ = b[1263:1256];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1828_ = b[1271:1264];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1828_ = b[1279:1272];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1828_ = b[1287:1280];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1828_ = b[1295:1288];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1828_ = b[1303:1296];
      256'b????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1828_ = b[1311:1304];
      256'b???????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1828_ = b[1319:1312];
      256'b??????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1828_ = b[1327:1320];
      256'b?????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1828_ = b[1335:1328];
      256'b????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1828_ = b[1343:1336];
      256'b???????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1828_ = b[1351:1344];
      256'b??????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1828_ = b[1359:1352];
      256'b?????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1828_ = b[1367:1360];
      256'b????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1828_ = b[1375:1368];
      256'b???????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1828_ = b[1383:1376];
      256'b??????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1828_ = b[1391:1384];
      256'b?????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1828_ = b[1399:1392];
      256'b????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1828_ = b[1407:1400];
      256'b???????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1828_ = b[1415:1408];
      256'b??????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1828_ = b[1423:1416];
      256'b?????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1828_ = b[1431:1424];
      256'b????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1828_ = b[1439:1432];
      256'b???????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1828_ = b[1447:1440];
      256'b??????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1828_ = b[1455:1448];
      256'b?????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1828_ = b[1463:1456];
      256'b????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1828_ = b[1471:1464];
      256'b???????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1828_ = b[1479:1472];
      256'b??????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1828_ = b[1487:1480];
      256'b?????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1828_ = b[1495:1488];
      256'b????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1828_ = b[1503:1496];
      256'b???????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1828_ = b[1511:1504];
      256'b??????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1828_ = b[1519:1512];
      256'b?????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1828_ = b[1527:1520];
      256'b????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1828_ = b[1535:1528];
      256'b???????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1828_ = b[1543:1536];
      256'b??????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1828_ = b[1551:1544];
      256'b?????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1828_ = b[1559:1552];
      256'b????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1828_ = b[1567:1560];
      256'b???????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1828_ = b[1575:1568];
      256'b??????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1828_ = b[1583:1576];
      256'b?????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1828_ = b[1591:1584];
      256'b????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1828_ = b[1599:1592];
      256'b???????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1828_ = b[1607:1600];
      256'b??????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1828_ = b[1615:1608];
      256'b?????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1828_ = b[1623:1616];
      256'b????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1828_ = b[1631:1624];
      256'b???????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1828_ = b[1639:1632];
      256'b??????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1828_ = b[1647:1640];
      256'b?????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1828_ = b[1655:1648];
      256'b????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1828_ = b[1663:1656];
      256'b???????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1828_ = b[1671:1664];
      256'b??????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1828_ = b[1679:1672];
      256'b?????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1828_ = b[1687:1680];
      256'b????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1828_ = b[1695:1688];
      256'b???????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1828_ = b[1703:1696];
      256'b??????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1828_ = b[1711:1704];
      256'b?????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1828_ = b[1719:1712];
      256'b????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1828_ = b[1727:1720];
      256'b???????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1828_ = b[1735:1728];
      256'b??????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1828_ = b[1743:1736];
      256'b?????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1828_ = b[1751:1744];
      256'b????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1828_ = b[1759:1752];
      256'b???????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1828_ = b[1767:1760];
      256'b??????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1828_ = b[1775:1768];
      256'b?????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1828_ = b[1783:1776];
      256'b????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1828_ = b[1791:1784];
      256'b???????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1828_ = b[1799:1792];
      256'b??????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1828_ = b[1807:1800];
      256'b?????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1828_ = b[1815:1808];
      256'b????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1828_ = b[1823:1816];
      256'b???????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1828_ = b[1831:1824];
      256'b??????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1828_ = b[1839:1832];
      256'b?????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1828_ = b[1847:1840];
      256'b????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1828_ = b[1855:1848];
      256'b???????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1828_ = b[1863:1856];
      256'b??????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1828_ = b[1871:1864];
      256'b?????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1828_ = b[1879:1872];
      256'b????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1828_ = b[1887:1880];
      256'b???????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1828_ = b[1895:1888];
      256'b??????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1828_ = b[1903:1896];
      256'b?????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1828_ = b[1911:1904];
      256'b????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1828_ = b[1919:1912];
      256'b???????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1828_ = b[1927:1920];
      256'b??????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1828_ = b[1935:1928];
      256'b?????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1828_ = b[1943:1936];
      256'b????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1828_ = b[1951:1944];
      256'b???????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1828_ = b[1959:1952];
      256'b??????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1828_ = b[1967:1960];
      256'b?????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1828_ = b[1975:1968];
      256'b????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1828_ = b[1983:1976];
      256'b???????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1828_ = b[1991:1984];
      256'b??????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1828_ = b[1999:1992];
      256'b?????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1828_ = b[2007:2000];
      256'b????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1828_ = b[2015:2008];
      256'b???1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1828_ = b[2023:2016];
      256'b??1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1828_ = b[2031:2024];
      256'b?1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1828_ = b[2039:2032];
      256'b1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _1828_ = b[2047:2040];
      default:
        _1828_ = a;
    endcase
  endfunction
  assign _0771_ = _1828_(\S4_0.S_3.out , 2048'h637c777bf26b6fc53001672bfed7ab76ca82c97dfa5947f0add4a2af9ca472c0b7fd9326363ff7cc34a5e5f171d8311504c723c31896059a071280e2eb27b27509832c1a1b6e5aa0523bd6b329e32f8453d100ed20fcb15b6acbbe394a4c58cfd0efaafb434d338545f9027f503c9fa851a3408f929d38f5bcb6da2110fff3d2cd0c13ec5f974417c4a77e3d645d197360814fdc222a908846eeb814de5e0bdbe0323a0a4906245cc2d3ac629195e479e7c8376d8dd54ea96c56f4ea657aae08ba78252e1ca6b4c6e8dd741f4bbd8b8a703eb5664803f60e613557b986c11d9ee1f8981169d98e949b1e87e9ce5528df8ca1890dbfe6426841992d0fb054bb16, { _0953_, _0952_, _0951_, _0950_, _0949_, _0948_, _0947_, _0946_, _0945_, _0943_, _0942_, _0941_, _0940_, _0939_, _0938_, _0937_, _0936_, _0935_, _0934_, _0932_, _0931_, _0930_, _0929_, _0928_, _0927_, _0926_, _0925_, _0924_, _0923_, _0921_, _0920_, _0919_, _0918_, _0917_, _0916_, _0915_, _0914_, _0913_, _0912_, _0910_, _0909_, _0908_, _0907_, _0906_, _0905_, _0904_, _0903_, _0902_, _0901_, _0899_, _0898_, _0897_, _0896_, _0895_, _0894_, _0893_, _0892_, _0891_, _0890_, _0888_, _0887_, _0886_, _0885_, _0884_, _0883_, _0882_, _0881_, _0880_, _0879_, _0877_, _0876_, _0875_, _0874_, _0873_, _0872_, _0871_, _0870_, _0869_, _0868_, _0866_, _0865_, _0864_, _0863_, _0862_, _0861_, _0860_, _0859_, _0858_, _0857_, _0855_, _0854_, _0853_, _0852_, _0851_, _0850_, _0849_, _0848_, _0847_, _0846_, _0844_, _0843_, _0842_, _0841_, _0840_, _0839_, _0838_, _0837_, _0836_, _0835_, _0833_, _0832_, _0831_, _0830_, _0829_, _0828_, _0827_, _0826_, _0825_, _0824_, _0822_, _0821_, _0820_, _0819_, _0818_, _0817_, _0816_, _0815_, _0814_, _0813_, _0811_, _0810_, _0809_, _0808_, _0807_, _0806_, _0805_, _0804_, _0803_, _0802_, _0801_, _0800_, _0799_, _0798_, _0797_, _0796_, _0795_, _0794_, _0793_, _0792_, _0791_, _0790_, _0789_, _0788_, _0787_, _0786_, _0785_, _0784_, _0783_, _0782_, _0781_, _0780_, _0779_, _0778_, _0777_, _0776_, _0775_, _0774_, _0773_, _0772_, _1027_, _1026_, _1025_, _1024_, _1023_, _1022_, _1021_, _1020_, _1019_, _1018_, _1017_, _1016_, _1015_, _1014_, _1013_, _1012_, _1011_, _1010_, _1009_, _1008_, _1007_, _1006_, _1005_, _1004_, _1003_, _1002_, _1001_, _1000_, _0999_, _0998_, _0997_, _0996_, _0995_, _0994_, _0993_, _0992_, _0991_, _0990_, _0989_, _0988_, _0987_, _0986_, _0985_, _0984_, _0983_, _0982_, _0981_, _0980_, _0979_, _0978_, _0977_, _0976_, _0975_, _0974_, _0973_, _0972_, _0971_, _0970_, _0969_, _0968_, _0967_, _0966_, _0965_, _0964_, _0963_, _0962_, _0961_, _0960_, _0959_, _0958_, _0957_, _0956_, _0955_, _0954_, _0944_, _0933_, _0922_, _0911_, _0900_, _0889_, _0878_, _0867_, _0856_, _0845_, _0834_, _0823_, _0812_ });
  assign _0792_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'h94;
  assign _0793_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'h93;
  assign _0794_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'h92;
  assign _0795_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'h91;
  assign _0796_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'h90;
  assign _0797_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'h8f;
  assign _0798_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'h8e;
  assign _0799_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'h8d;
  assign _0800_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'h8c;
  assign _0801_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'h8b;
  assign _0802_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'h8a;
  assign _0803_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'h89;
  assign _0804_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'h88;
  assign _0805_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'h87;
  assign _0806_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'h86;
  assign _0807_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'h85;
  assign _0808_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'h84;
  assign _0809_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'h83;
  assign _0810_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'h82;
  assign _0811_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'h81;
  assign _0812_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hff;
  assign _0813_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'h80;
  assign _0814_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h7f;
  assign _0815_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h7e;
  assign _0816_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h7d;
  assign _0817_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h7c;
  assign _0818_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h7b;
  assign _0819_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h7a;
  assign _0820_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h79;
  assign _0821_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h78;
  assign _0822_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h77;
  assign _0823_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hfe;
  assign _0824_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h76;
  assign _0825_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h75;
  assign _0826_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h74;
  assign _0827_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h73;
  assign _0828_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h72;
  assign _0829_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h71;
  assign _0830_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h70;
  assign _0831_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h6f;
  assign _0832_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h6e;
  assign _0833_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h6d;
  assign _0834_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hfd;
  assign _0835_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h6c;
  assign _0836_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h6b;
  assign _0837_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h6a;
  assign _0838_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h69;
  assign _0839_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h68;
  assign _0840_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h67;
  assign _0841_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h66;
  assign _0842_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h65;
  assign _0843_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h64;
  assign _0844_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h63;
  assign _0845_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hfc;
  assign _0846_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h62;
  assign _0847_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h61;
  assign _0848_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h60;
  assign _0849_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h5f;
  assign _0850_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h5e;
  assign _0851_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h5d;
  assign _0852_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h5c;
  assign _0853_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h5b;
  assign _0854_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h5a;
  assign _0855_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h59;
  assign _0856_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hfb;
  assign _0857_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h58;
  assign _0858_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h57;
  assign _0859_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h56;
  assign _0860_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h55;
  assign _0861_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h54;
  assign _0862_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h53;
  assign _0863_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h52;
  assign _0864_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h51;
  assign _0865_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h50;
  assign _0866_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h4f;
  assign _0867_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hfa;
  assign _0868_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h4e;
  assign _0869_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h4d;
  assign _0870_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h4c;
  assign _0871_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h4b;
  assign _0872_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h4a;
  assign _0873_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h49;
  assign _0874_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h48;
  assign _0875_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h47;
  assign _0876_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h46;
  assign _0877_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h45;
  assign _0878_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hf9;
  assign _0879_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h44;
  assign _0880_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h43;
  assign _0881_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h42;
  assign _0882_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h41;
  assign _0883_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 7'h40;
  assign _0884_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 6'h3f;
  assign _0885_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 6'h3e;
  assign _0886_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 6'h3d;
  assign _0887_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 6'h3c;
  assign _0888_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 6'h3b;
  assign _0889_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hf8;
  assign _0890_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 6'h3a;
  assign _0891_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 6'h39;
  assign _0892_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 6'h38;
  assign _0893_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 6'h37;
  assign _0894_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 6'h36;
  assign _0895_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 6'h35;
  assign _0896_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 6'h34;
  assign _0897_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 6'h33;
  assign _0898_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 6'h32;
  assign _0899_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 6'h31;
  assign _0900_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hf7;
  assign _0901_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 6'h30;
  assign _0902_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 6'h2f;
  assign _0903_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 6'h2e;
  assign _0904_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 6'h2d;
  assign _0905_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 6'h2c;
  assign _0906_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 6'h2b;
  assign _0907_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 6'h2a;
  assign _0908_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 6'h29;
  assign _0909_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 6'h28;
  assign _0910_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 6'h27;
  assign _0911_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hf6;
  assign _0912_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 6'h26;
  assign _0913_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 6'h25;
  assign _0914_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 6'h24;
  assign _0915_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 6'h23;
  assign _0916_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 6'h22;
  assign _0917_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 6'h21;
  assign _0918_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 6'h20;
  assign _0919_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 5'h1f;
  assign _0920_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 5'h1e;
  assign _0921_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 5'h1d;
  assign _0922_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hf5;
  assign _0923_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 5'h1c;
  assign _0924_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 5'h1b;
  assign _0925_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 5'h1a;
  assign _0926_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 5'h19;
  assign _0927_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 5'h18;
  assign _0928_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 5'h17;
  assign _0929_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 5'h16;
  assign _0930_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 5'h15;
  assign _0931_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 5'h14;
  assign _0932_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 5'h13;
  assign _0933_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hf4;
  assign _0934_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 5'h12;
  assign _0935_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 5'h11;
  assign _0936_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 5'h10;
  assign _0937_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 4'hf;
  assign _0938_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 4'he;
  assign _0939_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 4'hd;
  assign _0940_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 4'hc;
  assign _0941_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 4'hb;
  assign _0942_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 4'ha;
  assign _0943_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 4'h9;
  assign _0944_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hf3;
  assign _0945_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 4'h8;
  assign _0946_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 3'h7;
  assign _0947_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 3'h6;
  assign _0948_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 3'h5;
  assign _0949_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 3'h4;
  assign _0950_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 2'h3;
  assign _0951_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 2'h2;
  assign _0952_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 1'h1;
  assign _0953_ = ! (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) in[31:24];
  assign _0954_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hf2;
  assign _0955_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hf1;
  assign _0956_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hf0;
  assign _0957_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hef;
  assign _0958_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hee;
  assign _0959_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hed;
  assign _0960_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hec;
  assign _0961_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'heb;
  assign _0962_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hea;
  assign _0963_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'he9;
  assign _0964_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'he8;
  assign _0965_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'he7;
  assign _0966_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'he6;
  assign _0967_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'he5;
  assign _0968_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'he4;
  assign _0969_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'he3;
  assign _0970_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'he2;
  assign _0971_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'he1;
  assign _0972_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'he0;
  assign _0973_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hdf;
  assign _0974_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hde;
  assign _0975_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hdd;
  assign _0976_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hdc;
  assign _0977_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hdb;
  assign _0978_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hda;
  assign _0979_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hd9;
  assign _0980_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hd8;
  assign _0981_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hd7;
  assign _0982_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hd6;
  assign _0983_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hd5;
  assign _0984_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hd4;
  assign _0985_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hd3;
  assign _0986_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hd2;
  assign _0987_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hd1;
  assign _0988_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hd0;
  assign _0989_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hcf;
  assign _0990_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hce;
  assign _0991_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hcd;
  assign _0992_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hcc;
  assign _0993_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hcb;
  assign _0994_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hca;
  assign _0995_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hc9;
  assign _0996_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hc8;
  assign _0997_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hc7;
  assign _0998_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hc6;
  assign _0999_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hc5;
  assign _1000_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hc4;
  assign _1001_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hc3;
  assign _1002_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hc2;
  assign _1003_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hc1;
  assign _1004_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hc0;
  assign _1005_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hbf;
  assign _1006_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hbe;
  assign _1007_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hbd;
  assign _1008_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hbc;
  assign _1009_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hbb;
  assign _1010_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hba;
  assign _1011_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hb9;
  assign _1012_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hb8;
  assign _1013_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hb7;
  assign _1014_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hb6;
  assign _1015_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hb5;
  assign _1016_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hb4;
  assign _1017_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hb3;
  assign _1018_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hb2;
  assign _1019_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hb1;
  assign _1020_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hb0;
  assign _1021_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'haf;
  assign _1022_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hae;
  assign _1023_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'had;
  assign _1024_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hac;
  assign _1025_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'hab;
  assign _1026_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'haa;
  assign _1027_ = in[31:24] == (* src = "expand_key_128.v:28|S4.v:26|S.v:12" *) 8'ha9;
  assign v0[31:24] = in[127:120] ^ (* src = "expand_key_128.v:20" *) rcon;
  assign v1 = { v0[31:24], in[119:96] } ^ (* src = "expand_key_128.v:21" *) in[95:64];
  assign v2 = v1 ^ (* src = "expand_key_128.v:22" *) in[63:32];
  assign v3 = v2 ^ (* src = "expand_key_128.v:23" *) in[31:0];
  assign k0b = k0a ^ (* src = "expand_key_128.v:31" *) { \S4_0.S_0.out , \S4_0.S_1.out , \S4_0.S_2.out , \S4_0.S_3.out  };
  assign k1b = k1a ^ (* src = "expand_key_128.v:32" *) { \S4_0.S_0.out , \S4_0.S_1.out , \S4_0.S_2.out , \S4_0.S_3.out  };
  assign k2b = k2a ^ (* src = "expand_key_128.v:33" *) { \S4_0.S_0.out , \S4_0.S_1.out , \S4_0.S_2.out , \S4_0.S_3.out  };
  assign k3b = k3a ^ (* src = "expand_key_128.v:34" *) { \S4_0.S_0.out , \S4_0.S_1.out , \S4_0.S_2.out , \S4_0.S_3.out  };
  assign \S4_0.S_0.clk  = clk;
  assign \S4_0.S_0.in  = in[23:16];
  assign \S4_0.S_1.clk  = clk;
  assign \S4_0.S_1.in  = in[15:8];
  assign \S4_0.S_2.clk  = clk;
  assign \S4_0.S_2.in  = in[7:0];
  assign \S4_0.S_3.clk  = clk;
  assign \S4_0.S_3.in  = in[31:24];
  assign \S4_0.clk  = clk;
  assign \S4_0.in  = { in[23:0], in[31:24] };
  assign \S4_0.out  = { \S4_0.S_0.out , \S4_0.S_1.out , \S4_0.S_2.out , \S4_0.S_3.out  };
  assign k0 = in[127:96];
  assign k1 = in[95:64];
  assign k2 = in[63:32];
  assign k3 = in[31:0];
  assign k4a = { \S4_0.S_0.out , \S4_0.S_1.out , \S4_0.S_2.out , \S4_0.S_3.out  };
  assign out_2 = { k0b, k1b, k2b, k3b };
  assign v0[23:0] = in[119:96];
endmodule
