module NV_BLKBOX_BUFFER(Y, A);
  (* src = "./vmod/vlibs/NV_BLKBOX_BUFFER.v:14" *)
  input A;
  (* src = "./vmod/vlibs/NV_BLKBOX_BUFFER.v:13" *)
  output Y;
  assign Y = A;
endmodule
