module accum(clk, data, rst, start, finish, sum, timer);
  input [0:0] clk ;
  input [2:0] data ;
  input [0:0] rst ;
  input [0:0] start ;
  output [0:0] finish ;
  output [2:0] sum ;
  output [2:0] timer ;
// moduleRegs
  reg [2:0] cnt ;
// regWithFunc
endmodule
