module read_eg_arb(req0, req1, req2, req3, req4, req5, req6, req7, req8, req9, wt0, wt1, wt2, wt3, wt4, wt5, wt6, wt7, wt8, wt9, clk, reset_, gnt0, gnt1, gnt2, gnt3, gnt4, gnt5, gnt6, gnt7, gnt8, gnt9);
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2498" *)
  wire [9:0] _000_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2498" *)
  wire [7:0] _001_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2001" *)
  wire [9:0] _002_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2001" *)
  wire [7:0] _003_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2001" *)
  wire [9:0] _004_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2001" *)
  wire [7:0] _005_;
  wire [8:0] _006_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2001" *)
  wire [7:0] _007_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2001" *)
  wire [9:0] _008_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2001" *)
  wire [7:0] _009_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2001" *)
  wire [9:0] _010_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2001" *)
  wire [7:0] _011_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2001" *)
  wire [9:0] _012_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2001" *)
  wire [7:0] _013_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2001" *)
  wire [9:0] _014_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2001" *)
  wire [7:0] _015_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2001" *)
  wire [9:0] _016_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2001" *)
  wire [7:0] _017_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2001" *)
  wire [9:0] _018_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2001" *)
  wire [7:0] _019_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2001" *)
  wire [9:0] _020_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2001" *)
  wire [7:0] _021_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2001" *)
  wire [9:0] _022_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2001" *)
  wire [7:0] _023_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2001" *)
  wire [9:0] _024_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2001" *)
  wire [7:0] _025_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2001" *)
  wire [9:0] _026_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2001" *)
  wire [7:0] _027_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2001" *)
  wire [9:0] _028_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2001" *)
  wire [7:0] _029_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2001" *)
  wire [9:0] _030_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2001" *)
  wire [7:0] _031_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2001" *)
  wire [9:0] _032_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2001" *)
  wire [7:0] _033_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2001" *)
  wire [9:0] _034_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2001" *)
  wire [7:0] _035_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2001" *)
  wire [9:0] _036_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2001" *)
  wire [7:0] _037_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2001" *)
  wire [9:0] _038_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2001" *)
  wire [7:0] _039_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2001" *)
  wire [9:0] _040_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2001" *)
  wire [7:0] _041_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2001" *)
  wire [9:0] _042_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2001" *)
  wire [7:0] _043_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2001" *)
  wire [9:0] _044_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2001" *)
  wire [7:0] _045_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2001" *)
  wire [7:0] _046_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2001" *)
  wire [9:0] _047_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2001" *)
  wire [7:0] _048_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2001" *)
  wire [9:0] _049_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2001" *)
  wire [7:0] _050_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2001" *)
  wire [9:0] _051_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2001" *)
  wire [7:0] _052_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2001" *)
  wire [9:0] _053_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2001" *)
  wire [7:0] _054_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2001" *)
  wire [9:0] _055_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2001" *)
  wire [7:0] _056_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2001" *)
  wire [9:0] _057_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2001" *)
  wire [7:0] _058_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2001" *)
  wire [9:0] _059_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2001" *)
  wire [7:0] _060_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2001" *)
  wire [9:0] _061_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2001" *)
  wire [7:0] _062_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2001" *)
  wire [9:0] _063_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2001" *)
  wire [7:0] _064_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2001" *)
  wire [9:0] _065_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2001" *)
  wire [7:0] _066_;
  wire [1:0] _067_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2001" *)
  wire [7:0] _068_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2001" *)
  wire [9:0] _069_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2001" *)
  wire [7:0] _070_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2001" *)
  wire [9:0] _071_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2001" *)
  wire [7:0] _072_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2001" *)
  wire [9:0] _073_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2001" *)
  wire [7:0] _074_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2001" *)
  wire [9:0] _075_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2001" *)
  wire [7:0] _076_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2001" *)
  wire [9:0] _077_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2001" *)
  wire [7:0] _078_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2001" *)
  wire [9:0] _079_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2001" *)
  wire [7:0] _080_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2001" *)
  wire [9:0] _081_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2001" *)
  wire [7:0] _082_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2001" *)
  wire [9:0] _083_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2001" *)
  wire [7:0] _084_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2001" *)
  wire [9:0] _085_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2001" *)
  wire [7:0] _086_;
  wire [2:0] _087_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2001" *)
  wire [7:0] _088_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2001" *)
  wire [9:0] _089_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2001" *)
  wire [7:0] _090_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2001" *)
  wire [9:0] _091_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2001" *)
  wire [7:0] _092_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2001" *)
  wire [9:0] _093_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2001" *)
  wire [7:0] _094_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2001" *)
  wire [9:0] _095_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2001" *)
  wire [7:0] _096_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2001" *)
  wire [9:0] _097_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2001" *)
  wire [7:0] _098_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2001" *)
  wire [9:0] _099_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2001" *)
  wire [7:0] _100_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2001" *)
  wire [9:0] _101_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2001" *)
  wire [7:0] _102_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2001" *)
  wire [9:0] _103_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2001" *)
  wire [7:0] _104_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2001" *)
  wire [9:0] _105_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2001" *)
  wire [7:0] _106_;
  wire [3:0] _107_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2001" *)
  wire [7:0] _108_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2001" *)
  wire [9:0] _109_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2001" *)
  wire [7:0] _110_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2001" *)
  wire [9:0] _111_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2001" *)
  wire [7:0] _112_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2001" *)
  wire [9:0] _113_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2001" *)
  wire [7:0] _114_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2001" *)
  wire [9:0] _115_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2001" *)
  wire [7:0] _116_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2001" *)
  wire [9:0] _117_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2001" *)
  wire [7:0] _118_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2001" *)
  wire [9:0] _119_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2001" *)
  wire [7:0] _120_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2001" *)
  wire [9:0] _121_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2001" *)
  wire [7:0] _122_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2001" *)
  wire [9:0] _123_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2001" *)
  wire [7:0] _124_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2001" *)
  wire [9:0] _125_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2001" *)
  wire [7:0] _126_;
  wire [4:0] _127_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2001" *)
  wire [7:0] _128_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2001" *)
  wire [9:0] _129_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2001" *)
  wire [7:0] _130_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2001" *)
  wire [9:0] _131_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2001" *)
  wire [7:0] _132_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2001" *)
  wire [9:0] _133_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2001" *)
  wire [7:0] _134_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2001" *)
  wire [9:0] _135_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2001" *)
  wire [7:0] _136_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2001" *)
  wire [9:0] _137_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2001" *)
  wire [7:0] _138_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2001" *)
  wire [9:0] _139_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2001" *)
  wire [7:0] _140_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2001" *)
  wire [9:0] _141_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2001" *)
  wire [7:0] _142_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2001" *)
  wire [9:0] _143_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2001" *)
  wire [7:0] _144_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2001" *)
  wire [9:0] _145_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2001" *)
  wire [7:0] _146_;
  wire [5:0] _147_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2001" *)
  wire [7:0] _148_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2001" *)
  wire [9:0] _149_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2001" *)
  wire [7:0] _150_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2001" *)
  wire [9:0] _151_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2001" *)
  wire [7:0] _152_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2001" *)
  wire [9:0] _153_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2001" *)
  wire [7:0] _154_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2001" *)
  wire [9:0] _155_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2001" *)
  wire [7:0] _156_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2001" *)
  wire [9:0] _157_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2001" *)
  wire [7:0] _158_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2001" *)
  wire [9:0] _159_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2001" *)
  wire [7:0] _160_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2001" *)
  wire [9:0] _161_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2001" *)
  wire [7:0] _162_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2001" *)
  wire [9:0] _163_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2001" *)
  wire [7:0] _164_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2001" *)
  wire [9:0] _165_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2001" *)
  wire [7:0] _166_;
  wire [6:0] _167_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2001" *)
  wire [7:0] _168_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2001" *)
  wire [9:0] _169_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2001" *)
  wire [7:0] _170_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2001" *)
  wire [9:0] _171_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2001" *)
  wire [7:0] _172_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2001" *)
  wire [9:0] _173_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2001" *)
  wire [7:0] _174_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2001" *)
  wire [9:0] _175_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2001" *)
  wire [7:0] _176_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2001" *)
  wire [9:0] _177_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2001" *)
  wire [7:0] _178_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2001" *)
  wire [9:0] _179_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2001" *)
  wire [7:0] _180_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2001" *)
  wire [9:0] _181_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2001" *)
  wire [7:0] _182_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2001" *)
  wire [9:0] _183_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2001" *)
  wire [7:0] _184_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2001" *)
  wire [9:0] _185_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2001" *)
  wire [7:0] _186_;
  wire [7:0] _187_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2001" *)
  wire [7:0] _188_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2001" *)
  wire [9:0] _189_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2001" *)
  wire [7:0] _190_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2001" *)
  wire [9:0] _191_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2001" *)
  wire [7:0] _192_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2001" *)
  wire [9:0] _193_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2001" *)
  wire [7:0] _194_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2001" *)
  wire [9:0] _195_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2001" *)
  wire [7:0] _196_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2001" *)
  wire [9:0] _197_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2001" *)
  wire [7:0] _198_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2001" *)
  wire [9:0] _199_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2001" *)
  wire [7:0] _200_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2001" *)
  wire [9:0] _201_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2001" *)
  wire [7:0] _202_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2018" *)
  wire [9:0] _203_;
  wire _204_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2018" *)
  wire _205_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2018" *)
  wire _206_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2503" *)
  wire _207_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2018" *)
  wire _208_;
  wire _209_;
  wire _210_;
  wire _211_;
  wire _212_;
  wire _213_;
  wire _214_;
  wire _215_;
  wire _216_;
  wire _217_;
  wire _218_;
  wire _219_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:1959" *)
  wire _220_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:1960" *)
  wire _221_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:1961" *)
  wire _222_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:1962" *)
  wire _223_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:1963" *)
  wire _224_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:1964" *)
  wire _225_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:1965" *)
  wire _226_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:1966" *)
  wire _227_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:1967" *)
  wire _228_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:1968" *)
  wire _229_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2018" *)
  wire _230_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2491" *)
  wire [7:0] _231_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:1928" *)
  input clk;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:1942" *)
  wire [9:0] gnt;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:1930" *)
  output gnt0;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:1931" *)
  output gnt1;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:1932" *)
  output gnt2;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:1933" *)
  output gnt3;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:1934" *)
  output gnt4;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:1935" *)
  output gnt5;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:1936" *)
  output gnt6;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:1937" *)
  output gnt7;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:1938" *)
  output gnt8;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:1939" *)
  output gnt9;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:1943" *)
  wire [9:0] gnt_pre;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:1947" *)
  wire [7:0] new_wt_left0;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:1948" *)
  wire [7:0] new_wt_left1;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:1949" *)
  wire [7:0] new_wt_left2;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:1950" *)
  wire [7:0] new_wt_left3;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:1951" *)
  wire [7:0] new_wt_left4;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:1952" *)
  wire [7:0] new_wt_left5;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:1953" *)
  wire [7:0] new_wt_left6;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:1954" *)
  wire [7:0] new_wt_left7;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:1955" *)
  wire [7:0] new_wt_left8;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:1956" *)
  wire [7:0] new_wt_left9;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:1957" *)
  wire [9:0] req;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:1908" *)
  input req0;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:1909" *)
  input req1;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:1910" *)
  input req2;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:1911" *)
  input req3;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:1912" *)
  input req4;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:1913" *)
  input req5;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:1914" *)
  input req6;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:1915" *)
  input req7;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:1916" *)
  input req8;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:1917" *)
  input req9;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:1929" *)
  input reset_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:1944" *)
  reg [9:0] wrr_gnt;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:1918" *)
  input [7:0] wt0;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:1919" *)
  input [7:0] wt1;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:1920" *)
  input [7:0] wt2;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:1921" *)
  input [7:0] wt3;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:1922" *)
  input [7:0] wt4;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:1923" *)
  input [7:0] wt5;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:1924" *)
  input [7:0] wt6;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:1925" *)
  input [7:0] wt7;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:1926" *)
  input [7:0] wt8;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:1927" *)
  input [7:0] wt9;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:1945" *)
  reg [7:0] wt_left;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:1946" *)
  wire [7:0] wt_left_nxt;
  assign req[9] = req9 & (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:1959" *) _220_;
  assign req[8] = req8 & (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:1960" *) _221_;
  assign req[7] = req7 & (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:1961" *) _222_;
  assign req[6] = req6 & (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:1962" *) _223_;
  assign req[5] = req5 & (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:1963" *) _224_;
  assign req[4] = req4 & (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:1964" *) _225_;
  assign req[3] = req3 & (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:1965" *) _226_;
  assign req[2] = req2 & (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:1966" *) _227_;
  assign req[1] = req1 & (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:1967" *) _228_;
  assign req[0] = req0 & (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:1968" *) _229_;
  assign _203_ = req & (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2018" *) wrr_gnt;
  assign _204_ = | { _209_, _219_ };
  assign _205_ = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2018" *) wt_left;
  assign _206_ = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2018" *) _230_;
  assign _207_ = | (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2503" *) req;
  assign _208_ = _205_ | (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2018" *) _206_;
  always @(posedge clk or negedge reset_)
    if (!reset_)
      wrr_gnt <= 10'b0000000000;
    else
      wrr_gnt <= _000_;
  always @(posedge clk or negedge reset_)
    if (!reset_)
      wt_left <= 8'b00000000;
    else
      wt_left <= _001_;
  assign _001_ = _207_ ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2503" *) wt_left_nxt : wt_left;
  assign _000_ = _207_ ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2503" *) gnt : wrr_gnt;
  assign _209_ = wrr_gnt == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2440|./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2019" *) 10'b1000000000;
  assign _024_ = req[8] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2473" *) 10'b0100000000 : _026_;
  assign _023_ = req[7] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2469" *) new_wt_left7 : _025_;
  assign _019_ = req[5] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2461" *) new_wt_left5 : _021_;
  assign _017_ = req[4] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2457" *) new_wt_left4 : _019_;
  assign _016_ = req[4] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2457" *) 10'b0000010000 : _018_;
  assign _015_ = req[3] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2453" *) new_wt_left3 : _017_;
  assign _014_ = req[3] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2453" *) 10'b0000001000 : _016_;
  assign _013_ = req[2] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2449" *) new_wt_left2 : _015_;
  assign _012_ = req[2] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2449" *) 10'b0000000100 : _014_;
  assign _011_ = req[1] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2445" *) new_wt_left1 : _013_;
  assign _010_ = req[1] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2445" *) 10'b0000000010 : _012_;
  assign _009_ = req[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2441" *) new_wt_left0 : _011_;
  assign _008_ = req[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2441" *) 10'b0000000001 : _010_;
  assign _007_ = req[8] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2435" *) new_wt_left8 : wt_left;
  assign _210_ = wrr_gnt == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2398|./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2019" *) 9'b100000000;
  assign _006_ = req[8] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2435" *) 9'b100000000 : 9'b000000000;
  assign _005_ = req[7] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2431" *) new_wt_left7 : _007_;
  assign _004_ = req[7] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2431" *) 10'b0010000000 : { 1'b0, _006_ };
  assign _003_ = req[6] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2427" *) new_wt_left6 : _005_;
  assign _002_ = req[6] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2427" *) 10'b0001000000 : _004_;
  assign _202_ = req[5] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2423" *) new_wt_left5 : _003_;
  assign _201_ = req[5] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2423" *) 10'b0000100000 : _002_;
  assign _200_ = req[4] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2419" *) new_wt_left4 : _202_;
  assign _199_ = req[4] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2419" *) 10'b0000010000 : _201_;
  assign _198_ = req[3] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2415" *) new_wt_left3 : _200_;
  assign _197_ = req[3] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2415" *) 10'b0000001000 : _199_;
  assign _196_ = req[2] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2411" *) new_wt_left2 : _198_;
  assign _195_ = req[2] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2411" *) 10'b0000000100 : _197_;
  assign _194_ = req[1] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2407" *) new_wt_left1 : _196_;
  assign _193_ = req[1] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2407" *) 10'b0000000010 : _195_;
  assign _192_ = req[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2403" *) new_wt_left0 : _194_;
  assign _191_ = req[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2403" *) 10'b0000000001 : _193_;
  assign _190_ = req[9] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2399" *) new_wt_left9 : _192_;
  assign _189_ = req[9] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2399" *) 10'b1000000000 : _191_;
  assign _188_ = req[7] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2393" *) new_wt_left7 : wt_left;
  assign _211_ = wrr_gnt == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2356|./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2019" *) 8'b10000000;
  assign _187_ = req[7] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2393" *) 8'b10000000 : 8'b00000000;
  assign _186_ = req[6] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2389" *) new_wt_left6 : _188_;
  assign _185_ = req[6] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2389" *) 10'b0001000000 : { 2'b00, _187_ };
  assign _184_ = req[5] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2385" *) new_wt_left5 : _186_;
  assign _183_ = req[5] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2385" *) 10'b0000100000 : _185_;
  assign _182_ = req[4] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2381" *) new_wt_left4 : _184_;
  assign _181_ = req[4] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2381" *) 10'b0000010000 : _183_;
  assign _180_ = req[3] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2377" *) new_wt_left3 : _182_;
  assign _179_ = req[3] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2377" *) 10'b0000001000 : _181_;
  assign _178_ = req[2] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2373" *) new_wt_left2 : _180_;
  assign _177_ = req[2] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2373" *) 10'b0000000100 : _179_;
  assign _176_ = req[1] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2369" *) new_wt_left1 : _178_;
  assign _175_ = req[1] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2369" *) 10'b0000000010 : _177_;
  assign _174_ = req[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2365" *) new_wt_left0 : _176_;
  assign _173_ = req[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2365" *) 10'b0000000001 : _175_;
  assign _172_ = req[9] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2361" *) new_wt_left9 : _174_;
  assign _171_ = req[9] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2361" *) 10'b1000000000 : _173_;
  assign _170_ = req[8] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2357" *) new_wt_left8 : _172_;
  assign _169_ = req[8] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2357" *) 10'b0100000000 : _171_;
  assign _168_ = req[6] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2351" *) new_wt_left6 : wt_left;
  assign _212_ = wrr_gnt == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2314|./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2019" *) 7'b1000000;
  assign _167_ = req[6] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2351" *) 7'b1000000 : 7'b0000000;
  assign _166_ = req[5] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2347" *) new_wt_left5 : _168_;
  assign _165_ = req[5] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2347" *) 10'b0000100000 : { 3'b000, _167_ };
  assign _164_ = req[4] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2343" *) new_wt_left4 : _166_;
  assign _163_ = req[4] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2343" *) 10'b0000010000 : _165_;
  assign _162_ = req[3] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2339" *) new_wt_left3 : _164_;
  assign _161_ = req[3] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2339" *) 10'b0000001000 : _163_;
  assign _160_ = req[2] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2335" *) new_wt_left2 : _162_;
  assign _159_ = req[2] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2335" *) 10'b0000000100 : _161_;
  assign _158_ = req[1] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2331" *) new_wt_left1 : _160_;
  assign _157_ = req[1] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2331" *) 10'b0000000010 : _159_;
  assign _156_ = req[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2327" *) new_wt_left0 : _158_;
  assign _155_ = req[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2327" *) 10'b0000000001 : _157_;
  assign _154_ = req[9] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2323" *) new_wt_left9 : _156_;
  assign _153_ = req[9] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2323" *) 10'b1000000000 : _155_;
  assign _152_ = req[8] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2319" *) new_wt_left8 : _154_;
  assign _151_ = req[8] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2319" *) 10'b0100000000 : _153_;
  assign _150_ = req[7] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2315" *) new_wt_left7 : _152_;
  assign _149_ = req[7] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2315" *) 10'b0010000000 : _151_;
  assign _148_ = req[5] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2309" *) new_wt_left5 : wt_left;
  assign _213_ = wrr_gnt == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2272|./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2019" *) 6'b100000;
  assign _147_ = req[5] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2309" *) 6'b100000 : 6'b000000;
  assign _146_ = req[4] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2305" *) new_wt_left4 : _148_;
  assign _145_ = req[4] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2305" *) 10'b0000010000 : { 4'b0000, _147_ };
  assign _144_ = req[3] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2301" *) new_wt_left3 : _146_;
  assign _143_ = req[3] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2301" *) 10'b0000001000 : _145_;
  assign _142_ = req[2] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2297" *) new_wt_left2 : _144_;
  assign _141_ = req[2] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2297" *) 10'b0000000100 : _143_;
  assign _140_ = req[1] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2293" *) new_wt_left1 : _142_;
  assign _139_ = req[1] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2293" *) 10'b0000000010 : _141_;
  assign _138_ = req[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2289" *) new_wt_left0 : _140_;
  assign _137_ = req[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2289" *) 10'b0000000001 : _139_;
  assign _136_ = req[9] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2285" *) new_wt_left9 : _138_;
  assign _135_ = req[9] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2285" *) 10'b1000000000 : _137_;
  assign _134_ = req[8] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2281" *) new_wt_left8 : _136_;
  assign _133_ = req[8] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2281" *) 10'b0100000000 : _135_;
  assign _132_ = req[7] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2277" *) new_wt_left7 : _134_;
  assign _131_ = req[7] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2277" *) 10'b0010000000 : _133_;
  assign _130_ = req[6] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2273" *) new_wt_left6 : _132_;
  assign _129_ = req[6] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2273" *) 10'b0001000000 : _131_;
  assign _128_ = req[4] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2267" *) new_wt_left4 : wt_left;
  assign _214_ = wrr_gnt == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2230|./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2019" *) 5'b10000;
  assign _127_ = req[4] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2267" *) 5'b10000 : 5'b00000;
  assign _126_ = req[3] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2263" *) new_wt_left3 : _128_;
  assign _125_ = req[3] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2263" *) 10'b0000001000 : { 5'b00000, _127_ };
  assign _124_ = req[2] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2259" *) new_wt_left2 : _126_;
  assign _123_ = req[2] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2259" *) 10'b0000000100 : _125_;
  assign _122_ = req[1] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2255" *) new_wt_left1 : _124_;
  assign _121_ = req[1] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2255" *) 10'b0000000010 : _123_;
  assign _120_ = req[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2251" *) new_wt_left0 : _122_;
  assign _119_ = req[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2251" *) 10'b0000000001 : _121_;
  assign _118_ = req[9] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2247" *) new_wt_left9 : _120_;
  assign _117_ = req[9] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2247" *) 10'b1000000000 : _119_;
  assign _116_ = req[8] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2243" *) new_wt_left8 : _118_;
  assign _115_ = req[8] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2243" *) 10'b0100000000 : _117_;
  assign _114_ = req[7] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2239" *) new_wt_left7 : _116_;
  assign _113_ = req[7] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2239" *) 10'b0010000000 : _115_;
  assign _112_ = req[6] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2235" *) new_wt_left6 : _114_;
  assign _111_ = req[6] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2235" *) 10'b0001000000 : _113_;
  assign _110_ = req[5] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2231" *) new_wt_left5 : _112_;
  assign _109_ = req[5] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2231" *) 10'b0000100000 : _111_;
  assign _108_ = req[3] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2225" *) new_wt_left3 : wt_left;
  assign _215_ = wrr_gnt == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2188|./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2019" *) 4'b1000;
  assign _107_ = req[3] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2225" *) 4'b1000 : 4'b0000;
  assign _106_ = req[2] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2221" *) new_wt_left2 : _108_;
  assign _105_ = req[2] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2221" *) 10'b0000000100 : { 6'b000000, _107_ };
  assign _104_ = req[1] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2217" *) new_wt_left1 : _106_;
  assign _103_ = req[1] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2217" *) 10'b0000000010 : _105_;
  assign _102_ = req[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2213" *) new_wt_left0 : _104_;
  assign _101_ = req[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2213" *) 10'b0000000001 : _103_;
  assign _100_ = req[9] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2209" *) new_wt_left9 : _102_;
  assign _099_ = req[9] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2209" *) 10'b1000000000 : _101_;
  assign _098_ = req[8] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2205" *) new_wt_left8 : _100_;
  assign _097_ = req[8] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2205" *) 10'b0100000000 : _099_;
  assign _096_ = req[7] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2201" *) new_wt_left7 : _098_;
  assign _095_ = req[7] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2201" *) 10'b0010000000 : _097_;
  assign _094_ = req[6] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2197" *) new_wt_left6 : _096_;
  assign _093_ = req[6] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2197" *) 10'b0001000000 : _095_;
  assign _092_ = req[5] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2193" *) new_wt_left5 : _094_;
  assign _091_ = req[5] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2193" *) 10'b0000100000 : _093_;
  assign _090_ = req[4] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2189" *) new_wt_left4 : _092_;
  assign _089_ = req[4] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2189" *) 10'b0000010000 : _091_;
  assign _088_ = req[2] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2183" *) new_wt_left2 : wt_left;
  assign _216_ = wrr_gnt == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2146|./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2019" *) 3'b100;
  assign _087_ = req[2] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2183" *) 3'b100 : 3'b000;
  assign _086_ = req[1] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2179" *) new_wt_left1 : _088_;
  assign _085_ = req[1] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2179" *) 10'b0000000010 : { 7'b0000000, _087_ };
  assign _084_ = req[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2175" *) new_wt_left0 : _086_;
  assign _083_ = req[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2175" *) 10'b0000000001 : _085_;
  assign _082_ = req[9] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2171" *) new_wt_left9 : _084_;
  assign _081_ = req[9] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2171" *) 10'b1000000000 : _083_;
  assign _080_ = req[8] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2167" *) new_wt_left8 : _082_;
  assign _079_ = req[8] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2167" *) 10'b0100000000 : _081_;
  assign _078_ = req[7] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2163" *) new_wt_left7 : _080_;
  assign _077_ = req[7] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2163" *) 10'b0010000000 : _079_;
  assign _076_ = req[6] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2159" *) new_wt_left6 : _078_;
  assign _075_ = req[6] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2159" *) 10'b0001000000 : _077_;
  assign _074_ = req[5] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2155" *) new_wt_left5 : _076_;
  assign _073_ = req[5] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2155" *) 10'b0000100000 : _075_;
  assign _072_ = req[4] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2151" *) new_wt_left4 : _074_;
  assign _071_ = req[4] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2151" *) 10'b0000010000 : _073_;
  assign _070_ = req[3] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2147" *) new_wt_left3 : _072_;
  assign _069_ = req[3] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2147" *) 10'b0000001000 : _071_;
  assign _068_ = req[1] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2141" *) new_wt_left1 : wt_left;
  assign _217_ = wrr_gnt == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2104|./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2019" *) 2'b10;
  assign _067_ = req[1] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2141" *) 2'b10 : 2'b00;
  assign _066_ = req[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2137" *) new_wt_left0 : _068_;
  assign _065_ = req[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2137" *) 10'b0000000001 : { 8'b00000000, _067_ };
  assign _064_ = req[9] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2133" *) new_wt_left9 : _066_;
  assign _063_ = req[9] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2133" *) 10'b1000000000 : _065_;
  assign _060_ = req[8] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2129" *) new_wt_left8 : _064_;
  assign _059_ = req[8] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2129" *) 10'b0100000000 : _063_;
  assign _058_ = req[7] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2125" *) new_wt_left7 : _060_;
  assign _057_ = req[7] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2125" *) 10'b0010000000 : _059_;
  assign _056_ = req[6] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2121" *) new_wt_left6 : _058_;
  assign _055_ = req[6] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2121" *) 10'b0001000000 : _057_;
  assign _054_ = req[5] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2117" *) new_wt_left5 : _056_;
  assign _053_ = req[5] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2117" *) 10'b0000100000 : _055_;
  assign _052_ = req[4] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2113" *) new_wt_left4 : _054_;
  assign _051_ = req[4] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2113" *) 10'b0000010000 : _053_;
  assign _050_ = req[3] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2109" *) new_wt_left3 : _052_;
  assign _049_ = req[3] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2109" *) 10'b0000001000 : _051_;
  assign _048_ = req[2] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2105" *) new_wt_left2 : _050_;
  assign _047_ = req[2] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2105" *) 10'b0000000100 : _049_;
  assign _046_ = req[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2099" *) new_wt_left0 : wt_left;
  assign _218_ = wrr_gnt == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2062|./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2019" *) 1'b1;
  assign _045_ = req[9] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2095" *) new_wt_left9 : _046_;
  assign _044_ = req[9] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2095" *) 10'b1000000000 : { 9'b000000000, req[0] };
  assign _043_ = req[8] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2091" *) new_wt_left8 : _045_;
  assign _042_ = req[8] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2091" *) 10'b0100000000 : _044_;
  assign _041_ = req[7] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2087" *) new_wt_left7 : _043_;
  assign _040_ = req[7] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2087" *) 10'b0010000000 : _042_;
  assign _039_ = req[6] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2083" *) new_wt_left6 : _041_;
  assign _038_ = req[6] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2083" *) 10'b0001000000 : _040_;
  assign _037_ = req[5] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2079" *) new_wt_left5 : _039_;
  assign _036_ = req[5] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2079" *) 10'b0000100000 : _038_;
  assign _035_ = req[4] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2075" *) new_wt_left4 : _037_;
  assign _034_ = req[4] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2075" *) 10'b0000010000 : _036_;
  assign _033_ = req[3] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2071" *) new_wt_left3 : _035_;
  assign _032_ = req[3] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2071" *) 10'b0000001000 : _034_;
  assign _031_ = req[2] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2067" *) new_wt_left2 : _033_;
  assign _030_ = req[2] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2067" *) 10'b0000000100 : _032_;
  assign _029_ = req[1] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2063" *) new_wt_left1 : _031_;
  assign _028_ = req[1] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2063" *) 10'b0000000010 : _030_;
  assign _027_ = req[9] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2057" *) new_wt_left9 : wt_left;
  assign _219_ = ! (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2020|./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2019" *) wrr_gnt;
  assign _026_ = req[9] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2057" *) 10'b1000000000 : 10'b0000000000;
  assign _025_ = req[8] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2053" *) new_wt_left8 : _027_;
  assign _022_ = req[7] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2049" *) 10'b0010000000 : _024_;
  assign _021_ = req[6] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2045" *) new_wt_left6 : _023_;
  assign _020_ = req[6] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2045" *) 10'b0001000000 : _022_;
  assign _018_ = req[5] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2041" *) 10'b0000100000 : _020_;
  function [7:0] _462_;
    input [7:0] a;
    input [79:0] b;
    input [9:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2440|./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2019" *)
    (* parallel_case *)
    casez (s)
      10'b?????????1:
        _462_ = b[7:0];
      10'b????????1?:
        _462_ = b[15:8];
      10'b???????1??:
        _462_ = b[23:16];
      10'b??????1???:
        _462_ = b[31:24];
      10'b?????1????:
        _462_ = b[39:32];
      10'b????1?????:
        _462_ = b[47:40];
      10'b???1??????:
        _462_ = b[55:48];
      10'b??1???????:
        _462_ = b[63:56];
      10'b?1????????:
        _462_ = b[71:64];
      10'b1?????????:
        _462_ = b[79:72];
      default:
        _462_ = a;
    endcase
  endfunction
  assign _062_ = _462_(8'b00000000, { _029_, _048_, _070_, _090_, _110_, _130_, _150_, _170_, _190_, _009_ }, { _218_, _217_, _216_, _215_, _214_, _213_, _212_, _211_, _210_, _204_ });
  function [9:0] _463_;
    input [9:0] a;
    input [99:0] b;
    input [9:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2440|./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2019" *)
    (* parallel_case *)
    casez (s)
      10'b?????????1:
        _463_ = b[9:0];
      10'b????????1?:
        _463_ = b[19:10];
      10'b???????1??:
        _463_ = b[29:20];
      10'b??????1???:
        _463_ = b[39:30];
      10'b?????1????:
        _463_ = b[49:40];
      10'b????1?????:
        _463_ = b[59:50];
      10'b???1??????:
        _463_ = b[69:60];
      10'b??1???????:
        _463_ = b[79:70];
      10'b?1????????:
        _463_ = b[89:80];
      10'b1?????????:
        _463_ = b[99:90];
      default:
        _463_ = a;
    endcase
  endfunction
  assign _061_ = _463_(10'b0000000000, { _028_, _047_, _069_, _089_, _109_, _129_, _149_, _169_, _189_, _008_ }, { _218_, _217_, _216_, _215_, _214_, _213_, _212_, _211_, _210_, _204_ });
  assign wt_left_nxt = _208_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2018" *) _062_ : _231_;
  assign gnt = _208_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2018" *) _061_ : wrr_gnt;
  assign _220_ = | (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:1959" *) { wt9[0], wt9[1], wt9[2], wt9[3], wt9[4], wt9[5], wt9[6], wt9[7] };
  assign _221_ = | (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:1960" *) { wt8[0], wt8[1], wt8[2], wt8[3], wt8[4], wt8[5], wt8[6], wt8[7] };
  assign _222_ = | (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:1961" *) { wt7[0], wt7[1], wt7[2], wt7[3], wt7[4], wt7[5], wt7[6], wt7[7] };
  assign _223_ = | (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:1962" *) { wt6[0], wt6[1], wt6[2], wt6[3], wt6[4], wt6[5], wt6[6], wt6[7] };
  assign _224_ = | (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:1963" *) { wt5[0], wt5[1], wt5[2], wt5[3], wt5[4], wt5[5], wt5[6], wt5[7] };
  assign _225_ = | (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:1964" *) { wt4[0], wt4[1], wt4[2], wt4[3], wt4[4], wt4[5], wt4[6], wt4[7] };
  assign _226_ = | (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:1965" *) { wt3[0], wt3[1], wt3[2], wt3[3], wt3[4], wt3[5], wt3[6], wt3[7] };
  assign _227_ = | (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:1966" *) { wt2[0], wt2[1], wt2[2], wt2[3], wt2[4], wt2[5], wt2[6], wt2[7] };
  assign _228_ = | (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:1967" *) { wt1[0], wt1[1], wt1[2], wt1[3], wt1[4], wt1[5], wt1[6], wt1[7] };
  assign _229_ = | (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:1968" *) { wt0[0], wt0[1], wt0[2], wt0[3], wt0[4], wt0[5], wt0[6], wt0[7] };
  assign _230_ = | (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2018" *) { _203_[0], _203_[1], _203_[2], _203_[3], _203_[4], _203_[5], _203_[6], _203_[7], _203_[8], _203_[9] };
  assign new_wt_left0 = wt0 - (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:1991" *) 1'b1;
  assign new_wt_left1 = wt1 - (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:1992" *) 1'b1;
  assign new_wt_left2 = wt2 - (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:1993" *) 1'b1;
  assign new_wt_left3 = wt3 - (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:1994" *) 1'b1;
  assign new_wt_left4 = wt4 - (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:1995" *) 1'b1;
  assign new_wt_left5 = wt5 - (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:1996" *) 1'b1;
  assign new_wt_left6 = wt6 - (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:1997" *) 1'b1;
  assign new_wt_left7 = wt7 - (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:1998" *) 1'b1;
  assign new_wt_left8 = wt8 - (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:1999" *) 1'b1;
  assign new_wt_left9 = wt9 - (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2000" *) 1'b1;
  assign _231_ = wt_left - (* src = "./vmod/nvdla/nocif/NV_NVDLA_XXIF_libs.v:2491" *) 1'b1;
  assign gnt0 = gnt[0];
  assign gnt1 = gnt[1];
  assign gnt2 = gnt[2];
  assign gnt3 = gnt[3];
  assign gnt4 = gnt[4];
  assign gnt5 = gnt[5];
  assign gnt6 = gnt[6];
  assign gnt7 = gnt[7];
  assign gnt8 = gnt[8];
  assign gnt9 = gnt[9];
  assign gnt_pre = gnt;
endmodule
