module OR2D1(A1, A2, Z);
  (* src = "./vmod/vlibs/OR2D1.v:14" *)
  input A1;
  (* src = "./vmod/vlibs/OR2D1.v:15" *)
  input A2;
  (* src = "./vmod/vlibs/OR2D1.v:16" *)
  output Z;
  assign Z = A1 | (* src = "./vmod/vlibs/OR2D1.v:17" *) A2;
endmodule
