module \$paramod\SDP_Y_CORE_mgc_in_wire_v1\rscid=17\width=32 (d, z);
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:376" *)
  output [31:0] d;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:377" *)
  input [31:0] z;
  assign d = z;
endmodule
