module FP32_ADD_leading_sign_49_0(mantissa, rtn);
  (* src = "./vmod/vlibs/HLS_fp32_add.v:257" *)
  wire _000_;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:271" *)
  wire _001_;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:271" *)
  wire _002_;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:284" *)
  wire _003_;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:290" *)
  wire _004_;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:291" *)
  wire _005_;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:291" *)
  wire _006_;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:293" *)
  wire _007_;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:294" *)
  wire _008_;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:295" *)
  wire _009_;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:295" *)
  wire _010_;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:295" *)
  wire _011_;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:296" *)
  wire _012_;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:299" *)
  wire _013_;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:300" *)
  wire _014_;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:300" *)
  wire _015_;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:301" *)
  wire _016_;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:302" *)
  wire _017_;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:303" *)
  wire _018_;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:304" *)
  wire _019_;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:304" *)
  wire _020_;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:304" *)
  wire _021_;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:304" *)
  wire _022_;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:306" *)
  wire _023_;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:307" *)
  wire _024_;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:307" *)
  wire _025_;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:307" *)
  wire _026_;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:308" *)
  wire _027_;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:311" *)
  wire _028_;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:311" *)
  wire _029_;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:312" *)
  wire _030_;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:312" *)
  wire _031_;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:312" *)
  wire _032_;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:313" *)
  wire _033_;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:314" *)
  wire _034_;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:314" *)
  wire _035_;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:315" *)
  wire _036_;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:315" *)
  wire _037_;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:315" *)
  wire _038_;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:315" *)
  wire _039_;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:316" *)
  wire _040_;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:316" *)
  wire _041_;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:317" *)
  wire _042_;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:317" *)
  wire _043_;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:319" *)
  wire _044_;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:319" *)
  wire _045_;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:319" *)
  wire _046_;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:319" *)
  wire _047_;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:319" *)
  wire _048_;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:319" *)
  wire _049_;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:320" *)
  wire _050_;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:320" *)
  wire _051_;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:249" *)
  wire _052_;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:256" *)
  wire _053_;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:262" *)
  wire _054_;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:270" *)
  wire _055_;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:276" *)
  wire _056_;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:283" *)
  wire _057_;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:245" *)
  wire _058_;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:246" *)
  wire _059_;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:247" *)
  wire _060_;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:251" *)
  wire _061_;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:252" *)
  wire _062_;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:253" *)
  wire _063_;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:258" *)
  wire _064_;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:259" *)
  wire _065_;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:260" *)
  wire _066_;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:264" *)
  wire _067_;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:265" *)
  wire _068_;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:266" *)
  wire _069_;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:272" *)
  wire _070_;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:273" *)
  wire _071_;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:274" *)
  wire _072_;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:278" *)
  wire _073_;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:279" *)
  wire _074_;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:280" *)
  wire _075_;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:310" *)
  wire _076_;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:311" *)
  wire _077_;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:311" *)
  wire _078_;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:312" *)
  wire _079_;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:313" *)
  wire _080_;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:314" *)
  wire _081_;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:314" *)
  wire _082_;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:315" *)
  wire _083_;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:316" *)
  wire _084_;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:317" *)
  wire _085_;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:318" *)
  wire _086_;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:318" *)
  wire _087_;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:288" *)
  wire _088_;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:290" *)
  wire _089_;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:291" *)
  wire _090_;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:291" *)
  wire _091_;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:291" *)
  wire _092_;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:293" *)
  wire _093_;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:294" *)
  wire _094_;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:294" *)
  wire _095_;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:295" *)
  wire _096_;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:295" *)
  wire _097_;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:295" *)
  wire _098_;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:296" *)
  wire _099_;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:300" *)
  wire _100_;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:300" *)
  wire _101_;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:303" *)
  wire _102_;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:304" *)
  wire _103_;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:304" *)
  wire _104_;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:304" *)
  wire _105_;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:307" *)
  wire _106_;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:307" *)
  wire _107_;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:307" *)
  wire _108_;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:308" *)
  wire _109_;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:310" *)
  wire _110_;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:310" *)
  wire _111_;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:311" *)
  wire _112_;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:311" *)
  wire _113_;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:311" *)
  wire _114_;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:311" *)
  wire _115_;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:312" *)
  wire _116_;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:312" *)
  wire _117_;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:312" *)
  wire _118_;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:312" *)
  wire _119_;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:313" *)
  wire _120_;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:313" *)
  wire _121_;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:314" *)
  wire _122_;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:314" *)
  wire _123_;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:314" *)
  wire _124_;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:314" *)
  wire _125_;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:315" *)
  wire _126_;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:315" *)
  wire _127_;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:315" *)
  wire _128_;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:315" *)
  wire _129_;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:315" *)
  wire _130_;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:316" *)
  wire _131_;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:316" *)
  wire _132_;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:316" *)
  wire _133_;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:317" *)
  wire _134_;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:317" *)
  wire _135_;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:318" *)
  wire _136_;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:318" *)
  wire _137_;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:318" *)
  wire _138_;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:319" *)
  wire _139_;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:319" *)
  wire _140_;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:319" *)
  wire _141_;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:319" *)
  wire _142_;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:319" *)
  wire _143_;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:319" *)
  wire _144_;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:288" *)
  wire _145_;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:290" *)
  wire _146_;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:293" *)
  wire _147_;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:294" *)
  wire _148_;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:295" *)
  wire _149_;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:296" *)
  wire _150_;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:298" *)
  wire _151_;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:300" *)
  wire _152_;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:302" *)
  wire _153_;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:303" *)
  wire _154_;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:305" *)
  wire _155_;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:307" *)
  wire _156_;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:308" *)
  wire _157_;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:310" *)
  wire _158_;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:311" *)
  wire _159_;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:311" *)
  wire _160_;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:312" *)
  wire _161_;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:313" *)
  wire _162_;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:314" *)
  wire _163_;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:314" *)
  wire _164_;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:315" *)
  wire _165_;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:316" *)
  wire _166_;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:317" *)
  wire _167_;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:318" *)
  wire _168_;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:318" *)
  wire _169_;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:319" *)
  wire _170_;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:243" *)
  wire IntLeadZero_49U_leading_sign_49_0_rtn_IntLeadZero_49U_leading_sign_49_0_rtn_or_1_nl;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:240" *)
  wire IntLeadZero_49U_leading_sign_49_0_rtn_and_187_nl;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:239" *)
  wire IntLeadZero_49U_leading_sign_49_0_rtn_and_189_nl;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:241" *)
  wire IntLeadZero_49U_leading_sign_49_0_rtn_and_194_nl;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:242" *)
  wire IntLeadZero_49U_leading_sign_49_0_rtn_and_195_nl;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:224" *)
  wire IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_106_2_sdt_1;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:212" *)
  wire IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_110_3_sdt_3;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:225" *)
  wire IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_118_2_sdt_1;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:213" *)
  wire IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_118_2_sdt_2;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:226" *)
  wire IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_126_2_sdt_1;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:214" *)
  wire IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_134_4_sdt_4;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:216" *)
  wire IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_14_2_sdt_1;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:204" *)
  wire IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_18_3_sdt_3;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:217" *)
  wire IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_26_2_sdt_1;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:205" *)
  wire IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_26_2_sdt_2;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:218" *)
  wire IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_34_2_sdt_1;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:206" *)
  wire IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_42_4_sdt_4;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:219" *)
  wire IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_50_2_sdt_1;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:207" *)
  wire IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_50_2_sdt_2;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:220" *)
  wire IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_58_2_sdt_1;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:208" *)
  wire IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_62_3_sdt_3;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:215" *)
  wire IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_6_2_sdt_1;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:203" *)
  wire IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_6_2_sdt_2;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:221" *)
  wire IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_70_2_sdt_1;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:209" *)
  wire IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_70_2_sdt_2;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:222" *)
  wire IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_78_2_sdt_1;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:210" *)
  wire IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_90_5_sdt_5;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:223" *)
  wire IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_98_2_sdt_1;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:211" *)
  wire IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_98_2_sdt_2;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:231" *)
  wire c_h_1_12;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:232" *)
  wire c_h_1_13;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:233" *)
  wire c_h_1_14;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:234" *)
  wire c_h_1_17;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:227" *)
  wire c_h_1_2;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:235" *)
  wire c_h_1_20;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:236" *)
  wire c_h_1_21;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:237" *)
  wire c_h_1_22;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:238" *)
  wire c_h_1_23;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:228" *)
  wire c_h_1_5;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:229" *)
  wire c_h_1_6;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:230" *)
  wire c_h_1_9;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:200" *)
  input [48:0] mantissa;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:201" *)
  output [5:0] rtn;
  assign c_h_1_2 = IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_6_2_sdt_1 & (* src = "./vmod/vlibs/HLS_fp32_add.v:248" *) IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_6_2_sdt_2;
  assign IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_18_3_sdt_3 = _052_ & (* src = "./vmod/vlibs/HLS_fp32_add.v:250" *) IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_14_2_sdt_1;
  assign c_h_1_5 = IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_26_2_sdt_1 & (* src = "./vmod/vlibs/HLS_fp32_add.v:254" *) IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_26_2_sdt_2;
  assign c_h_1_6 = c_h_1_2 & (* src = "./vmod/vlibs/HLS_fp32_add.v:255" *) IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_18_3_sdt_3;
  assign _000_ = _053_ & (* src = "./vmod/vlibs/HLS_fp32_add.v:257" *) IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_34_2_sdt_1;
  assign IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_42_4_sdt_4 = _000_ & (* src = "./vmod/vlibs/HLS_fp32_add.v:257" *) c_h_1_5;
  assign c_h_1_9 = IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_50_2_sdt_1 & (* src = "./vmod/vlibs/HLS_fp32_add.v:261" *) IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_50_2_sdt_2;
  assign IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_62_3_sdt_3 = _054_ & (* src = "./vmod/vlibs/HLS_fp32_add.v:263" *) IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_58_2_sdt_1;
  assign c_h_1_12 = IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_70_2_sdt_1 & (* src = "./vmod/vlibs/HLS_fp32_add.v:267" *) IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_70_2_sdt_2;
  assign c_h_1_13 = c_h_1_9 & (* src = "./vmod/vlibs/HLS_fp32_add.v:268" *) IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_62_3_sdt_3;
  assign c_h_1_14 = c_h_1_6 & (* src = "./vmod/vlibs/HLS_fp32_add.v:269" *) IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_42_4_sdt_4;
  assign _001_ = _055_ & (* src = "./vmod/vlibs/HLS_fp32_add.v:271" *) IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_78_2_sdt_1;
  assign _002_ = _001_ & (* src = "./vmod/vlibs/HLS_fp32_add.v:271" *) c_h_1_12;
  assign IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_90_5_sdt_5 = _002_ & (* src = "./vmod/vlibs/HLS_fp32_add.v:271" *) c_h_1_13;
  assign c_h_1_17 = IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_98_2_sdt_1 & (* src = "./vmod/vlibs/HLS_fp32_add.v:275" *) IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_98_2_sdt_2;
  assign IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_110_3_sdt_3 = _056_ & (* src = "./vmod/vlibs/HLS_fp32_add.v:277" *) IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_106_2_sdt_1;
  assign c_h_1_20 = IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_118_2_sdt_1 & (* src = "./vmod/vlibs/HLS_fp32_add.v:281" *) IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_118_2_sdt_2;
  assign c_h_1_21 = c_h_1_17 & (* src = "./vmod/vlibs/HLS_fp32_add.v:282" *) IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_110_3_sdt_3;
  assign _003_ = _057_ & (* src = "./vmod/vlibs/HLS_fp32_add.v:284" *) IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_126_2_sdt_1;
  assign IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_134_4_sdt_4 = _003_ & (* src = "./vmod/vlibs/HLS_fp32_add.v:284" *) c_h_1_20;
  assign c_h_1_22 = c_h_1_21 & (* src = "./vmod/vlibs/HLS_fp32_add.v:285" *) IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_134_4_sdt_4;
  assign c_h_1_23 = c_h_1_14 & (* src = "./vmod/vlibs/HLS_fp32_add.v:286" *) IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_90_5_sdt_5;
  assign IntLeadZero_49U_leading_sign_49_0_rtn_and_189_nl = c_h_1_14 & (* src = "./vmod/vlibs/HLS_fp32_add.v:288" *) _145_;
  assign _004_ = c_h_1_6 & (* src = "./vmod/vlibs/HLS_fp32_add.v:290" *) _146_;
  assign _005_ = c_h_1_21 & (* src = "./vmod/vlibs/HLS_fp32_add.v:291" *) _090_;
  assign _006_ = _091_ & (* src = "./vmod/vlibs/HLS_fp32_add.v:291" *) c_h_1_23;
  assign IntLeadZero_49U_leading_sign_49_0_rtn_and_187_nl = _004_ & (* src = "./vmod/vlibs/HLS_fp32_add.v:291" *) _092_;
  assign _007_ = c_h_1_2 & (* src = "./vmod/vlibs/HLS_fp32_add.v:293" *) _147_;
  assign _008_ = c_h_1_9 & (* src = "./vmod/vlibs/HLS_fp32_add.v:294" *) _148_;
  assign _009_ = _095_ & (* src = "./vmod/vlibs/HLS_fp32_add.v:295" *) c_h_1_14;
  assign _010_ = _007_ & (* src = "./vmod/vlibs/HLS_fp32_add.v:295" *) _096_;
  assign _011_ = c_h_1_17 & (* src = "./vmod/vlibs/HLS_fp32_add.v:295" *) _149_;
  assign _012_ = _150_ & (* src = "./vmod/vlibs/HLS_fp32_add.v:296" *) c_h_1_23;
  assign IntLeadZero_49U_leading_sign_49_0_rtn_and_194_nl = _010_ & (* src = "./vmod/vlibs/HLS_fp32_add.v:296" *) _099_;
  assign _013_ = IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_6_2_sdt_1 & (* src = "./vmod/vlibs/HLS_fp32_add.v:299" *) _151_;
  assign _014_ = IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_26_2_sdt_1 & (* src = "./vmod/vlibs/HLS_fp32_add.v:300" *) _152_;
  assign _015_ = _100_ & (* src = "./vmod/vlibs/HLS_fp32_add.v:300" *) c_h_1_6;
  assign _016_ = _013_ & (* src = "./vmod/vlibs/HLS_fp32_add.v:301" *) _101_;
  assign _017_ = IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_50_2_sdt_1 & (* src = "./vmod/vlibs/HLS_fp32_add.v:302" *) _153_;
  assign _018_ = IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_70_2_sdt_1 & (* src = "./vmod/vlibs/HLS_fp32_add.v:303" *) _154_;
  assign _019_ = _102_ & (* src = "./vmod/vlibs/HLS_fp32_add.v:304" *) c_h_1_13;
  assign _020_ = _017_ & (* src = "./vmod/vlibs/HLS_fp32_add.v:304" *) _103_;
  assign _021_ = _104_ & (* src = "./vmod/vlibs/HLS_fp32_add.v:304" *) c_h_1_14;
  assign _022_ = _016_ & (* src = "./vmod/vlibs/HLS_fp32_add.v:304" *) _105_;
  assign _023_ = IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_98_2_sdt_1 & (* src = "./vmod/vlibs/HLS_fp32_add.v:306" *) _155_;
  assign _024_ = IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_118_2_sdt_1 & (* src = "./vmod/vlibs/HLS_fp32_add.v:307" *) _156_;
  assign _025_ = _106_ & (* src = "./vmod/vlibs/HLS_fp32_add.v:307" *) c_h_1_21;
  assign _026_ = _023_ & (* src = "./vmod/vlibs/HLS_fp32_add.v:307" *) _107_;
  assign _027_ = _157_ & (* src = "./vmod/vlibs/HLS_fp32_add.v:308" *) c_h_1_23;
  assign IntLeadZero_49U_leading_sign_49_0_rtn_and_195_nl = _022_ & (* src = "./vmod/vlibs/HLS_fp32_add.v:308" *) _109_;
  assign _028_ = _159_ & (* src = "./vmod/vlibs/HLS_fp32_add.v:311" *) c_h_1_2;
  assign _029_ = _111_ & (* src = "./vmod/vlibs/HLS_fp32_add.v:311" *) _113_;
  assign _030_ = _161_ & (* src = "./vmod/vlibs/HLS_fp32_add.v:312" *) c_h_1_5;
  assign _031_ = _115_ & (* src = "./vmod/vlibs/HLS_fp32_add.v:312" *) _117_;
  assign _032_ = _118_ & (* src = "./vmod/vlibs/HLS_fp32_add.v:312" *) c_h_1_6;
  assign _033_ = _029_ & (* src = "./vmod/vlibs/HLS_fp32_add.v:313" *) _119_;
  assign _034_ = _163_ & (* src = "./vmod/vlibs/HLS_fp32_add.v:314" *) c_h_1_9;
  assign _035_ = _121_ & (* src = "./vmod/vlibs/HLS_fp32_add.v:314" *) _123_;
  assign _036_ = _165_ & (* src = "./vmod/vlibs/HLS_fp32_add.v:315" *) c_h_1_12;
  assign _037_ = _125_ & (* src = "./vmod/vlibs/HLS_fp32_add.v:315" *) _127_;
  assign _038_ = _128_ & (* src = "./vmod/vlibs/HLS_fp32_add.v:315" *) c_h_1_13;
  assign _039_ = _035_ & (* src = "./vmod/vlibs/HLS_fp32_add.v:315" *) _129_;
  assign _040_ = _130_ & (* src = "./vmod/vlibs/HLS_fp32_add.v:316" *) c_h_1_14;
  assign _041_ = _033_ & (* src = "./vmod/vlibs/HLS_fp32_add.v:316" *) _131_;
  assign _042_ = _167_ & (* src = "./vmod/vlibs/HLS_fp32_add.v:317" *) c_h_1_17;
  assign _043_ = _133_ & (* src = "./vmod/vlibs/HLS_fp32_add.v:317" *) _135_;
  assign _044_ = _169_ & (* src = "./vmod/vlibs/HLS_fp32_add.v:319" *) c_h_1_20;
  assign _045_ = _137_ & (* src = "./vmod/vlibs/HLS_fp32_add.v:319" *) _139_;
  assign _046_ = _140_ & (* src = "./vmod/vlibs/HLS_fp32_add.v:319" *) c_h_1_21;
  assign _047_ = _043_ & (* src = "./vmod/vlibs/HLS_fp32_add.v:319" *) _141_;
  assign _048_ = _170_ & (* src = "./vmod/vlibs/HLS_fp32_add.v:319" *) c_h_1_23;
  assign _049_ = _041_ & (* src = "./vmod/vlibs/HLS_fp32_add.v:319" *) _143_;
  assign _050_ = _144_ & (* src = "./vmod/vlibs/HLS_fp32_add.v:320" *) c_h_1_22;
  assign _051_ = _050_ & (* src = "./vmod/vlibs/HLS_fp32_add.v:320" *) c_h_1_23;
  assign _052_ = ! (* src = "./vmod/vlibs/HLS_fp32_add.v:249" *) mantissa[42:41];
  assign _053_ = ! (* src = "./vmod/vlibs/HLS_fp32_add.v:256" *) mantissa[34:33];
  assign _054_ = ! (* src = "./vmod/vlibs/HLS_fp32_add.v:262" *) mantissa[26:25];
  assign _055_ = ! (* src = "./vmod/vlibs/HLS_fp32_add.v:270" *) mantissa[18:17];
  assign _056_ = ! (* src = "./vmod/vlibs/HLS_fp32_add.v:276" *) mantissa[10:9];
  assign _057_ = ! (* src = "./vmod/vlibs/HLS_fp32_add.v:283" *) mantissa[2:1];
  assign _058_ = | (* src = "./vmod/vlibs/HLS_fp32_add.v:245" *) mantissa[46:45];
  assign _059_ = | (* src = "./vmod/vlibs/HLS_fp32_add.v:246" *) mantissa[48:47];
  assign _060_ = | (* src = "./vmod/vlibs/HLS_fp32_add.v:247" *) mantissa[44:43];
  assign _061_ = | (* src = "./vmod/vlibs/HLS_fp32_add.v:251" *) mantissa[38:37];
  assign _062_ = | (* src = "./vmod/vlibs/HLS_fp32_add.v:252" *) mantissa[40:39];
  assign _063_ = | (* src = "./vmod/vlibs/HLS_fp32_add.v:253" *) mantissa[36:35];
  assign _064_ = | (* src = "./vmod/vlibs/HLS_fp32_add.v:258" *) mantissa[30:29];
  assign _065_ = | (* src = "./vmod/vlibs/HLS_fp32_add.v:259" *) mantissa[32:31];
  assign _066_ = | (* src = "./vmod/vlibs/HLS_fp32_add.v:260" *) mantissa[28:27];
  assign _067_ = | (* src = "./vmod/vlibs/HLS_fp32_add.v:264" *) mantissa[22:21];
  assign _068_ = | (* src = "./vmod/vlibs/HLS_fp32_add.v:265" *) mantissa[24:23];
  assign _069_ = | (* src = "./vmod/vlibs/HLS_fp32_add.v:266" *) mantissa[20:19];
  assign _070_ = | (* src = "./vmod/vlibs/HLS_fp32_add.v:272" *) mantissa[14:13];
  assign _071_ = | (* src = "./vmod/vlibs/HLS_fp32_add.v:273" *) mantissa[16:15];
  assign _072_ = | (* src = "./vmod/vlibs/HLS_fp32_add.v:274" *) mantissa[12:11];
  assign _073_ = | (* src = "./vmod/vlibs/HLS_fp32_add.v:278" *) mantissa[6:5];
  assign _074_ = | (* src = "./vmod/vlibs/HLS_fp32_add.v:279" *) mantissa[8:7];
  assign _075_ = | (* src = "./vmod/vlibs/HLS_fp32_add.v:280" *) mantissa[4:3];
  assign _076_ = mantissa[47:46] != (* src = "./vmod/vlibs/HLS_fp32_add.v:310" *) 1'b1;
  assign _077_ = mantissa[43:42] != (* src = "./vmod/vlibs/HLS_fp32_add.v:311" *) 1'b1;
  assign _078_ = mantissa[39:38] != (* src = "./vmod/vlibs/HLS_fp32_add.v:311" *) 1'b1;
  assign _079_ = mantissa[35:34] != (* src = "./vmod/vlibs/HLS_fp32_add.v:312" *) 1'b1;
  assign _080_ = mantissa[31:30] != (* src = "./vmod/vlibs/HLS_fp32_add.v:313" *) 1'b1;
  assign _081_ = mantissa[27:26] != (* src = "./vmod/vlibs/HLS_fp32_add.v:314" *) 1'b1;
  assign _082_ = mantissa[23:22] != (* src = "./vmod/vlibs/HLS_fp32_add.v:314" *) 1'b1;
  assign _083_ = mantissa[19:18] != (* src = "./vmod/vlibs/HLS_fp32_add.v:315" *) 1'b1;
  assign _084_ = mantissa[15:14] != (* src = "./vmod/vlibs/HLS_fp32_add.v:316" *) 1'b1;
  assign _085_ = mantissa[11:10] != (* src = "./vmod/vlibs/HLS_fp32_add.v:317" *) 1'b1;
  assign _086_ = mantissa[7:6] != (* src = "./vmod/vlibs/HLS_fp32_add.v:318" *) 1'b1;
  assign _087_ = mantissa[3:2] != (* src = "./vmod/vlibs/HLS_fp32_add.v:318" *) 1'b1;
  assign IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_6_2_sdt_2 = ~ (* src = "./vmod/vlibs/HLS_fp32_add.v:245" *) _058_;
  assign IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_6_2_sdt_1 = ~ (* src = "./vmod/vlibs/HLS_fp32_add.v:246" *) _059_;
  assign IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_14_2_sdt_1 = ~ (* src = "./vmod/vlibs/HLS_fp32_add.v:247" *) _060_;
  assign IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_26_2_sdt_2 = ~ (* src = "./vmod/vlibs/HLS_fp32_add.v:251" *) _061_;
  assign IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_26_2_sdt_1 = ~ (* src = "./vmod/vlibs/HLS_fp32_add.v:252" *) _062_;
  assign IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_34_2_sdt_1 = ~ (* src = "./vmod/vlibs/HLS_fp32_add.v:253" *) _063_;
  assign IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_50_2_sdt_2 = ~ (* src = "./vmod/vlibs/HLS_fp32_add.v:258" *) _064_;
  assign IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_50_2_sdt_1 = ~ (* src = "./vmod/vlibs/HLS_fp32_add.v:259" *) _065_;
  assign IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_58_2_sdt_1 = ~ (* src = "./vmod/vlibs/HLS_fp32_add.v:260" *) _066_;
  assign IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_70_2_sdt_2 = ~ (* src = "./vmod/vlibs/HLS_fp32_add.v:264" *) _067_;
  assign IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_70_2_sdt_1 = ~ (* src = "./vmod/vlibs/HLS_fp32_add.v:265" *) _068_;
  assign IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_78_2_sdt_1 = ~ (* src = "./vmod/vlibs/HLS_fp32_add.v:266" *) _069_;
  assign IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_98_2_sdt_2 = ~ (* src = "./vmod/vlibs/HLS_fp32_add.v:272" *) _070_;
  assign IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_98_2_sdt_1 = ~ (* src = "./vmod/vlibs/HLS_fp32_add.v:273" *) _071_;
  assign IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_106_2_sdt_1 = ~ (* src = "./vmod/vlibs/HLS_fp32_add.v:274" *) _072_;
  assign IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_118_2_sdt_2 = ~ (* src = "./vmod/vlibs/HLS_fp32_add.v:278" *) _073_;
  assign IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_118_2_sdt_1 = ~ (* src = "./vmod/vlibs/HLS_fp32_add.v:279" *) _074_;
  assign IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_126_2_sdt_1 = ~ (* src = "./vmod/vlibs/HLS_fp32_add.v:280" *) _075_;
  assign _088_ = ~ (* src = "./vmod/vlibs/HLS_fp32_add.v:288" *) IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_90_5_sdt_5;
  assign _089_ = ~ (* src = "./vmod/vlibs/HLS_fp32_add.v:290" *) IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_42_4_sdt_4;
  assign _090_ = ~ (* src = "./vmod/vlibs/HLS_fp32_add.v:291" *) IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_134_4_sdt_4;
  assign _091_ = ~ (* src = "./vmod/vlibs/HLS_fp32_add.v:291" *) _005_;
  assign _092_ = ~ (* src = "./vmod/vlibs/HLS_fp32_add.v:291" *) _006_;
  assign _093_ = ~ (* src = "./vmod/vlibs/HLS_fp32_add.v:293" *) IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_18_3_sdt_3;
  assign _094_ = ~ (* src = "./vmod/vlibs/HLS_fp32_add.v:294" *) IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_62_3_sdt_3;
  assign _095_ = ~ (* src = "./vmod/vlibs/HLS_fp32_add.v:294" *) _008_;
  assign _096_ = ~ (* src = "./vmod/vlibs/HLS_fp32_add.v:295" *) _009_;
  assign _097_ = ~ (* src = "./vmod/vlibs/HLS_fp32_add.v:295" *) IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_110_3_sdt_3;
  assign _098_ = ~ (* src = "./vmod/vlibs/HLS_fp32_add.v:295" *) _011_;
  assign _099_ = ~ (* src = "./vmod/vlibs/HLS_fp32_add.v:296" *) _012_;
  assign _100_ = ~ (* src = "./vmod/vlibs/HLS_fp32_add.v:300" *) _014_;
  assign _101_ = ~ (* src = "./vmod/vlibs/HLS_fp32_add.v:300" *) _015_;
  assign _102_ = ~ (* src = "./vmod/vlibs/HLS_fp32_add.v:303" *) _018_;
  assign _103_ = ~ (* src = "./vmod/vlibs/HLS_fp32_add.v:304" *) _019_;
  assign _104_ = ~ (* src = "./vmod/vlibs/HLS_fp32_add.v:304" *) _020_;
  assign _105_ = ~ (* src = "./vmod/vlibs/HLS_fp32_add.v:304" *) _021_;
  assign _106_ = ~ (* src = "./vmod/vlibs/HLS_fp32_add.v:307" *) _024_;
  assign _107_ = ~ (* src = "./vmod/vlibs/HLS_fp32_add.v:307" *) _025_;
  assign _108_ = ~ (* src = "./vmod/vlibs/HLS_fp32_add.v:307" *) _026_;
  assign _109_ = ~ (* src = "./vmod/vlibs/HLS_fp32_add.v:308" *) _027_;
  assign _110_ = ~ (* src = "./vmod/vlibs/HLS_fp32_add.v:310" *) _076_;
  assign _111_ = ~ (* src = "./vmod/vlibs/HLS_fp32_add.v:310" *) _158_;
  assign _112_ = ~ (* src = "./vmod/vlibs/HLS_fp32_add.v:311" *) _077_;
  assign _113_ = ~ (* src = "./vmod/vlibs/HLS_fp32_add.v:311" *) _028_;
  assign _114_ = ~ (* src = "./vmod/vlibs/HLS_fp32_add.v:311" *) _078_;
  assign _115_ = ~ (* src = "./vmod/vlibs/HLS_fp32_add.v:311" *) _160_;
  assign _116_ = ~ (* src = "./vmod/vlibs/HLS_fp32_add.v:312" *) _079_;
  assign _117_ = ~ (* src = "./vmod/vlibs/HLS_fp32_add.v:312" *) _030_;
  assign _118_ = ~ (* src = "./vmod/vlibs/HLS_fp32_add.v:312" *) _031_;
  assign _119_ = ~ (* src = "./vmod/vlibs/HLS_fp32_add.v:312" *) _032_;
  assign _120_ = ~ (* src = "./vmod/vlibs/HLS_fp32_add.v:313" *) _080_;
  assign _121_ = ~ (* src = "./vmod/vlibs/HLS_fp32_add.v:313" *) _162_;
  assign _122_ = ~ (* src = "./vmod/vlibs/HLS_fp32_add.v:314" *) _081_;
  assign _123_ = ~ (* src = "./vmod/vlibs/HLS_fp32_add.v:314" *) _034_;
  assign _124_ = ~ (* src = "./vmod/vlibs/HLS_fp32_add.v:314" *) _082_;
  assign _125_ = ~ (* src = "./vmod/vlibs/HLS_fp32_add.v:314" *) _164_;
  assign _126_ = ~ (* src = "./vmod/vlibs/HLS_fp32_add.v:315" *) _083_;
  assign _127_ = ~ (* src = "./vmod/vlibs/HLS_fp32_add.v:315" *) _036_;
  assign _128_ = ~ (* src = "./vmod/vlibs/HLS_fp32_add.v:315" *) _037_;
  assign _129_ = ~ (* src = "./vmod/vlibs/HLS_fp32_add.v:315" *) _038_;
  assign _130_ = ~ (* src = "./vmod/vlibs/HLS_fp32_add.v:315" *) _039_;
  assign _131_ = ~ (* src = "./vmod/vlibs/HLS_fp32_add.v:316" *) _040_;
  assign _132_ = ~ (* src = "./vmod/vlibs/HLS_fp32_add.v:316" *) _084_;
  assign _133_ = ~ (* src = "./vmod/vlibs/HLS_fp32_add.v:316" *) _166_;
  assign _134_ = ~ (* src = "./vmod/vlibs/HLS_fp32_add.v:317" *) _085_;
  assign _135_ = ~ (* src = "./vmod/vlibs/HLS_fp32_add.v:317" *) _042_;
  assign _136_ = ~ (* src = "./vmod/vlibs/HLS_fp32_add.v:318" *) _086_;
  assign _137_ = ~ (* src = "./vmod/vlibs/HLS_fp32_add.v:318" *) _168_;
  assign _138_ = ~ (* src = "./vmod/vlibs/HLS_fp32_add.v:318" *) _087_;
  assign _139_ = ~ (* src = "./vmod/vlibs/HLS_fp32_add.v:319" *) _044_;
  assign _140_ = ~ (* src = "./vmod/vlibs/HLS_fp32_add.v:319" *) _045_;
  assign _141_ = ~ (* src = "./vmod/vlibs/HLS_fp32_add.v:319" *) _046_;
  assign _142_ = ~ (* src = "./vmod/vlibs/HLS_fp32_add.v:319" *) _047_;
  assign _143_ = ~ (* src = "./vmod/vlibs/HLS_fp32_add.v:319" *) _048_;
  assign _144_ = ~ (* src = "./vmod/vlibs/HLS_fp32_add.v:319" *) mantissa[0];
  assign _145_ = c_h_1_22 | (* src = "./vmod/vlibs/HLS_fp32_add.v:288" *) _088_;
  assign _146_ = c_h_1_13 | (* src = "./vmod/vlibs/HLS_fp32_add.v:290" *) _089_;
  assign _147_ = c_h_1_5 | (* src = "./vmod/vlibs/HLS_fp32_add.v:293" *) _093_;
  assign _148_ = c_h_1_12 | (* src = "./vmod/vlibs/HLS_fp32_add.v:294" *) _094_;
  assign _149_ = c_h_1_20 | (* src = "./vmod/vlibs/HLS_fp32_add.v:295" *) _097_;
  assign _150_ = _098_ | (* src = "./vmod/vlibs/HLS_fp32_add.v:296" *) c_h_1_22;
  assign _151_ = IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_14_2_sdt_1 | (* src = "./vmod/vlibs/HLS_fp32_add.v:298" *) _058_;
  assign _152_ = IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_34_2_sdt_1 | (* src = "./vmod/vlibs/HLS_fp32_add.v:300" *) _061_;
  assign _153_ = IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_58_2_sdt_1 | (* src = "./vmod/vlibs/HLS_fp32_add.v:302" *) _064_;
  assign _154_ = IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_78_2_sdt_1 | (* src = "./vmod/vlibs/HLS_fp32_add.v:303" *) _067_;
  assign _155_ = IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_106_2_sdt_1 | (* src = "./vmod/vlibs/HLS_fp32_add.v:305" *) _070_;
  assign _156_ = IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_126_2_sdt_1 | (* src = "./vmod/vlibs/HLS_fp32_add.v:307" *) _073_;
  assign _157_ = _108_ | (* src = "./vmod/vlibs/HLS_fp32_add.v:308" *) c_h_1_22;
  assign _158_ = mantissa[48] | (* src = "./vmod/vlibs/HLS_fp32_add.v:310" *) _110_;
  assign _159_ = mantissa[44] | (* src = "./vmod/vlibs/HLS_fp32_add.v:311" *) _112_;
  assign _160_ = mantissa[40] | (* src = "./vmod/vlibs/HLS_fp32_add.v:311" *) _114_;
  assign _161_ = mantissa[36] | (* src = "./vmod/vlibs/HLS_fp32_add.v:312" *) _116_;
  assign _162_ = mantissa[32] | (* src = "./vmod/vlibs/HLS_fp32_add.v:313" *) _120_;
  assign _163_ = mantissa[28] | (* src = "./vmod/vlibs/HLS_fp32_add.v:314" *) _122_;
  assign _164_ = mantissa[24] | (* src = "./vmod/vlibs/HLS_fp32_add.v:314" *) _124_;
  assign _165_ = mantissa[20] | (* src = "./vmod/vlibs/HLS_fp32_add.v:315" *) _126_;
  assign _166_ = mantissa[16] | (* src = "./vmod/vlibs/HLS_fp32_add.v:316" *) _132_;
  assign _167_ = mantissa[12] | (* src = "./vmod/vlibs/HLS_fp32_add.v:317" *) _134_;
  assign _168_ = mantissa[8] | (* src = "./vmod/vlibs/HLS_fp32_add.v:318" *) _136_;
  assign _169_ = mantissa[4] | (* src = "./vmod/vlibs/HLS_fp32_add.v:318" *) _138_;
  assign _170_ = _142_ | (* src = "./vmod/vlibs/HLS_fp32_add.v:319" *) c_h_1_22;
  assign IntLeadZero_49U_leading_sign_49_0_rtn_IntLeadZero_49U_leading_sign_49_0_rtn_or_1_nl = _049_ | (* src = "./vmod/vlibs/HLS_fp32_add.v:320" *) _051_;
  assign rtn = { c_h_1_23, IntLeadZero_49U_leading_sign_49_0_rtn_and_189_nl, IntLeadZero_49U_leading_sign_49_0_rtn_and_187_nl, IntLeadZero_49U_leading_sign_49_0_rtn_and_194_nl, IntLeadZero_49U_leading_sign_49_0_rtn_and_195_nl, IntLeadZero_49U_leading_sign_49_0_rtn_IntLeadZero_49U_leading_sign_49_0_rtn_or_1_nl };
endmodule
