module SDP_X_leading_sign_49_0(mantissa, rtn);
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:467" *)
  wire _000_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:481" *)
  wire _001_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:481" *)
  wire _002_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:494" *)
  wire _003_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:500" *)
  wire _004_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:501" *)
  wire _005_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:501" *)
  wire _006_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:503" *)
  wire _007_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:504" *)
  wire _008_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:505" *)
  wire _009_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:505" *)
  wire _010_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:505" *)
  wire _011_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:506" *)
  wire _012_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:509" *)
  wire _013_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:510" *)
  wire _014_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:510" *)
  wire _015_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:511" *)
  wire _016_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:512" *)
  wire _017_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:513" *)
  wire _018_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:514" *)
  wire _019_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:514" *)
  wire _020_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:514" *)
  wire _021_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:514" *)
  wire _022_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:516" *)
  wire _023_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:517" *)
  wire _024_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:517" *)
  wire _025_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:517" *)
  wire _026_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:518" *)
  wire _027_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:521" *)
  wire _028_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:521" *)
  wire _029_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:522" *)
  wire _030_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:522" *)
  wire _031_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:522" *)
  wire _032_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:523" *)
  wire _033_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:524" *)
  wire _034_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:524" *)
  wire _035_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:525" *)
  wire _036_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:525" *)
  wire _037_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:525" *)
  wire _038_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:525" *)
  wire _039_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:526" *)
  wire _040_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:526" *)
  wire _041_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:527" *)
  wire _042_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:527" *)
  wire _043_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:529" *)
  wire _044_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:529" *)
  wire _045_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:529" *)
  wire _046_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:529" *)
  wire _047_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:529" *)
  wire _048_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:529" *)
  wire _049_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:530" *)
  wire _050_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:530" *)
  wire _051_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:459" *)
  wire _052_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:466" *)
  wire _053_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:472" *)
  wire _054_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:480" *)
  wire _055_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:486" *)
  wire _056_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:493" *)
  wire _057_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:455" *)
  wire _058_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:456" *)
  wire _059_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:457" *)
  wire _060_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:461" *)
  wire _061_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:462" *)
  wire _062_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:463" *)
  wire _063_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:468" *)
  wire _064_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:469" *)
  wire _065_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:470" *)
  wire _066_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:474" *)
  wire _067_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:475" *)
  wire _068_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:476" *)
  wire _069_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:482" *)
  wire _070_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:483" *)
  wire _071_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:484" *)
  wire _072_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:488" *)
  wire _073_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:489" *)
  wire _074_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:490" *)
  wire _075_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:520" *)
  wire _076_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:521" *)
  wire _077_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:521" *)
  wire _078_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:522" *)
  wire _079_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:523" *)
  wire _080_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:524" *)
  wire _081_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:524" *)
  wire _082_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:525" *)
  wire _083_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:526" *)
  wire _084_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:527" *)
  wire _085_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:528" *)
  wire _086_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:528" *)
  wire _087_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:498" *)
  wire _088_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:500" *)
  wire _089_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:501" *)
  wire _090_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:501" *)
  wire _091_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:501" *)
  wire _092_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:503" *)
  wire _093_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:504" *)
  wire _094_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:504" *)
  wire _095_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:505" *)
  wire _096_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:505" *)
  wire _097_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:505" *)
  wire _098_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:506" *)
  wire _099_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:510" *)
  wire _100_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:510" *)
  wire _101_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:513" *)
  wire _102_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:514" *)
  wire _103_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:514" *)
  wire _104_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:514" *)
  wire _105_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:517" *)
  wire _106_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:517" *)
  wire _107_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:517" *)
  wire _108_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:518" *)
  wire _109_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:520" *)
  wire _110_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:520" *)
  wire _111_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:521" *)
  wire _112_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:521" *)
  wire _113_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:521" *)
  wire _114_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:521" *)
  wire _115_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:522" *)
  wire _116_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:522" *)
  wire _117_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:522" *)
  wire _118_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:522" *)
  wire _119_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:523" *)
  wire _120_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:523" *)
  wire _121_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:524" *)
  wire _122_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:524" *)
  wire _123_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:524" *)
  wire _124_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:524" *)
  wire _125_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:525" *)
  wire _126_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:525" *)
  wire _127_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:525" *)
  wire _128_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:525" *)
  wire _129_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:525" *)
  wire _130_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:526" *)
  wire _131_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:526" *)
  wire _132_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:526" *)
  wire _133_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:527" *)
  wire _134_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:527" *)
  wire _135_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:528" *)
  wire _136_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:528" *)
  wire _137_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:528" *)
  wire _138_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:529" *)
  wire _139_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:529" *)
  wire _140_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:529" *)
  wire _141_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:529" *)
  wire _142_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:529" *)
  wire _143_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:529" *)
  wire _144_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:498" *)
  wire _145_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:500" *)
  wire _146_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:503" *)
  wire _147_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:504" *)
  wire _148_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:505" *)
  wire _149_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:506" *)
  wire _150_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:508" *)
  wire _151_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:510" *)
  wire _152_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:512" *)
  wire _153_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:513" *)
  wire _154_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:515" *)
  wire _155_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:517" *)
  wire _156_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:518" *)
  wire _157_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:520" *)
  wire _158_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:521" *)
  wire _159_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:521" *)
  wire _160_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:522" *)
  wire _161_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:523" *)
  wire _162_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:524" *)
  wire _163_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:524" *)
  wire _164_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:525" *)
  wire _165_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:526" *)
  wire _166_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:527" *)
  wire _167_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:528" *)
  wire _168_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:528" *)
  wire _169_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:529" *)
  wire _170_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:453" *)
  wire IntLeadZero_49U_leading_sign_49_0_rtn_IntLeadZero_49U_leading_sign_49_0_rtn_or_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:450" *)
  wire IntLeadZero_49U_leading_sign_49_0_rtn_and_187_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:449" *)
  wire IntLeadZero_49U_leading_sign_49_0_rtn_and_189_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:451" *)
  wire IntLeadZero_49U_leading_sign_49_0_rtn_and_194_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:452" *)
  wire IntLeadZero_49U_leading_sign_49_0_rtn_and_195_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:434" *)
  wire IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_106_2_sdt_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:422" *)
  wire IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_110_3_sdt_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:435" *)
  wire IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_118_2_sdt_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:423" *)
  wire IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_118_2_sdt_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:436" *)
  wire IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_126_2_sdt_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:424" *)
  wire IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_134_4_sdt_4;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:426" *)
  wire IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_14_2_sdt_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:414" *)
  wire IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_18_3_sdt_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:427" *)
  wire IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_26_2_sdt_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:415" *)
  wire IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_26_2_sdt_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:428" *)
  wire IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_34_2_sdt_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:416" *)
  wire IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_42_4_sdt_4;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:429" *)
  wire IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_50_2_sdt_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:417" *)
  wire IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_50_2_sdt_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:430" *)
  wire IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_58_2_sdt_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:418" *)
  wire IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_62_3_sdt_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:425" *)
  wire IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_6_2_sdt_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:413" *)
  wire IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_6_2_sdt_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:431" *)
  wire IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_70_2_sdt_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:419" *)
  wire IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_70_2_sdt_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:432" *)
  wire IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_78_2_sdt_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:420" *)
  wire IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_90_5_sdt_5;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:433" *)
  wire IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_98_2_sdt_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:421" *)
  wire IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_98_2_sdt_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:441" *)
  wire c_h_1_12;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:442" *)
  wire c_h_1_13;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:443" *)
  wire c_h_1_14;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:444" *)
  wire c_h_1_17;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:437" *)
  wire c_h_1_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:445" *)
  wire c_h_1_20;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:446" *)
  wire c_h_1_21;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:447" *)
  wire c_h_1_22;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:448" *)
  wire c_h_1_23;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:438" *)
  wire c_h_1_5;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:439" *)
  wire c_h_1_6;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:440" *)
  wire c_h_1_9;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:410" *)
  input [48:0] mantissa;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:411" *)
  output [5:0] rtn;
  assign c_h_1_2 = IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_6_2_sdt_1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:458" *) IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_6_2_sdt_2;
  assign IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_18_3_sdt_3 = _052_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:460" *) IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_14_2_sdt_1;
  assign c_h_1_5 = IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_26_2_sdt_1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:464" *) IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_26_2_sdt_2;
  assign c_h_1_6 = c_h_1_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:465" *) IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_18_3_sdt_3;
  assign _000_ = _053_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:467" *) IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_34_2_sdt_1;
  assign IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_42_4_sdt_4 = _000_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:467" *) c_h_1_5;
  assign c_h_1_9 = IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_50_2_sdt_1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:471" *) IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_50_2_sdt_2;
  assign IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_62_3_sdt_3 = _054_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:473" *) IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_58_2_sdt_1;
  assign c_h_1_12 = IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_70_2_sdt_1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:477" *) IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_70_2_sdt_2;
  assign c_h_1_13 = c_h_1_9 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:478" *) IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_62_3_sdt_3;
  assign c_h_1_14 = c_h_1_6 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:479" *) IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_42_4_sdt_4;
  assign _001_ = _055_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:481" *) IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_78_2_sdt_1;
  assign _002_ = _001_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:481" *) c_h_1_12;
  assign IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_90_5_sdt_5 = _002_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:481" *) c_h_1_13;
  assign c_h_1_17 = IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_98_2_sdt_1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:485" *) IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_98_2_sdt_2;
  assign IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_110_3_sdt_3 = _056_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:487" *) IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_106_2_sdt_1;
  assign c_h_1_20 = IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_118_2_sdt_1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:491" *) IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_118_2_sdt_2;
  assign c_h_1_21 = c_h_1_17 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:492" *) IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_110_3_sdt_3;
  assign _003_ = _057_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:494" *) IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_126_2_sdt_1;
  assign IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_134_4_sdt_4 = _003_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:494" *) c_h_1_20;
  assign c_h_1_22 = c_h_1_21 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:495" *) IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_134_4_sdt_4;
  assign c_h_1_23 = c_h_1_14 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:496" *) IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_90_5_sdt_5;
  assign IntLeadZero_49U_leading_sign_49_0_rtn_and_189_nl = c_h_1_14 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:498" *) _145_;
  assign _004_ = c_h_1_6 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:500" *) _146_;
  assign _005_ = c_h_1_21 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:501" *) _090_;
  assign _006_ = _091_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:501" *) c_h_1_23;
  assign IntLeadZero_49U_leading_sign_49_0_rtn_and_187_nl = _004_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:501" *) _092_;
  assign _007_ = c_h_1_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:503" *) _147_;
  assign _008_ = c_h_1_9 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:504" *) _148_;
  assign _009_ = _095_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:505" *) c_h_1_14;
  assign _010_ = _007_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:505" *) _096_;
  assign _011_ = c_h_1_17 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:505" *) _149_;
  assign _012_ = _150_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:506" *) c_h_1_23;
  assign IntLeadZero_49U_leading_sign_49_0_rtn_and_194_nl = _010_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:506" *) _099_;
  assign _013_ = IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_6_2_sdt_1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:509" *) _151_;
  assign _014_ = IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_26_2_sdt_1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:510" *) _152_;
  assign _015_ = _100_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:510" *) c_h_1_6;
  assign _016_ = _013_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:511" *) _101_;
  assign _017_ = IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_50_2_sdt_1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:512" *) _153_;
  assign _018_ = IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_70_2_sdt_1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:513" *) _154_;
  assign _019_ = _102_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:514" *) c_h_1_13;
  assign _020_ = _017_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:514" *) _103_;
  assign _021_ = _104_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:514" *) c_h_1_14;
  assign _022_ = _016_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:514" *) _105_;
  assign _023_ = IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_98_2_sdt_1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:516" *) _155_;
  assign _024_ = IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_118_2_sdt_1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:517" *) _156_;
  assign _025_ = _106_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:517" *) c_h_1_21;
  assign _026_ = _023_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:517" *) _107_;
  assign _027_ = _157_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:518" *) c_h_1_23;
  assign IntLeadZero_49U_leading_sign_49_0_rtn_and_195_nl = _022_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:518" *) _109_;
  assign _028_ = _159_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:521" *) c_h_1_2;
  assign _029_ = _111_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:521" *) _113_;
  assign _030_ = _161_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:522" *) c_h_1_5;
  assign _031_ = _115_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:522" *) _117_;
  assign _032_ = _118_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:522" *) c_h_1_6;
  assign _033_ = _029_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:523" *) _119_;
  assign _034_ = _163_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:524" *) c_h_1_9;
  assign _035_ = _121_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:524" *) _123_;
  assign _036_ = _165_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:525" *) c_h_1_12;
  assign _037_ = _125_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:525" *) _127_;
  assign _038_ = _128_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:525" *) c_h_1_13;
  assign _039_ = _035_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:525" *) _129_;
  assign _040_ = _130_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:526" *) c_h_1_14;
  assign _041_ = _033_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:526" *) _131_;
  assign _042_ = _167_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:527" *) c_h_1_17;
  assign _043_ = _133_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:527" *) _135_;
  assign _044_ = _169_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:529" *) c_h_1_20;
  assign _045_ = _137_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:529" *) _139_;
  assign _046_ = _140_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:529" *) c_h_1_21;
  assign _047_ = _043_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:529" *) _141_;
  assign _048_ = _170_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:529" *) c_h_1_23;
  assign _049_ = _041_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:529" *) _143_;
  assign _050_ = _144_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:530" *) c_h_1_22;
  assign _051_ = _050_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:530" *) c_h_1_23;
  assign _052_ = ! (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:459" *) mantissa[42:41];
  assign _053_ = ! (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:466" *) mantissa[34:33];
  assign _054_ = ! (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:472" *) mantissa[26:25];
  assign _055_ = ! (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:480" *) mantissa[18:17];
  assign _056_ = ! (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:486" *) mantissa[10:9];
  assign _057_ = ! (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:493" *) mantissa[2:1];
  assign _058_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:455" *) mantissa[46:45];
  assign _059_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:456" *) mantissa[48:47];
  assign _060_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:457" *) mantissa[44:43];
  assign _061_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:461" *) mantissa[38:37];
  assign _062_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:462" *) mantissa[40:39];
  assign _063_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:463" *) mantissa[36:35];
  assign _064_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:468" *) mantissa[30:29];
  assign _065_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:469" *) mantissa[32:31];
  assign _066_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:470" *) mantissa[28:27];
  assign _067_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:474" *) mantissa[22:21];
  assign _068_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:475" *) mantissa[24:23];
  assign _069_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:476" *) mantissa[20:19];
  assign _070_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:482" *) mantissa[14:13];
  assign _071_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:483" *) mantissa[16:15];
  assign _072_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:484" *) mantissa[12:11];
  assign _073_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:488" *) mantissa[6:5];
  assign _074_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:489" *) mantissa[8:7];
  assign _075_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:490" *) mantissa[4:3];
  assign _076_ = mantissa[47:46] != (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:520" *) 1'b1;
  assign _077_ = mantissa[43:42] != (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:521" *) 1'b1;
  assign _078_ = mantissa[39:38] != (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:521" *) 1'b1;
  assign _079_ = mantissa[35:34] != (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:522" *) 1'b1;
  assign _080_ = mantissa[31:30] != (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:523" *) 1'b1;
  assign _081_ = mantissa[27:26] != (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:524" *) 1'b1;
  assign _082_ = mantissa[23:22] != (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:524" *) 1'b1;
  assign _083_ = mantissa[19:18] != (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:525" *) 1'b1;
  assign _084_ = mantissa[15:14] != (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:526" *) 1'b1;
  assign _085_ = mantissa[11:10] != (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:527" *) 1'b1;
  assign _086_ = mantissa[7:6] != (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:528" *) 1'b1;
  assign _087_ = mantissa[3:2] != (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:528" *) 1'b1;
  assign IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_6_2_sdt_2 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:455" *) _058_;
  assign IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_6_2_sdt_1 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:456" *) _059_;
  assign IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_14_2_sdt_1 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:457" *) _060_;
  assign IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_26_2_sdt_2 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:461" *) _061_;
  assign IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_26_2_sdt_1 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:462" *) _062_;
  assign IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_34_2_sdt_1 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:463" *) _063_;
  assign IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_50_2_sdt_2 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:468" *) _064_;
  assign IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_50_2_sdt_1 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:469" *) _065_;
  assign IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_58_2_sdt_1 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:470" *) _066_;
  assign IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_70_2_sdt_2 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:474" *) _067_;
  assign IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_70_2_sdt_1 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:475" *) _068_;
  assign IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_78_2_sdt_1 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:476" *) _069_;
  assign IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_98_2_sdt_2 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:482" *) _070_;
  assign IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_98_2_sdt_1 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:483" *) _071_;
  assign IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_106_2_sdt_1 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:484" *) _072_;
  assign IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_118_2_sdt_2 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:488" *) _073_;
  assign IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_118_2_sdt_1 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:489" *) _074_;
  assign IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_126_2_sdt_1 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:490" *) _075_;
  assign _088_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:498" *) IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_90_5_sdt_5;
  assign _089_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:500" *) IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_42_4_sdt_4;
  assign _090_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:501" *) IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_134_4_sdt_4;
  assign _091_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:501" *) _005_;
  assign _092_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:501" *) _006_;
  assign _093_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:503" *) IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_18_3_sdt_3;
  assign _094_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:504" *) IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_62_3_sdt_3;
  assign _095_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:504" *) _008_;
  assign _096_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:505" *) _009_;
  assign _097_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:505" *) IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_110_3_sdt_3;
  assign _098_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:505" *) _011_;
  assign _099_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:506" *) _012_;
  assign _100_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:510" *) _014_;
  assign _101_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:510" *) _015_;
  assign _102_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:513" *) _018_;
  assign _103_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:514" *) _019_;
  assign _104_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:514" *) _020_;
  assign _105_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:514" *) _021_;
  assign _106_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:517" *) _024_;
  assign _107_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:517" *) _025_;
  assign _108_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:517" *) _026_;
  assign _109_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:518" *) _027_;
  assign _110_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:520" *) _076_;
  assign _111_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:520" *) _158_;
  assign _112_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:521" *) _077_;
  assign _113_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:521" *) _028_;
  assign _114_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:521" *) _078_;
  assign _115_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:521" *) _160_;
  assign _116_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:522" *) _079_;
  assign _117_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:522" *) _030_;
  assign _118_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:522" *) _031_;
  assign _119_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:522" *) _032_;
  assign _120_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:523" *) _080_;
  assign _121_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:523" *) _162_;
  assign _122_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:524" *) _081_;
  assign _123_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:524" *) _034_;
  assign _124_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:524" *) _082_;
  assign _125_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:524" *) _164_;
  assign _126_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:525" *) _083_;
  assign _127_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:525" *) _036_;
  assign _128_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:525" *) _037_;
  assign _129_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:525" *) _038_;
  assign _130_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:525" *) _039_;
  assign _131_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:526" *) _040_;
  assign _132_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:526" *) _084_;
  assign _133_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:526" *) _166_;
  assign _134_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:527" *) _085_;
  assign _135_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:527" *) _042_;
  assign _136_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:528" *) _086_;
  assign _137_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:528" *) _168_;
  assign _138_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:528" *) _087_;
  assign _139_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:529" *) _044_;
  assign _140_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:529" *) _045_;
  assign _141_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:529" *) _046_;
  assign _142_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:529" *) _047_;
  assign _143_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:529" *) _048_;
  assign _144_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:529" *) mantissa[0];
  assign _145_ = c_h_1_22 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:498" *) _088_;
  assign _146_ = c_h_1_13 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:500" *) _089_;
  assign _147_ = c_h_1_5 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:503" *) _093_;
  assign _148_ = c_h_1_12 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:504" *) _094_;
  assign _149_ = c_h_1_20 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:505" *) _097_;
  assign _150_ = _098_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:506" *) c_h_1_22;
  assign _151_ = IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_14_2_sdt_1 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:508" *) _058_;
  assign _152_ = IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_34_2_sdt_1 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:510" *) _061_;
  assign _153_ = IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_58_2_sdt_1 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:512" *) _064_;
  assign _154_ = IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_78_2_sdt_1 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:513" *) _067_;
  assign _155_ = IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_106_2_sdt_1 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:515" *) _070_;
  assign _156_ = IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_126_2_sdt_1 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:517" *) _073_;
  assign _157_ = _108_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:518" *) c_h_1_22;
  assign _158_ = mantissa[48] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:520" *) _110_;
  assign _159_ = mantissa[44] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:521" *) _112_;
  assign _160_ = mantissa[40] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:521" *) _114_;
  assign _161_ = mantissa[36] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:522" *) _116_;
  assign _162_ = mantissa[32] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:523" *) _120_;
  assign _163_ = mantissa[28] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:524" *) _122_;
  assign _164_ = mantissa[24] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:524" *) _124_;
  assign _165_ = mantissa[20] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:525" *) _126_;
  assign _166_ = mantissa[16] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:526" *) _132_;
  assign _167_ = mantissa[12] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:527" *) _134_;
  assign _168_ = mantissa[8] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:528" *) _136_;
  assign _169_ = mantissa[4] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:528" *) _138_;
  assign _170_ = _142_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:529" *) c_h_1_22;
  assign IntLeadZero_49U_leading_sign_49_0_rtn_IntLeadZero_49U_leading_sign_49_0_rtn_or_1_nl = _049_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:530" *) _051_;
  assign rtn = { c_h_1_23, IntLeadZero_49U_leading_sign_49_0_rtn_and_189_nl, IntLeadZero_49U_leading_sign_49_0_rtn_and_187_nl, IntLeadZero_49U_leading_sign_49_0_rtn_and_194_nl, IntLeadZero_49U_leading_sign_49_0_rtn_and_195_nl, IntLeadZero_49U_leading_sign_49_0_rtn_IntLeadZero_49U_leading_sign_49_0_rtn_or_1_nl };
endmodule
