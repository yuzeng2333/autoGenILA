module bar__DOT__i1(
__START__,
clk,
rst,
__ILA_bar_decode_of_i1__,
__ILA_bar_valid__,
data,
rst,
start,
timer,
__COUNTER_start__n0
);
input            __START__;
input            clk;
input            rst;
output            __ILA_bar_decode_of_i1__;
output            __ILA_bar_valid__;
output reg      [2:0] data;
output reg            rst;
output reg            start;
output reg      [2:0] timer;
output reg      [7:0] __COUNTER_start__n0;
wire            __ILA_bar_decode_of_i1__;
wire            __ILA_bar_valid__;
wire            __START__;
wire      [2:0] bv_3_0_n1;
wire      [2:0] bv_3_1_n78;
wire      [2:0] bv_3_6_n111;
wire      [2:0] bv_3_7_n3;
wire            clk;
(* keep *) wire      [2:0] data_randinit;
wire            n10;
wire            n100;
wire            n101;
wire      [2:0] n102;
wire      [2:0] n103;
wire            n104;
wire            n105;
wire            n106;
wire      [2:0] n107;
wire      [2:0] n108;
wire            n109;
wire      [2:0] n11;
wire            n110;
wire      [2:0] n112;
wire            n113;
wire      [2:0] n114;
wire      [2:0] n115;
wire      [2:0] n116;
wire      [2:0] n117;
wire      [2:0] n118;
wire            n119;
wire      [2:0] n12;
wire      [2:0] n120;
wire      [2:0] n121;
wire      [2:0] n122;
wire      [2:0] n123;
wire      [2:0] n124;
wire      [2:0] n125;
wire            n126;
wire      [2:0] n127;
wire      [2:0] n128;
wire      [2:0] n129;
wire      [2:0] n13;
wire      [2:0] n130;
wire      [2:0] n131;
wire      [2:0] n132;
wire            n133;
wire      [2:0] n134;
wire      [2:0] n135;
wire      [2:0] n136;
wire      [2:0] n137;
wire      [2:0] n138;
wire      [2:0] n139;
wire      [2:0] n14;
wire            n140;
wire      [2:0] n141;
wire      [2:0] n142;
wire      [2:0] n143;
wire      [2:0] n144;
wire      [2:0] n145;
wire      [2:0] n146;
wire            n147;
wire      [2:0] n148;
wire      [2:0] n149;
wire            n15;
wire      [2:0] n150;
wire      [2:0] n151;
wire      [2:0] n152;
wire      [2:0] n153;
wire            n154;
wire      [2:0] n155;
wire      [2:0] n156;
wire      [2:0] n157;
wire      [2:0] n158;
wire      [2:0] n159;
wire      [2:0] n16;
wire      [2:0] n17;
wire            n18;
wire            n19;
wire            n2;
wire      [2:0] n20;
wire      [2:0] n21;
wire            n22;
wire      [2:0] n23;
wire      [2:0] n24;
wire      [2:0] n25;
wire      [2:0] n26;
wire            n27;
wire      [2:0] n28;
wire      [2:0] n29;
wire            n30;
wire            n31;
wire      [2:0] n32;
wire      [2:0] n33;
wire            n34;
wire      [2:0] n35;
wire      [2:0] n36;
wire      [2:0] n37;
wire      [2:0] n38;
wire            n39;
wire      [2:0] n4;
wire      [2:0] n40;
wire      [2:0] n41;
wire            n42;
wire            n43;
wire      [2:0] n44;
wire      [2:0] n45;
wire            n46;
wire      [2:0] n47;
wire      [2:0] n48;
wire      [2:0] n49;
wire      [2:0] n5;
wire      [2:0] n50;
wire            n51;
wire      [2:0] n52;
wire      [2:0] n53;
wire            n54;
wire            n55;
wire      [2:0] n56;
wire      [2:0] n57;
wire            n58;
wire      [2:0] n59;
wire            n6;
wire      [2:0] n60;
wire      [2:0] n61;
wire      [2:0] n62;
wire            n63;
wire      [2:0] n64;
wire      [2:0] n65;
wire            n66;
wire            n67;
wire      [2:0] n68;
wire      [2:0] n69;
wire            n7;
wire            n70;
wire      [2:0] n71;
wire      [2:0] n72;
wire      [2:0] n73;
wire      [2:0] n74;
wire            n75;
wire      [2:0] n76;
wire      [2:0] n77;
wire            n79;
wire      [2:0] n8;
wire            n80;
wire            n81;
wire      [2:0] n82;
wire      [2:0] n83;
wire            n84;
wire            n85;
wire            n86;
wire      [2:0] n87;
wire      [2:0] n88;
wire            n89;
wire      [2:0] n9;
wire            n90;
wire            n91;
wire      [2:0] n92;
wire      [2:0] n93;
wire            n94;
wire            n95;
wire            n96;
wire      [2:0] n97;
wire      [2:0] n98;
wire            n99;
wire            rst;
(* keep *) wire            rst_randinit;
(* keep *) wire            start_randinit;
(* keep *) wire      [2:0] timer_randinit;
assign __ILA_bar_valid__ = 1'b1 ;
assign __ILA_bar_decode_of_i1__ = 1'b1 ;
assign bv_3_0_n1 = 3'h0 ;
assign n2 =  ( data ) == ( bv_3_0_n1 )  ;
assign bv_3_7_n3 = 3'h7 ;
assign n4 =  ( bv_3_7_n3 ) + ( data )  ;
assign n5 =  ( n2 ) ? ( data ) : ( n4 ) ;
assign n6 =  ( n5 ) == ( bv_3_0_n1 )  ;
assign n7 =  ( data ) == ( bv_3_0_n1 )  ;
assign n8 =  ( bv_3_7_n3 ) + ( data )  ;
assign n9 =  ( n7 ) ? ( data ) : ( n8 ) ;
assign n10 =  ( data ) == ( bv_3_0_n1 )  ;
assign n11 =  ( bv_3_7_n3 ) + ( data )  ;
assign n12 =  ( n10 ) ? ( data ) : ( n11 ) ;
assign n13 =  ( bv_3_7_n3 ) + ( n12 )  ;
assign n14 =  ( n6 ) ? ( n9 ) : ( n13 ) ;
assign n15 =  ( n14 ) == ( bv_3_0_n1 )  ;
assign n16 =  ( bv_3_7_n3 ) + ( n14 )  ;
assign n17 =  ( n15 ) ? ( n14 ) : ( n16 ) ;
assign n18 =  ( n17 ) == ( bv_3_0_n1 )  ;
assign n19 =  ( n14 ) == ( bv_3_0_n1 )  ;
assign n20 =  ( bv_3_7_n3 ) + ( n14 )  ;
assign n21 =  ( n19 ) ? ( n14 ) : ( n20 ) ;
assign n22 =  ( n14 ) == ( bv_3_0_n1 )  ;
assign n23 =  ( bv_3_7_n3 ) + ( n14 )  ;
assign n24 =  ( n22 ) ? ( n14 ) : ( n23 ) ;
assign n25 =  ( bv_3_7_n3 ) + ( n24 )  ;
assign n26 =  ( n18 ) ? ( n21 ) : ( n25 ) ;
assign n27 =  ( n26 ) == ( bv_3_0_n1 )  ;
assign n28 =  ( bv_3_7_n3 ) + ( n26 )  ;
assign n29 =  ( n27 ) ? ( n26 ) : ( n28 ) ;
assign n30 =  ( n29 ) == ( bv_3_0_n1 )  ;
assign n31 =  ( n26 ) == ( bv_3_0_n1 )  ;
assign n32 =  ( bv_3_7_n3 ) + ( n26 )  ;
assign n33 =  ( n31 ) ? ( n26 ) : ( n32 ) ;
assign n34 =  ( n26 ) == ( bv_3_0_n1 )  ;
assign n35 =  ( bv_3_7_n3 ) + ( n26 )  ;
assign n36 =  ( n34 ) ? ( n26 ) : ( n35 ) ;
assign n37 =  ( bv_3_7_n3 ) + ( n36 )  ;
assign n38 =  ( n30 ) ? ( n33 ) : ( n37 ) ;
assign n39 =  ( n38 ) == ( bv_3_0_n1 )  ;
assign n40 =  ( bv_3_7_n3 ) + ( n38 )  ;
assign n41 =  ( n39 ) ? ( n38 ) : ( n40 ) ;
assign n42 =  ( n41 ) == ( bv_3_0_n1 )  ;
assign n43 =  ( n38 ) == ( bv_3_0_n1 )  ;
assign n44 =  ( bv_3_7_n3 ) + ( n38 )  ;
assign n45 =  ( n43 ) ? ( n38 ) : ( n44 ) ;
assign n46 =  ( n38 ) == ( bv_3_0_n1 )  ;
assign n47 =  ( bv_3_7_n3 ) + ( n38 )  ;
assign n48 =  ( n46 ) ? ( n38 ) : ( n47 ) ;
assign n49 =  ( bv_3_7_n3 ) + ( n48 )  ;
assign n50 =  ( n42 ) ? ( n45 ) : ( n49 ) ;
assign n51 =  ( n50 ) == ( bv_3_0_n1 )  ;
assign n52 =  ( bv_3_7_n3 ) + ( n50 )  ;
assign n53 =  ( n51 ) ? ( n50 ) : ( n52 ) ;
assign n54 =  ( n53 ) == ( bv_3_0_n1 )  ;
assign n55 =  ( n50 ) == ( bv_3_0_n1 )  ;
assign n56 =  ( bv_3_7_n3 ) + ( n50 )  ;
assign n57 =  ( n55 ) ? ( n50 ) : ( n56 ) ;
assign n58 =  ( n50 ) == ( bv_3_0_n1 )  ;
assign n59 =  ( bv_3_7_n3 ) + ( n50 )  ;
assign n60 =  ( n58 ) ? ( n50 ) : ( n59 ) ;
assign n61 =  ( bv_3_7_n3 ) + ( n60 )  ;
assign n62 =  ( n54 ) ? ( n57 ) : ( n61 ) ;
assign n63 =  ( n62 ) == ( bv_3_0_n1 )  ;
assign n64 =  ( bv_3_7_n3 ) + ( n62 )  ;
assign n65 =  ( n63 ) ? ( n62 ) : ( n64 ) ;
assign n66 =  ( n65 ) == ( bv_3_0_n1 )  ;
assign n67 =  ( n62 ) == ( bv_3_0_n1 )  ;
assign n68 =  ( bv_3_7_n3 ) + ( n62 )  ;
assign n69 =  ( n67 ) ? ( n62 ) : ( n68 ) ;
assign n70 =  ( n62 ) == ( bv_3_0_n1 )  ;
assign n71 =  ( bv_3_7_n3 ) + ( n62 )  ;
assign n72 =  ( n70 ) ? ( n62 ) : ( n71 ) ;
assign n73 =  ( bv_3_7_n3 ) + ( n72 )  ;
assign n74 =  ( n66 ) ? ( n69 ) : ( n73 ) ;
assign n75 =  ( n74 ) == ( bv_3_0_n1 )  ;
assign n76 =  ( bv_3_7_n3 ) + ( n74 )  ;
assign n77 =  ( n75 ) ? ( n74 ) : ( n76 ) ;
assign bv_3_1_n78 = 3'h1 ;
assign n79 =  ( n77 ) == ( bv_3_1_n78 )  ;
assign n80 =  ( n74 ) == ( bv_3_1_n78 )  ;
assign n81 =  ( n62 ) == ( bv_3_0_n1 )  ;
assign n82 =  ( bv_3_7_n3 ) + ( n62 )  ;
assign n83 =  ( n81 ) ? ( n62 ) : ( n82 ) ;
assign n84 =  ( n83 ) == ( bv_3_1_n78 )  ;
assign n85 =  ( n62 ) == ( bv_3_1_n78 )  ;
assign n86 =  ( n50 ) == ( bv_3_0_n1 )  ;
assign n87 =  ( bv_3_7_n3 ) + ( n50 )  ;
assign n88 =  ( n86 ) ? ( n50 ) : ( n87 ) ;
assign n89 =  ( n88 ) == ( bv_3_1_n78 )  ;
assign n90 =  ( n50 ) == ( bv_3_1_n78 )  ;
assign n91 =  ( n38 ) == ( bv_3_0_n1 )  ;
assign n92 =  ( bv_3_7_n3 ) + ( n38 )  ;
assign n93 =  ( n91 ) ? ( n38 ) : ( n92 ) ;
assign n94 =  ( n93 ) == ( bv_3_1_n78 )  ;
assign n95 =  ( n38 ) == ( bv_3_1_n78 )  ;
assign n96 =  ( n26 ) == ( bv_3_0_n1 )  ;
assign n97 =  ( bv_3_7_n3 ) + ( n26 )  ;
assign n98 =  ( n96 ) ? ( n26 ) : ( n97 ) ;
assign n99 =  ( n98 ) == ( bv_3_1_n78 )  ;
assign n100 =  ( n26 ) == ( bv_3_1_n78 )  ;
assign n101 =  ( n14 ) == ( bv_3_0_n1 )  ;
assign n102 =  ( bv_3_7_n3 ) + ( n14 )  ;
assign n103 =  ( n101 ) ? ( n14 ) : ( n102 ) ;
assign n104 =  ( n103 ) == ( bv_3_1_n78 )  ;
assign n105 =  ( n14 ) == ( bv_3_1_n78 )  ;
assign n106 =  ( data ) == ( bv_3_0_n1 )  ;
assign n107 =  ( bv_3_7_n3 ) + ( data )  ;
assign n108 =  ( n106 ) ? ( data ) : ( n107 ) ;
assign n109 =  ( n108 ) == ( bv_3_1_n78 )  ;
assign n110 =  ( data ) == ( bv_3_1_n78 )  ;
assign bv_3_6_n111 = 3'h6 ;
assign n112 =  ( n110 ) ? ( bv_3_6_n111 ) : ( bv_3_7_n3 ) ;
assign n113 =  ( data ) == ( bv_3_1_n78 )  ;
assign n114 =  ( n113 ) ? ( bv_3_6_n111 ) : ( bv_3_7_n3 ) ;
assign n115 =  ( bv_3_1_n78 ) + ( n114 )  ;
assign n116 =  ( n109 ) ? ( n112 ) : ( n115 ) ;
assign n117 =  ( bv_3_1_n78 ) + ( n116 )  ;
assign n118 =  ( n105 ) ? ( n116 ) : ( n117 ) ;
assign n119 =  ( n14 ) == ( bv_3_1_n78 )  ;
assign n120 =  ( bv_3_1_n78 ) + ( n116 )  ;
assign n121 =  ( n119 ) ? ( n116 ) : ( n120 ) ;
assign n122 =  ( bv_3_1_n78 ) + ( n121 )  ;
assign n123 =  ( n104 ) ? ( n118 ) : ( n122 ) ;
assign n124 =  ( bv_3_1_n78 ) + ( n123 )  ;
assign n125 =  ( n100 ) ? ( n123 ) : ( n124 ) ;
assign n126 =  ( n26 ) == ( bv_3_1_n78 )  ;
assign n127 =  ( bv_3_1_n78 ) + ( n123 )  ;
assign n128 =  ( n126 ) ? ( n123 ) : ( n127 ) ;
assign n129 =  ( bv_3_1_n78 ) + ( n128 )  ;
assign n130 =  ( n99 ) ? ( n125 ) : ( n129 ) ;
assign n131 =  ( bv_3_1_n78 ) + ( n130 )  ;
assign n132 =  ( n95 ) ? ( n130 ) : ( n131 ) ;
assign n133 =  ( n38 ) == ( bv_3_1_n78 )  ;
assign n134 =  ( bv_3_1_n78 ) + ( n130 )  ;
assign n135 =  ( n133 ) ? ( n130 ) : ( n134 ) ;
assign n136 =  ( bv_3_1_n78 ) + ( n135 )  ;
assign n137 =  ( n94 ) ? ( n132 ) : ( n136 ) ;
assign n138 =  ( bv_3_1_n78 ) + ( n137 )  ;
assign n139 =  ( n90 ) ? ( n137 ) : ( n138 ) ;
assign n140 =  ( n50 ) == ( bv_3_1_n78 )  ;
assign n141 =  ( bv_3_1_n78 ) + ( n137 )  ;
assign n142 =  ( n140 ) ? ( n137 ) : ( n141 ) ;
assign n143 =  ( bv_3_1_n78 ) + ( n142 )  ;
assign n144 =  ( n89 ) ? ( n139 ) : ( n143 ) ;
assign n145 =  ( bv_3_1_n78 ) + ( n144 )  ;
assign n146 =  ( n85 ) ? ( n144 ) : ( n145 ) ;
assign n147 =  ( n62 ) == ( bv_3_1_n78 )  ;
assign n148 =  ( bv_3_1_n78 ) + ( n144 )  ;
assign n149 =  ( n147 ) ? ( n144 ) : ( n148 ) ;
assign n150 =  ( bv_3_1_n78 ) + ( n149 )  ;
assign n151 =  ( n84 ) ? ( n146 ) : ( n150 ) ;
assign n152 =  ( bv_3_1_n78 ) + ( n151 )  ;
assign n153 =  ( n80 ) ? ( n151 ) : ( n152 ) ;
assign n154 =  ( n74 ) == ( bv_3_1_n78 )  ;
assign n155 =  ( bv_3_1_n78 ) + ( n151 )  ;
assign n156 =  ( n154 ) ? ( n151 ) : ( n155 ) ;
assign n157 =  ( bv_3_1_n78 ) + ( n156 )  ;
assign n158 =  ( n79 ) ? ( n153 ) : ( n157 ) ;
assign n159 =  ( bv_3_0_n1 ) + ( n158 )  ;
always @(posedge clk) begin
   if(rst) begin
       data <= data_randinit ;
       rst <= rst_randinit ;
       start <= start_randinit ;
       timer <= timer_randinit ;
       __COUNTER_start__n0 <= 0;
   end
   else if(__START__ && __ILA_bar_valid__) begin
       if ( __ILA_bar_decode_of_i1__ ) begin 
           __COUNTER_start__n0 <= 1; end
       else if( (__COUNTER_start__n0 >= 1 ) && ( __COUNTER_start__n0 < 255 )) begin
           __COUNTER_start__n0 <= __COUNTER_start__n0 + 1; end
       if (__ILA_bar_decode_of_i1__) begin
           data <= data ;
       end
       if (__ILA_bar_decode_of_i1__) begin
           rst <= rst ;
       end
       if (__ILA_bar_decode_of_i1__) begin
           start <= start ;
       end
       if (__ILA_bar_decode_of_i1__) begin
           timer <= n159 ;
       end
   end
end
endmodule
