module bar__DOT__i1(
clk,
rst,
__ILA_bar_decode_of_i1__,
__ILA_bar_valid__,
in,
rcon,
out_1,
__COUNTER_start__n0
);
input            clk;
input            rst;
output            __ILA_bar_decode_of_i1__;
output            __ILA_bar_valid__;
output reg    [127:0] in;
output reg      [7:0] rcon;
output reg    [127:0] out_1;
output reg      [7:0] __COUNTER_start__n0;
wire            __ILA_bar_decode_of_i1__;
wire            __ILA_bar_valid__;
wire    [127:0] bv_128_0_n1;
wire      [7:0] bv_8_0_n583;
wire      [7:0] bv_8_100_n417;
wire      [7:0] bv_8_101_n261;
wire      [7:0] bv_8_102_n176;
wire      [7:0] bv_8_103_n525;
wire      [7:0] bv_8_104_n39;
wire      [7:0] bv_8_105_n113;
wire      [7:0] bv_8_106_n516;
wire      [7:0] bv_8_107_n513;
wire      [7:0] bv_8_108_n272;
wire      [7:0] bv_8_109_n289;
wire      [7:0] bv_8_10_n343;
wire      [7:0] bv_8_110_n504;
wire      [7:0] bv_8_111_n501;
wire      [7:0] bv_8_112_n188;
wire      [7:0] bv_8_113_n495;
wire      [7:0] bv_8_114_n491;
wire      [7:0] bv_8_115_n408;
wire      [7:0] bv_8_116_n211;
wire      [7:0] bv_8_117_n484;
wire      [7:0] bv_8_118_n480;
wire      [7:0] bv_8_119_n477;
wire      [7:0] bv_8_11_n359;
wire      [7:0] bv_8_120_n243;
wire      [7:0] bv_8_121_n302;
wire      [7:0] bv_8_122_n257;
wire      [7:0] bv_8_123_n467;
wire      [7:0] bv_8_124_n463;
wire      [7:0] bv_8_125_n460;
wire      [7:0] bv_8_126_n423;
wire      [7:0] bv_8_127_n455;
wire      [7:0] bv_8_128_n452;
wire      [7:0] bv_8_129_n401;
wire      [7:0] bv_8_12_n450;
wire      [7:0] bv_8_130_n445;
wire      [7:0] bv_8_131_n442;
wire      [7:0] bv_8_132_n438;
wire      [7:0] bv_8_133_n435;
wire      [7:0] bv_8_134_n142;
wire      [7:0] bv_8_135_n91;
wire      [7:0] bv_8_136_n381;
wire      [7:0] bv_8_137_n59;
wire      [7:0] bv_8_138_n192;
wire      [7:0] bv_8_139_n195;
wire      [7:0] bv_8_13_n55;
wire      [7:0] bv_8_140_n67;
wire      [7:0] bv_8_141_n285;
wire      [7:0] bv_8_142_n105;
wire      [7:0] bv_8_143_n406;
wire      [7:0] bv_8_144_n385;
wire      [7:0] bv_8_145_n312;
wire      [7:0] bv_8_146_n396;
wire      [7:0] bv_8_147_n393;
wire      [7:0] bv_8_148_n102;
wire      [7:0] bv_8_149_n308;
wire      [7:0] bv_8_14_n161;
wire      [7:0] bv_8_150_n383;
wire      [7:0] bv_8_151_n379;
wire      [7:0] bv_8_152_n121;
wire      [7:0] bv_8_153_n31;
wire      [7:0] bv_8_154_n371;
wire      [7:0] bv_8_155_n98;
wire      [7:0] bv_8_156_n365;
wire      [7:0] bv_8_157_n361;
wire      [7:0] bv_8_158_n130;
wire      [7:0] bv_8_159_n355;
wire      [7:0] bv_8_15_n23;
wire      [7:0] bv_8_160_n352;
wire      [7:0] bv_8_161_n63;
wire      [7:0] bv_8_162_n345;
wire      [7:0] bv_8_163_n341;
wire      [7:0] bv_8_164_n337;
wire      [7:0] bv_8_165_n333;
wire      [7:0] bv_8_166_n228;
wire      [7:0] bv_8_167_n326;
wire      [7:0] bv_8_168_n323;
wire      [7:0] bv_8_169_n276;
wire      [7:0] bv_8_16_n465;
wire      [7:0] bv_8_170_n318;
wire      [7:0] bv_8_171_n314;
wire      [7:0] bv_8_172_n310;
wire      [7:0] bv_8_173_n306;
wire      [7:0] bv_8_174_n254;
wire      [7:0] bv_8_175_n300;
wire      [7:0] bv_8_176_n19;
wire      [7:0] bv_8_177_n295;
wire      [7:0] bv_8_178_n291;
wire      [7:0] bv_8_179_n287;
wire      [7:0] bv_8_17_n117;
wire      [7:0] bv_8_180_n224;
wire      [7:0] bv_8_181_n180;
wire      [7:0] bv_8_182_n278;
wire      [7:0] bv_8_183_n274;
wire      [7:0] bv_8_184_n270;
wire      [7:0] bv_8_185_n146;
wire      [7:0] bv_8_186_n247;
wire      [7:0] bv_8_187_n11;
wire      [7:0] bv_8_188_n259;
wire      [7:0] bv_8_189_n199;
wire      [7:0] bv_8_18_n644;
wire      [7:0] bv_8_190_n252;
wire      [7:0] bv_8_191_n51;
wire      [7:0] bv_8_192_n245;
wire      [7:0] bv_8_193_n138;
wire      [7:0] bv_8_194_n238;
wire      [7:0] bv_8_195_n234;
wire      [7:0] bv_8_196_n230;
wire      [7:0] bv_8_197_n226;
wire      [7:0] bv_8_198_n221;
wire      [7:0] bv_8_199_n219;
wire      [7:0] bv_8_19_n447;
wire      [7:0] bv_8_1_n753;
wire      [7:0] bv_8_200_n216;
wire      [7:0] bv_8_201_n213;
wire      [7:0] bv_8_202_n209;
wire      [7:0] bv_8_203_n205;
wire      [7:0] bv_8_204_n201;
wire      [7:0] bv_8_205_n197;
wire      [7:0] bv_8_206_n83;
wire      [7:0] bv_8_207_n190;
wire      [7:0] bv_8_208_n186;
wire      [7:0] bv_8_209_n182;
wire      [7:0] bv_8_20_n369;
wire      [7:0] bv_8_210_n178;
wire      [7:0] bv_8_211_n174;
wire      [7:0] bv_8_212_n170;
wire      [7:0] bv_8_213_n166;
wire      [7:0] bv_8_214_n163;
wire      [7:0] bv_8_215_n159;
wire      [7:0] bv_8_216_n155;
wire      [7:0] bv_8_217_n109;
wire      [7:0] bv_8_218_n148;
wire      [7:0] bv_8_219_n144;
wire      [7:0] bv_8_21_n674;
wire      [7:0] bv_8_220_n140;
wire      [7:0] bv_8_221_n136;
wire      [7:0] bv_8_222_n132;
wire      [7:0] bv_8_223_n71;
wire      [7:0] bv_8_224_n126;
wire      [7:0] bv_8_225_n123;
wire      [7:0] bv_8_226_n119;
wire      [7:0] bv_8_227_n115;
wire      [7:0] bv_8_228_n111;
wire      [7:0] bv_8_229_n107;
wire      [7:0] bv_8_22_n7;
wire      [7:0] bv_8_230_n47;
wire      [7:0] bv_8_231_n100;
wire      [7:0] bv_8_232_n96;
wire      [7:0] bv_8_233_n87;
wire      [7:0] bv_8_234_n89;
wire      [7:0] bv_8_235_n85;
wire      [7:0] bv_8_236_n81;
wire      [7:0] bv_8_237_n77;
wire      [7:0] bv_8_238_n73;
wire      [7:0] bv_8_239_n69;
wire      [7:0] bv_8_23_n430;
wire      [7:0] bv_8_240_n65;
wire      [7:0] bv_8_241_n61;
wire      [7:0] bv_8_242_n57;
wire      [7:0] bv_8_243_n53;
wire      [7:0] bv_8_244_n49;
wire      [7:0] bv_8_245_n45;
wire      [7:0] bv_8_246_n41;
wire      [7:0] bv_8_247_n37;
wire      [7:0] bv_8_248_n33;
wire      [7:0] bv_8_249_n29;
wire      [7:0] bv_8_24_n659;
wire      [7:0] bv_8_250_n25;
wire      [7:0] bv_8_251_n21;
wire      [7:0] bv_8_252_n17;
wire      [7:0] bv_8_253_n13;
wire      [7:0] bv_8_254_n9;
wire      [7:0] bv_8_255_n5;
wire      [7:0] bv_8_25_n411;
wire      [7:0] bv_8_26_n619;
wire      [7:0] bv_8_27_n616;
wire      [7:0] bv_8_28_n232;
wire      [7:0] bv_8_29_n134;
wire      [7:0] bv_8_2_n518;
wire      [7:0] bv_8_30_n94;
wire      [7:0] bv_8_31_n207;
wire      [7:0] bv_8_32_n576;
wire      [7:0] bv_8_33_n469;
wire      [7:0] bv_8_34_n391;
wire      [7:0] bv_8_35_n664;
wire      [7:0] bv_8_36_n331;
wire      [7:0] bv_8_37_n240;
wire      [7:0] bv_8_38_n693;
wire      [7:0] bv_8_39_n635;
wire      [7:0] bv_8_3_n168;
wire      [7:0] bv_8_40_n75;
wire      [7:0] bv_8_41_n597;
wire      [7:0] bv_8_42_n388;
wire      [7:0] bv_8_43_n682;
wire      [7:0] bv_8_44_n622;
wire      [7:0] bv_8_45_n27;
wire      [7:0] bv_8_46_n236;
wire      [7:0] bv_8_47_n592;
wire      [7:0] bv_8_48_n669;
wire      [7:0] bv_8_49_n666;
wire      [7:0] bv_8_4_n671;
wire      [7:0] bv_8_50_n350;
wire      [7:0] bv_8_51_n529;
wire      [7:0] bv_8_52_n657;
wire      [7:0] bv_8_53_n153;
wire      [7:0] bv_8_54_n651;
wire      [7:0] bv_8_55_n293;
wire      [7:0] bv_8_56_n482;
wire      [7:0] bv_8_57_n559;
wire      [7:0] bv_8_58_n347;
wire      [7:0] bv_8_59_n604;
wire      [7:0] bv_8_5_n653;
wire      [7:0] bv_8_60_n508;
wire      [7:0] bv_8_61_n420;
wire      [7:0] bv_8_62_n184;
wire      [7:0] bv_8_63_n629;
wire      [7:0] bv_8_64_n493;
wire      [7:0] bv_8_65_n35;
wire      [7:0] bv_8_66_n43;
wire      [7:0] bv_8_67_n535;
wire      [7:0] bv_8_68_n433;
wire      [7:0] bv_8_69_n523;
wire      [7:0] bv_8_6_n335;
wire      [7:0] bv_8_70_n377;
wire      [7:0] bv_8_71_n608;
wire      [7:0] bv_8_72_n172;
wire      [7:0] bv_8_73_n339;
wire      [7:0] bv_8_74_n555;
wire      [7:0] bv_8_75_n203;
wire      [7:0] bv_8_76_n552;
wire      [7:0] bv_8_77_n532;
wire      [7:0] bv_8_78_n280;
wire      [7:0] bv_8_79_n398;
wire      [7:0] bv_8_7_n647;
wire      [7:0] bv_8_80_n511;
wire      [7:0] bv_8_81_n499;
wire      [7:0] bv_8_82_n581;
wire      [7:0] bv_8_83_n578;
wire      [7:0] bv_8_84_n15;
wire      [7:0] bv_8_85_n79;
wire      [7:0] bv_8_86_n268;
wire      [7:0] bv_8_87_n150;
wire      [7:0] bv_8_88_n549;
wire      [7:0] bv_8_89_n564;
wire      [7:0] bv_8_8_n250;
wire      [7:0] bv_8_90_n561;
wire      [7:0] bv_8_91_n557;
wire      [7:0] bv_8_92_n328;
wire      [7:0] bv_8_93_n414;
wire      [7:0] bv_8_94_n363;
wire      [7:0] bv_8_95_n440;
wire      [7:0] bv_8_96_n404;
wire      [7:0] bv_8_97_n157;
wire      [7:0] bv_8_98_n316;
wire      [7:0] bv_8_99_n537;
wire      [7:0] bv_8_9_n627;
wire            clk;
wire            n10;
wire      [7:0] n1000;
wire      [7:0] n1001;
wire      [7:0] n1002;
wire      [7:0] n1003;
wire      [7:0] n1004;
wire      [7:0] n1005;
wire      [7:0] n1006;
wire      [7:0] n1007;
wire      [7:0] n1008;
wire      [7:0] n1009;
wire            n101;
wire      [7:0] n1010;
wire      [7:0] n1011;
wire      [7:0] n1012;
wire      [7:0] n1013;
wire      [7:0] n1014;
wire      [7:0] n1015;
wire      [7:0] n1016;
wire      [7:0] n1017;
wire      [7:0] n1018;
wire      [7:0] n1019;
wire      [7:0] n1020;
wire      [7:0] n1021;
wire      [7:0] n1022;
wire      [7:0] n1023;
wire      [7:0] n1024;
wire      [7:0] n1025;
wire      [7:0] n1026;
wire      [7:0] n1027;
wire      [7:0] n1028;
wire      [7:0] n1029;
wire      [7:0] n103;
wire      [7:0] n1030;
wire            n1031;
wire      [7:0] n1032;
wire            n1033;
wire      [7:0] n1034;
wire            n1035;
wire      [7:0] n1036;
wire            n1037;
wire      [7:0] n1038;
wire            n1039;
wire            n104;
wire      [7:0] n1040;
wire            n1041;
wire      [7:0] n1042;
wire            n1043;
wire      [7:0] n1044;
wire            n1045;
wire      [7:0] n1046;
wire            n1047;
wire      [7:0] n1048;
wire            n1049;
wire      [7:0] n1050;
wire            n1051;
wire      [7:0] n1052;
wire            n1053;
wire      [7:0] n1054;
wire            n1055;
wire      [7:0] n1056;
wire            n1057;
wire      [7:0] n1058;
wire            n1059;
wire      [7:0] n106;
wire      [7:0] n1060;
wire            n1061;
wire      [7:0] n1062;
wire            n1063;
wire      [7:0] n1064;
wire            n1065;
wire      [7:0] n1066;
wire            n1067;
wire      [7:0] n1068;
wire            n1069;
wire      [7:0] n1070;
wire            n1071;
wire      [7:0] n1072;
wire            n1073;
wire      [7:0] n1074;
wire            n1075;
wire      [7:0] n1076;
wire            n1077;
wire      [7:0] n1078;
wire            n1079;
wire            n108;
wire      [7:0] n1080;
wire            n1081;
wire      [7:0] n1082;
wire            n1083;
wire      [7:0] n1084;
wire            n1085;
wire      [7:0] n1086;
wire            n1087;
wire      [7:0] n1088;
wire            n1089;
wire      [7:0] n1090;
wire            n1091;
wire      [7:0] n1092;
wire            n1093;
wire      [7:0] n1094;
wire            n1095;
wire      [7:0] n1096;
wire            n1097;
wire      [7:0] n1098;
wire            n1099;
wire      [7:0] n110;
wire      [7:0] n1100;
wire            n1101;
wire      [7:0] n1102;
wire            n1103;
wire      [7:0] n1104;
wire            n1105;
wire      [7:0] n1106;
wire            n1107;
wire      [7:0] n1108;
wire            n1109;
wire      [7:0] n1110;
wire            n1111;
wire      [7:0] n1112;
wire            n1113;
wire      [7:0] n1114;
wire            n1115;
wire      [7:0] n1116;
wire            n1117;
wire      [7:0] n1118;
wire            n1119;
wire            n112;
wire      [7:0] n1120;
wire            n1121;
wire      [7:0] n1122;
wire            n1123;
wire      [7:0] n1124;
wire            n1125;
wire      [7:0] n1126;
wire            n1127;
wire      [7:0] n1128;
wire            n1129;
wire      [7:0] n1130;
wire            n1131;
wire      [7:0] n1132;
wire            n1133;
wire      [7:0] n1134;
wire            n1135;
wire      [7:0] n1136;
wire            n1137;
wire      [7:0] n1138;
wire            n1139;
wire      [7:0] n114;
wire      [7:0] n1140;
wire            n1141;
wire      [7:0] n1142;
wire            n1143;
wire      [7:0] n1144;
wire            n1145;
wire      [7:0] n1146;
wire            n1147;
wire      [7:0] n1148;
wire            n1149;
wire      [7:0] n1150;
wire            n1151;
wire      [7:0] n1152;
wire            n1153;
wire      [7:0] n1154;
wire            n1155;
wire      [7:0] n1156;
wire            n1157;
wire      [7:0] n1158;
wire            n1159;
wire            n116;
wire      [7:0] n1160;
wire            n1161;
wire      [7:0] n1162;
wire            n1163;
wire      [7:0] n1164;
wire            n1165;
wire      [7:0] n1166;
wire            n1167;
wire      [7:0] n1168;
wire            n1169;
wire      [7:0] n1170;
wire            n1171;
wire      [7:0] n1172;
wire            n1173;
wire      [7:0] n1174;
wire            n1175;
wire      [7:0] n1176;
wire            n1177;
wire      [7:0] n1178;
wire            n1179;
wire      [7:0] n118;
wire      [7:0] n1180;
wire            n1181;
wire      [7:0] n1182;
wire            n1183;
wire      [7:0] n1184;
wire            n1185;
wire      [7:0] n1186;
wire            n1187;
wire      [7:0] n1188;
wire            n1189;
wire      [7:0] n1190;
wire            n1191;
wire      [7:0] n1192;
wire            n1193;
wire      [7:0] n1194;
wire            n1195;
wire      [7:0] n1196;
wire            n1197;
wire      [7:0] n1198;
wire            n1199;
wire      [7:0] n12;
wire            n120;
wire      [7:0] n1200;
wire            n1201;
wire      [7:0] n1202;
wire            n1203;
wire      [7:0] n1204;
wire            n1205;
wire      [7:0] n1206;
wire            n1207;
wire      [7:0] n1208;
wire            n1209;
wire      [7:0] n1210;
wire            n1211;
wire      [7:0] n1212;
wire            n1213;
wire      [7:0] n1214;
wire            n1215;
wire      [7:0] n1216;
wire            n1217;
wire      [7:0] n1218;
wire            n1219;
wire      [7:0] n122;
wire      [7:0] n1220;
wire            n1221;
wire      [7:0] n1222;
wire            n1223;
wire      [7:0] n1224;
wire            n1225;
wire      [7:0] n1226;
wire            n1227;
wire      [7:0] n1228;
wire            n1229;
wire      [7:0] n1230;
wire            n1231;
wire      [7:0] n1232;
wire            n1233;
wire      [7:0] n1234;
wire            n1235;
wire      [7:0] n1236;
wire            n1237;
wire      [7:0] n1238;
wire            n1239;
wire            n124;
wire      [7:0] n1240;
wire            n1241;
wire      [7:0] n1242;
wire            n1243;
wire      [7:0] n1244;
wire            n1245;
wire      [7:0] n1246;
wire            n1247;
wire      [7:0] n1248;
wire            n1249;
wire      [7:0] n125;
wire      [7:0] n1250;
wire            n1251;
wire      [7:0] n1252;
wire            n1253;
wire      [7:0] n1254;
wire            n1255;
wire      [7:0] n1256;
wire            n1257;
wire      [7:0] n1258;
wire            n1259;
wire      [7:0] n1260;
wire            n1261;
wire      [7:0] n1262;
wire            n1263;
wire      [7:0] n1264;
wire            n1265;
wire      [7:0] n1266;
wire            n1267;
wire      [7:0] n1268;
wire            n1269;
wire            n127;
wire      [7:0] n1270;
wire            n1271;
wire      [7:0] n1272;
wire            n1273;
wire      [7:0] n1274;
wire            n1275;
wire      [7:0] n1276;
wire            n1277;
wire      [7:0] n1278;
wire            n1279;
wire      [7:0] n128;
wire      [7:0] n1280;
wire            n1281;
wire      [7:0] n1282;
wire            n1283;
wire      [7:0] n1284;
wire            n1285;
wire      [7:0] n1286;
wire            n1287;
wire      [7:0] n1288;
wire            n1289;
wire            n129;
wire      [7:0] n1290;
wire            n1291;
wire      [7:0] n1292;
wire            n1293;
wire      [7:0] n1294;
wire            n1295;
wire      [7:0] n1296;
wire            n1297;
wire      [7:0] n1298;
wire            n1299;
wire      [7:0] n1300;
wire            n1301;
wire      [7:0] n1302;
wire            n1303;
wire      [7:0] n1304;
wire            n1305;
wire      [7:0] n1306;
wire            n1307;
wire      [7:0] n1308;
wire            n1309;
wire      [7:0] n131;
wire      [7:0] n1310;
wire            n1311;
wire      [7:0] n1312;
wire            n1313;
wire      [7:0] n1314;
wire            n1315;
wire      [7:0] n1316;
wire            n1317;
wire      [7:0] n1318;
wire            n1319;
wire      [7:0] n1320;
wire            n1321;
wire      [7:0] n1322;
wire            n1323;
wire      [7:0] n1324;
wire            n1325;
wire      [7:0] n1326;
wire            n1327;
wire      [7:0] n1328;
wire            n1329;
wire            n133;
wire      [7:0] n1330;
wire            n1331;
wire      [7:0] n1332;
wire            n1333;
wire      [7:0] n1334;
wire            n1335;
wire      [7:0] n1336;
wire            n1337;
wire      [7:0] n1338;
wire            n1339;
wire      [7:0] n1340;
wire            n1341;
wire      [7:0] n1342;
wire            n1343;
wire      [7:0] n1344;
wire            n1345;
wire      [7:0] n1346;
wire            n1347;
wire      [7:0] n1348;
wire            n1349;
wire      [7:0] n135;
wire      [7:0] n1350;
wire            n1351;
wire      [7:0] n1352;
wire            n1353;
wire      [7:0] n1354;
wire            n1355;
wire      [7:0] n1356;
wire            n1357;
wire      [7:0] n1358;
wire            n1359;
wire      [7:0] n1360;
wire            n1361;
wire      [7:0] n1362;
wire            n1363;
wire      [7:0] n1364;
wire            n1365;
wire      [7:0] n1366;
wire            n1367;
wire      [7:0] n1368;
wire            n1369;
wire            n137;
wire      [7:0] n1370;
wire            n1371;
wire      [7:0] n1372;
wire            n1373;
wire      [7:0] n1374;
wire            n1375;
wire      [7:0] n1376;
wire            n1377;
wire      [7:0] n1378;
wire            n1379;
wire      [7:0] n1380;
wire            n1381;
wire      [7:0] n1382;
wire            n1383;
wire      [7:0] n1384;
wire            n1385;
wire      [7:0] n1386;
wire            n1387;
wire      [7:0] n1388;
wire            n1389;
wire      [7:0] n139;
wire      [7:0] n1390;
wire            n1391;
wire      [7:0] n1392;
wire            n1393;
wire      [7:0] n1394;
wire            n1395;
wire      [7:0] n1396;
wire            n1397;
wire      [7:0] n1398;
wire            n1399;
wire            n14;
wire      [7:0] n1400;
wire            n1401;
wire      [7:0] n1402;
wire            n1403;
wire      [7:0] n1404;
wire            n1405;
wire      [7:0] n1406;
wire            n1407;
wire      [7:0] n1408;
wire            n1409;
wire            n141;
wire      [7:0] n1410;
wire            n1411;
wire      [7:0] n1412;
wire            n1413;
wire      [7:0] n1414;
wire            n1415;
wire      [7:0] n1416;
wire            n1417;
wire      [7:0] n1418;
wire            n1419;
wire      [7:0] n1420;
wire            n1421;
wire      [7:0] n1422;
wire            n1423;
wire      [7:0] n1424;
wire            n1425;
wire      [7:0] n1426;
wire            n1427;
wire      [7:0] n1428;
wire            n1429;
wire      [7:0] n143;
wire      [7:0] n1430;
wire            n1431;
wire      [7:0] n1432;
wire            n1433;
wire      [7:0] n1434;
wire            n1435;
wire      [7:0] n1436;
wire            n1437;
wire      [7:0] n1438;
wire            n1439;
wire      [7:0] n1440;
wire            n1441;
wire      [7:0] n1442;
wire            n1443;
wire      [7:0] n1444;
wire            n1445;
wire      [7:0] n1446;
wire            n1447;
wire      [7:0] n1448;
wire            n1449;
wire            n145;
wire      [7:0] n1450;
wire            n1451;
wire      [7:0] n1452;
wire            n1453;
wire      [7:0] n1454;
wire            n1455;
wire      [7:0] n1456;
wire            n1457;
wire      [7:0] n1458;
wire            n1459;
wire      [7:0] n1460;
wire            n1461;
wire      [7:0] n1462;
wire            n1463;
wire      [7:0] n1464;
wire            n1465;
wire      [7:0] n1466;
wire            n1467;
wire      [7:0] n1468;
wire            n1469;
wire      [7:0] n147;
wire      [7:0] n1470;
wire            n1471;
wire      [7:0] n1472;
wire            n1473;
wire      [7:0] n1474;
wire            n1475;
wire      [7:0] n1476;
wire            n1477;
wire      [7:0] n1478;
wire            n1479;
wire      [7:0] n1480;
wire            n1481;
wire      [7:0] n1482;
wire            n1483;
wire      [7:0] n1484;
wire            n1485;
wire      [7:0] n1486;
wire            n1487;
wire      [7:0] n1488;
wire            n1489;
wire            n149;
wire      [7:0] n1490;
wire            n1491;
wire      [7:0] n1492;
wire            n1493;
wire      [7:0] n1494;
wire            n1495;
wire      [7:0] n1496;
wire            n1497;
wire      [7:0] n1498;
wire            n1499;
wire      [7:0] n1500;
wire            n1501;
wire      [7:0] n1502;
wire            n1503;
wire      [7:0] n1504;
wire            n1505;
wire      [7:0] n1506;
wire            n1507;
wire      [7:0] n1508;
wire            n1509;
wire      [7:0] n151;
wire      [7:0] n1510;
wire            n1511;
wire      [7:0] n1512;
wire            n1513;
wire      [7:0] n1514;
wire            n1515;
wire      [7:0] n1516;
wire            n1517;
wire      [7:0] n1518;
wire            n1519;
wire            n152;
wire      [7:0] n1520;
wire            n1521;
wire      [7:0] n1522;
wire            n1523;
wire      [7:0] n1524;
wire            n1525;
wire      [7:0] n1526;
wire            n1527;
wire      [7:0] n1528;
wire            n1529;
wire      [7:0] n1530;
wire            n1531;
wire      [7:0] n1532;
wire            n1533;
wire      [7:0] n1534;
wire            n1535;
wire      [7:0] n1536;
wire            n1537;
wire      [7:0] n1538;
wire            n1539;
wire      [7:0] n154;
wire      [7:0] n1540;
wire            n1541;
wire      [7:0] n1542;
wire      [7:0] n1543;
wire      [7:0] n1544;
wire      [7:0] n1545;
wire      [7:0] n1546;
wire      [7:0] n1547;
wire      [7:0] n1548;
wire      [7:0] n1549;
wire      [7:0] n1550;
wire      [7:0] n1551;
wire      [7:0] n1552;
wire      [7:0] n1553;
wire      [7:0] n1554;
wire      [7:0] n1555;
wire      [7:0] n1556;
wire      [7:0] n1557;
wire      [7:0] n1558;
wire      [7:0] n1559;
wire            n156;
wire      [7:0] n1560;
wire      [7:0] n1561;
wire      [7:0] n1562;
wire      [7:0] n1563;
wire      [7:0] n1564;
wire      [7:0] n1565;
wire      [7:0] n1566;
wire      [7:0] n1567;
wire      [7:0] n1568;
wire      [7:0] n1569;
wire      [7:0] n1570;
wire      [7:0] n1571;
wire      [7:0] n1572;
wire      [7:0] n1573;
wire      [7:0] n1574;
wire      [7:0] n1575;
wire      [7:0] n1576;
wire      [7:0] n1577;
wire      [7:0] n1578;
wire      [7:0] n1579;
wire      [7:0] n158;
wire      [7:0] n1580;
wire      [7:0] n1581;
wire      [7:0] n1582;
wire      [7:0] n1583;
wire      [7:0] n1584;
wire      [7:0] n1585;
wire      [7:0] n1586;
wire      [7:0] n1587;
wire      [7:0] n1588;
wire      [7:0] n1589;
wire      [7:0] n1590;
wire      [7:0] n1591;
wire      [7:0] n1592;
wire      [7:0] n1593;
wire      [7:0] n1594;
wire      [7:0] n1595;
wire      [7:0] n1596;
wire      [7:0] n1597;
wire      [7:0] n1598;
wire      [7:0] n1599;
wire      [7:0] n16;
wire            n160;
wire      [7:0] n1600;
wire      [7:0] n1601;
wire      [7:0] n1602;
wire      [7:0] n1603;
wire      [7:0] n1604;
wire      [7:0] n1605;
wire      [7:0] n1606;
wire      [7:0] n1607;
wire      [7:0] n1608;
wire      [7:0] n1609;
wire      [7:0] n1610;
wire      [7:0] n1611;
wire      [7:0] n1612;
wire      [7:0] n1613;
wire      [7:0] n1614;
wire      [7:0] n1615;
wire      [7:0] n1616;
wire      [7:0] n1617;
wire      [7:0] n1618;
wire      [7:0] n1619;
wire      [7:0] n162;
wire      [7:0] n1620;
wire      [7:0] n1621;
wire      [7:0] n1622;
wire      [7:0] n1623;
wire      [7:0] n1624;
wire      [7:0] n1625;
wire      [7:0] n1626;
wire      [7:0] n1627;
wire      [7:0] n1628;
wire      [7:0] n1629;
wire      [7:0] n1630;
wire      [7:0] n1631;
wire      [7:0] n1632;
wire      [7:0] n1633;
wire      [7:0] n1634;
wire      [7:0] n1635;
wire      [7:0] n1636;
wire      [7:0] n1637;
wire      [7:0] n1638;
wire      [7:0] n1639;
wire            n164;
wire      [7:0] n1640;
wire      [7:0] n1641;
wire      [7:0] n1642;
wire      [7:0] n1643;
wire      [7:0] n1644;
wire      [7:0] n1645;
wire      [7:0] n1646;
wire      [7:0] n1647;
wire      [7:0] n1648;
wire      [7:0] n1649;
wire      [7:0] n165;
wire      [7:0] n1650;
wire      [7:0] n1651;
wire      [7:0] n1652;
wire      [7:0] n1653;
wire      [7:0] n1654;
wire      [7:0] n1655;
wire      [7:0] n1656;
wire      [7:0] n1657;
wire      [7:0] n1658;
wire      [7:0] n1659;
wire      [7:0] n1660;
wire      [7:0] n1661;
wire      [7:0] n1662;
wire      [7:0] n1663;
wire      [7:0] n1664;
wire      [7:0] n1665;
wire      [7:0] n1666;
wire      [7:0] n1667;
wire      [7:0] n1668;
wire      [7:0] n1669;
wire            n167;
wire      [7:0] n1670;
wire      [7:0] n1671;
wire      [7:0] n1672;
wire      [7:0] n1673;
wire      [7:0] n1674;
wire      [7:0] n1675;
wire      [7:0] n1676;
wire      [7:0] n1677;
wire      [7:0] n1678;
wire      [7:0] n1679;
wire      [7:0] n1680;
wire      [7:0] n1681;
wire      [7:0] n1682;
wire      [7:0] n1683;
wire      [7:0] n1684;
wire      [7:0] n1685;
wire      [7:0] n1686;
wire      [7:0] n1687;
wire      [7:0] n1688;
wire      [7:0] n1689;
wire      [7:0] n169;
wire      [7:0] n1690;
wire      [7:0] n1691;
wire      [7:0] n1692;
wire      [7:0] n1693;
wire      [7:0] n1694;
wire      [7:0] n1695;
wire      [7:0] n1696;
wire      [7:0] n1697;
wire      [7:0] n1698;
wire      [7:0] n1699;
wire      [7:0] n1700;
wire      [7:0] n1701;
wire      [7:0] n1702;
wire      [7:0] n1703;
wire      [7:0] n1704;
wire      [7:0] n1705;
wire      [7:0] n1706;
wire      [7:0] n1707;
wire      [7:0] n1708;
wire      [7:0] n1709;
wire            n171;
wire      [7:0] n1710;
wire      [7:0] n1711;
wire      [7:0] n1712;
wire      [7:0] n1713;
wire      [7:0] n1714;
wire      [7:0] n1715;
wire      [7:0] n1716;
wire      [7:0] n1717;
wire      [7:0] n1718;
wire      [7:0] n1719;
wire      [7:0] n1720;
wire      [7:0] n1721;
wire      [7:0] n1722;
wire      [7:0] n1723;
wire      [7:0] n1724;
wire      [7:0] n1725;
wire      [7:0] n1726;
wire      [7:0] n1727;
wire      [7:0] n1728;
wire      [7:0] n1729;
wire      [7:0] n173;
wire      [7:0] n1730;
wire      [7:0] n1731;
wire      [7:0] n1732;
wire      [7:0] n1733;
wire      [7:0] n1734;
wire      [7:0] n1735;
wire      [7:0] n1736;
wire      [7:0] n1737;
wire      [7:0] n1738;
wire      [7:0] n1739;
wire      [7:0] n1740;
wire      [7:0] n1741;
wire      [7:0] n1742;
wire      [7:0] n1743;
wire      [7:0] n1744;
wire      [7:0] n1745;
wire      [7:0] n1746;
wire      [7:0] n1747;
wire      [7:0] n1748;
wire      [7:0] n1749;
wire            n175;
wire      [7:0] n1750;
wire      [7:0] n1751;
wire      [7:0] n1752;
wire      [7:0] n1753;
wire      [7:0] n1754;
wire      [7:0] n1755;
wire      [7:0] n1756;
wire      [7:0] n1757;
wire      [7:0] n1758;
wire      [7:0] n1759;
wire      [7:0] n1760;
wire      [7:0] n1761;
wire      [7:0] n1762;
wire      [7:0] n1763;
wire      [7:0] n1764;
wire      [7:0] n1765;
wire      [7:0] n1766;
wire      [7:0] n1767;
wire      [7:0] n1768;
wire      [7:0] n1769;
wire      [7:0] n177;
wire      [7:0] n1770;
wire      [7:0] n1771;
wire      [7:0] n1772;
wire      [7:0] n1773;
wire      [7:0] n1774;
wire      [7:0] n1775;
wire      [7:0] n1776;
wire      [7:0] n1777;
wire      [7:0] n1778;
wire      [7:0] n1779;
wire      [7:0] n1780;
wire      [7:0] n1781;
wire      [7:0] n1782;
wire      [7:0] n1783;
wire      [7:0] n1784;
wire      [7:0] n1785;
wire      [7:0] n1786;
wire      [7:0] n1787;
wire      [7:0] n1788;
wire      [7:0] n1789;
wire            n179;
wire      [7:0] n1790;
wire      [7:0] n1791;
wire      [7:0] n1792;
wire      [7:0] n1793;
wire      [7:0] n1794;
wire      [7:0] n1795;
wire      [7:0] n1796;
wire      [7:0] n1797;
wire      [7:0] n1798;
wire     [15:0] n1799;
wire            n18;
wire      [7:0] n1800;
wire      [7:0] n1801;
wire            n1802;
wire      [7:0] n1803;
wire            n1804;
wire      [7:0] n1805;
wire            n1806;
wire      [7:0] n1807;
wire            n1808;
wire      [7:0] n1809;
wire      [7:0] n181;
wire            n1810;
wire      [7:0] n1811;
wire            n1812;
wire      [7:0] n1813;
wire            n1814;
wire      [7:0] n1815;
wire            n1816;
wire      [7:0] n1817;
wire            n1818;
wire      [7:0] n1819;
wire            n1820;
wire      [7:0] n1821;
wire            n1822;
wire      [7:0] n1823;
wire            n1824;
wire      [7:0] n1825;
wire            n1826;
wire      [7:0] n1827;
wire            n1828;
wire      [7:0] n1829;
wire            n183;
wire            n1830;
wire      [7:0] n1831;
wire            n1832;
wire      [7:0] n1833;
wire            n1834;
wire      [7:0] n1835;
wire            n1836;
wire      [7:0] n1837;
wire            n1838;
wire      [7:0] n1839;
wire            n1840;
wire      [7:0] n1841;
wire            n1842;
wire      [7:0] n1843;
wire            n1844;
wire      [7:0] n1845;
wire            n1846;
wire      [7:0] n1847;
wire            n1848;
wire      [7:0] n1849;
wire      [7:0] n185;
wire            n1850;
wire      [7:0] n1851;
wire            n1852;
wire      [7:0] n1853;
wire            n1854;
wire      [7:0] n1855;
wire            n1856;
wire      [7:0] n1857;
wire            n1858;
wire      [7:0] n1859;
wire            n1860;
wire      [7:0] n1861;
wire            n1862;
wire      [7:0] n1863;
wire            n1864;
wire      [7:0] n1865;
wire            n1866;
wire      [7:0] n1867;
wire            n1868;
wire      [7:0] n1869;
wire            n187;
wire            n1870;
wire      [7:0] n1871;
wire            n1872;
wire      [7:0] n1873;
wire            n1874;
wire      [7:0] n1875;
wire            n1876;
wire      [7:0] n1877;
wire            n1878;
wire      [7:0] n1879;
wire            n1880;
wire      [7:0] n1881;
wire            n1882;
wire      [7:0] n1883;
wire            n1884;
wire      [7:0] n1885;
wire            n1886;
wire      [7:0] n1887;
wire            n1888;
wire      [7:0] n1889;
wire      [7:0] n189;
wire            n1890;
wire      [7:0] n1891;
wire            n1892;
wire      [7:0] n1893;
wire            n1894;
wire      [7:0] n1895;
wire            n1896;
wire      [7:0] n1897;
wire            n1898;
wire      [7:0] n1899;
wire            n1900;
wire      [7:0] n1901;
wire            n1902;
wire      [7:0] n1903;
wire            n1904;
wire      [7:0] n1905;
wire            n1906;
wire      [7:0] n1907;
wire            n1908;
wire      [7:0] n1909;
wire            n191;
wire            n1910;
wire      [7:0] n1911;
wire            n1912;
wire      [7:0] n1913;
wire            n1914;
wire      [7:0] n1915;
wire            n1916;
wire      [7:0] n1917;
wire            n1918;
wire      [7:0] n1919;
wire            n1920;
wire      [7:0] n1921;
wire            n1922;
wire      [7:0] n1923;
wire            n1924;
wire      [7:0] n1925;
wire            n1926;
wire      [7:0] n1927;
wire            n1928;
wire      [7:0] n1929;
wire      [7:0] n193;
wire            n1930;
wire      [7:0] n1931;
wire            n1932;
wire      [7:0] n1933;
wire            n1934;
wire      [7:0] n1935;
wire            n1936;
wire      [7:0] n1937;
wire            n1938;
wire      [7:0] n1939;
wire            n194;
wire            n1940;
wire      [7:0] n1941;
wire            n1942;
wire      [7:0] n1943;
wire            n1944;
wire      [7:0] n1945;
wire            n1946;
wire      [7:0] n1947;
wire            n1948;
wire      [7:0] n1949;
wire            n1950;
wire      [7:0] n1951;
wire            n1952;
wire      [7:0] n1953;
wire            n1954;
wire      [7:0] n1955;
wire            n1956;
wire      [7:0] n1957;
wire            n1958;
wire      [7:0] n1959;
wire      [7:0] n196;
wire            n1960;
wire      [7:0] n1961;
wire            n1962;
wire      [7:0] n1963;
wire            n1964;
wire      [7:0] n1965;
wire            n1966;
wire      [7:0] n1967;
wire            n1968;
wire      [7:0] n1969;
wire            n1970;
wire      [7:0] n1971;
wire            n1972;
wire      [7:0] n1973;
wire            n1974;
wire      [7:0] n1975;
wire            n1976;
wire      [7:0] n1977;
wire            n1978;
wire      [7:0] n1979;
wire            n198;
wire            n1980;
wire      [7:0] n1981;
wire            n1982;
wire      [7:0] n1983;
wire            n1984;
wire      [7:0] n1985;
wire            n1986;
wire      [7:0] n1987;
wire            n1988;
wire      [7:0] n1989;
wire            n1990;
wire      [7:0] n1991;
wire            n1992;
wire      [7:0] n1993;
wire            n1994;
wire      [7:0] n1995;
wire            n1996;
wire      [7:0] n1997;
wire            n1998;
wire      [7:0] n1999;
wire      [7:0] n2;
wire      [7:0] n20;
wire      [7:0] n200;
wire            n2000;
wire      [7:0] n2001;
wire            n2002;
wire      [7:0] n2003;
wire            n2004;
wire      [7:0] n2005;
wire            n2006;
wire      [7:0] n2007;
wire            n2008;
wire      [7:0] n2009;
wire            n2010;
wire      [7:0] n2011;
wire            n2012;
wire      [7:0] n2013;
wire            n2014;
wire      [7:0] n2015;
wire            n2016;
wire      [7:0] n2017;
wire            n2018;
wire      [7:0] n2019;
wire            n202;
wire            n2020;
wire      [7:0] n2021;
wire            n2022;
wire      [7:0] n2023;
wire            n2024;
wire      [7:0] n2025;
wire            n2026;
wire      [7:0] n2027;
wire            n2028;
wire      [7:0] n2029;
wire            n2030;
wire      [7:0] n2031;
wire            n2032;
wire      [7:0] n2033;
wire            n2034;
wire      [7:0] n2035;
wire            n2036;
wire      [7:0] n2037;
wire            n2038;
wire      [7:0] n2039;
wire      [7:0] n204;
wire            n2040;
wire      [7:0] n2041;
wire            n2042;
wire      [7:0] n2043;
wire            n2044;
wire      [7:0] n2045;
wire            n2046;
wire      [7:0] n2047;
wire            n2048;
wire      [7:0] n2049;
wire            n2050;
wire      [7:0] n2051;
wire            n2052;
wire      [7:0] n2053;
wire            n2054;
wire      [7:0] n2055;
wire            n2056;
wire      [7:0] n2057;
wire            n2058;
wire      [7:0] n2059;
wire            n206;
wire            n2060;
wire      [7:0] n2061;
wire            n2062;
wire      [7:0] n2063;
wire            n2064;
wire      [7:0] n2065;
wire            n2066;
wire      [7:0] n2067;
wire            n2068;
wire      [7:0] n2069;
wire            n2070;
wire      [7:0] n2071;
wire            n2072;
wire      [7:0] n2073;
wire            n2074;
wire      [7:0] n2075;
wire            n2076;
wire      [7:0] n2077;
wire            n2078;
wire      [7:0] n2079;
wire      [7:0] n208;
wire            n2080;
wire      [7:0] n2081;
wire            n2082;
wire      [7:0] n2083;
wire            n2084;
wire      [7:0] n2085;
wire            n2086;
wire      [7:0] n2087;
wire            n2088;
wire      [7:0] n2089;
wire            n2090;
wire      [7:0] n2091;
wire            n2092;
wire      [7:0] n2093;
wire            n2094;
wire      [7:0] n2095;
wire            n2096;
wire      [7:0] n2097;
wire            n2098;
wire      [7:0] n2099;
wire            n210;
wire            n2100;
wire      [7:0] n2101;
wire            n2102;
wire      [7:0] n2103;
wire            n2104;
wire      [7:0] n2105;
wire            n2106;
wire      [7:0] n2107;
wire            n2108;
wire      [7:0] n2109;
wire            n2110;
wire      [7:0] n2111;
wire            n2112;
wire      [7:0] n2113;
wire            n2114;
wire      [7:0] n2115;
wire            n2116;
wire      [7:0] n2117;
wire            n2118;
wire      [7:0] n2119;
wire      [7:0] n212;
wire            n2120;
wire      [7:0] n2121;
wire            n2122;
wire      [7:0] n2123;
wire            n2124;
wire      [7:0] n2125;
wire            n2126;
wire      [7:0] n2127;
wire            n2128;
wire      [7:0] n2129;
wire            n2130;
wire      [7:0] n2131;
wire            n2132;
wire      [7:0] n2133;
wire            n2134;
wire      [7:0] n2135;
wire            n2136;
wire      [7:0] n2137;
wire            n2138;
wire      [7:0] n2139;
wire            n214;
wire            n2140;
wire      [7:0] n2141;
wire            n2142;
wire      [7:0] n2143;
wire            n2144;
wire      [7:0] n2145;
wire            n2146;
wire      [7:0] n2147;
wire            n2148;
wire      [7:0] n2149;
wire      [7:0] n215;
wire            n2150;
wire      [7:0] n2151;
wire            n2152;
wire      [7:0] n2153;
wire            n2154;
wire      [7:0] n2155;
wire            n2156;
wire      [7:0] n2157;
wire            n2158;
wire      [7:0] n2159;
wire            n2160;
wire      [7:0] n2161;
wire            n2162;
wire      [7:0] n2163;
wire            n2164;
wire      [7:0] n2165;
wire            n2166;
wire      [7:0] n2167;
wire            n2168;
wire      [7:0] n2169;
wire            n217;
wire            n2170;
wire      [7:0] n2171;
wire            n2172;
wire      [7:0] n2173;
wire            n2174;
wire      [7:0] n2175;
wire            n2176;
wire      [7:0] n2177;
wire            n2178;
wire      [7:0] n2179;
wire      [7:0] n218;
wire            n2180;
wire      [7:0] n2181;
wire            n2182;
wire      [7:0] n2183;
wire            n2184;
wire      [7:0] n2185;
wire            n2186;
wire      [7:0] n2187;
wire            n2188;
wire      [7:0] n2189;
wire            n2190;
wire      [7:0] n2191;
wire            n2192;
wire      [7:0] n2193;
wire            n2194;
wire      [7:0] n2195;
wire            n2196;
wire      [7:0] n2197;
wire            n2198;
wire      [7:0] n2199;
wire            n22;
wire            n220;
wire            n2200;
wire      [7:0] n2201;
wire            n2202;
wire      [7:0] n2203;
wire            n2204;
wire      [7:0] n2205;
wire            n2206;
wire      [7:0] n2207;
wire            n2208;
wire      [7:0] n2209;
wire            n2210;
wire      [7:0] n2211;
wire            n2212;
wire      [7:0] n2213;
wire            n2214;
wire      [7:0] n2215;
wire            n2216;
wire      [7:0] n2217;
wire            n2218;
wire      [7:0] n2219;
wire      [7:0] n222;
wire            n2220;
wire      [7:0] n2221;
wire            n2222;
wire      [7:0] n2223;
wire            n2224;
wire      [7:0] n2225;
wire            n2226;
wire      [7:0] n2227;
wire            n2228;
wire      [7:0] n2229;
wire            n223;
wire            n2230;
wire      [7:0] n2231;
wire            n2232;
wire      [7:0] n2233;
wire            n2234;
wire      [7:0] n2235;
wire            n2236;
wire      [7:0] n2237;
wire            n2238;
wire      [7:0] n2239;
wire            n2240;
wire      [7:0] n2241;
wire            n2242;
wire      [7:0] n2243;
wire            n2244;
wire      [7:0] n2245;
wire            n2246;
wire      [7:0] n2247;
wire            n2248;
wire      [7:0] n2249;
wire      [7:0] n225;
wire            n2250;
wire      [7:0] n2251;
wire            n2252;
wire      [7:0] n2253;
wire            n2254;
wire      [7:0] n2255;
wire            n2256;
wire      [7:0] n2257;
wire            n2258;
wire      [7:0] n2259;
wire            n2260;
wire      [7:0] n2261;
wire            n2262;
wire      [7:0] n2263;
wire            n2264;
wire      [7:0] n2265;
wire            n2266;
wire      [7:0] n2267;
wire            n2268;
wire      [7:0] n2269;
wire            n227;
wire            n2270;
wire      [7:0] n2271;
wire            n2272;
wire      [7:0] n2273;
wire            n2274;
wire      [7:0] n2275;
wire            n2276;
wire      [7:0] n2277;
wire            n2278;
wire      [7:0] n2279;
wire            n2280;
wire      [7:0] n2281;
wire            n2282;
wire      [7:0] n2283;
wire            n2284;
wire      [7:0] n2285;
wire            n2286;
wire      [7:0] n2287;
wire            n2288;
wire      [7:0] n2289;
wire      [7:0] n229;
wire            n2290;
wire      [7:0] n2291;
wire            n2292;
wire      [7:0] n2293;
wire            n2294;
wire      [7:0] n2295;
wire            n2296;
wire      [7:0] n2297;
wire            n2298;
wire      [7:0] n2299;
wire            n2300;
wire      [7:0] n2301;
wire            n2302;
wire      [7:0] n2303;
wire            n2304;
wire      [7:0] n2305;
wire            n2306;
wire      [7:0] n2307;
wire            n2308;
wire      [7:0] n2309;
wire            n231;
wire            n2310;
wire      [7:0] n2311;
wire            n2312;
wire      [7:0] n2313;
wire      [7:0] n2314;
wire      [7:0] n2315;
wire      [7:0] n2316;
wire      [7:0] n2317;
wire      [7:0] n2318;
wire      [7:0] n2319;
wire      [7:0] n2320;
wire      [7:0] n2321;
wire      [7:0] n2322;
wire      [7:0] n2323;
wire      [7:0] n2324;
wire      [7:0] n2325;
wire      [7:0] n2326;
wire      [7:0] n2327;
wire      [7:0] n2328;
wire      [7:0] n2329;
wire      [7:0] n233;
wire      [7:0] n2330;
wire      [7:0] n2331;
wire      [7:0] n2332;
wire      [7:0] n2333;
wire      [7:0] n2334;
wire      [7:0] n2335;
wire      [7:0] n2336;
wire      [7:0] n2337;
wire      [7:0] n2338;
wire      [7:0] n2339;
wire      [7:0] n2340;
wire      [7:0] n2341;
wire      [7:0] n2342;
wire      [7:0] n2343;
wire      [7:0] n2344;
wire      [7:0] n2345;
wire      [7:0] n2346;
wire      [7:0] n2347;
wire      [7:0] n2348;
wire      [7:0] n2349;
wire            n235;
wire      [7:0] n2350;
wire      [7:0] n2351;
wire      [7:0] n2352;
wire      [7:0] n2353;
wire      [7:0] n2354;
wire      [7:0] n2355;
wire      [7:0] n2356;
wire      [7:0] n2357;
wire      [7:0] n2358;
wire      [7:0] n2359;
wire      [7:0] n2360;
wire      [7:0] n2361;
wire      [7:0] n2362;
wire      [7:0] n2363;
wire      [7:0] n2364;
wire      [7:0] n2365;
wire      [7:0] n2366;
wire      [7:0] n2367;
wire      [7:0] n2368;
wire      [7:0] n2369;
wire      [7:0] n237;
wire      [7:0] n2370;
wire      [7:0] n2371;
wire      [7:0] n2372;
wire      [7:0] n2373;
wire      [7:0] n2374;
wire      [7:0] n2375;
wire      [7:0] n2376;
wire      [7:0] n2377;
wire      [7:0] n2378;
wire      [7:0] n2379;
wire      [7:0] n2380;
wire      [7:0] n2381;
wire      [7:0] n2382;
wire      [7:0] n2383;
wire      [7:0] n2384;
wire      [7:0] n2385;
wire      [7:0] n2386;
wire      [7:0] n2387;
wire      [7:0] n2388;
wire      [7:0] n2389;
wire            n239;
wire      [7:0] n2390;
wire      [7:0] n2391;
wire      [7:0] n2392;
wire      [7:0] n2393;
wire      [7:0] n2394;
wire      [7:0] n2395;
wire      [7:0] n2396;
wire      [7:0] n2397;
wire      [7:0] n2398;
wire      [7:0] n2399;
wire      [7:0] n24;
wire      [7:0] n2400;
wire      [7:0] n2401;
wire      [7:0] n2402;
wire      [7:0] n2403;
wire      [7:0] n2404;
wire      [7:0] n2405;
wire      [7:0] n2406;
wire      [7:0] n2407;
wire      [7:0] n2408;
wire      [7:0] n2409;
wire      [7:0] n241;
wire      [7:0] n2410;
wire      [7:0] n2411;
wire      [7:0] n2412;
wire      [7:0] n2413;
wire      [7:0] n2414;
wire      [7:0] n2415;
wire      [7:0] n2416;
wire      [7:0] n2417;
wire      [7:0] n2418;
wire      [7:0] n2419;
wire            n242;
wire      [7:0] n2420;
wire      [7:0] n2421;
wire      [7:0] n2422;
wire      [7:0] n2423;
wire      [7:0] n2424;
wire      [7:0] n2425;
wire      [7:0] n2426;
wire      [7:0] n2427;
wire      [7:0] n2428;
wire      [7:0] n2429;
wire      [7:0] n2430;
wire      [7:0] n2431;
wire      [7:0] n2432;
wire      [7:0] n2433;
wire      [7:0] n2434;
wire      [7:0] n2435;
wire      [7:0] n2436;
wire      [7:0] n2437;
wire      [7:0] n2438;
wire      [7:0] n2439;
wire      [7:0] n244;
wire      [7:0] n2440;
wire      [7:0] n2441;
wire      [7:0] n2442;
wire      [7:0] n2443;
wire      [7:0] n2444;
wire      [7:0] n2445;
wire      [7:0] n2446;
wire      [7:0] n2447;
wire      [7:0] n2448;
wire      [7:0] n2449;
wire      [7:0] n2450;
wire      [7:0] n2451;
wire      [7:0] n2452;
wire      [7:0] n2453;
wire      [7:0] n2454;
wire      [7:0] n2455;
wire      [7:0] n2456;
wire      [7:0] n2457;
wire      [7:0] n2458;
wire      [7:0] n2459;
wire            n246;
wire      [7:0] n2460;
wire      [7:0] n2461;
wire      [7:0] n2462;
wire      [7:0] n2463;
wire      [7:0] n2464;
wire      [7:0] n2465;
wire      [7:0] n2466;
wire      [7:0] n2467;
wire      [7:0] n2468;
wire      [7:0] n2469;
wire      [7:0] n2470;
wire      [7:0] n2471;
wire      [7:0] n2472;
wire      [7:0] n2473;
wire      [7:0] n2474;
wire      [7:0] n2475;
wire      [7:0] n2476;
wire      [7:0] n2477;
wire      [7:0] n2478;
wire      [7:0] n2479;
wire      [7:0] n248;
wire      [7:0] n2480;
wire      [7:0] n2481;
wire      [7:0] n2482;
wire      [7:0] n2483;
wire      [7:0] n2484;
wire      [7:0] n2485;
wire      [7:0] n2486;
wire      [7:0] n2487;
wire      [7:0] n2488;
wire      [7:0] n2489;
wire            n249;
wire      [7:0] n2490;
wire      [7:0] n2491;
wire      [7:0] n2492;
wire      [7:0] n2493;
wire      [7:0] n2494;
wire      [7:0] n2495;
wire      [7:0] n2496;
wire      [7:0] n2497;
wire      [7:0] n2498;
wire      [7:0] n2499;
wire      [7:0] n2500;
wire      [7:0] n2501;
wire      [7:0] n2502;
wire      [7:0] n2503;
wire      [7:0] n2504;
wire      [7:0] n2505;
wire      [7:0] n2506;
wire      [7:0] n2507;
wire      [7:0] n2508;
wire      [7:0] n2509;
wire      [7:0] n251;
wire      [7:0] n2510;
wire      [7:0] n2511;
wire      [7:0] n2512;
wire      [7:0] n2513;
wire      [7:0] n2514;
wire      [7:0] n2515;
wire      [7:0] n2516;
wire      [7:0] n2517;
wire      [7:0] n2518;
wire      [7:0] n2519;
wire      [7:0] n2520;
wire      [7:0] n2521;
wire      [7:0] n2522;
wire      [7:0] n2523;
wire      [7:0] n2524;
wire      [7:0] n2525;
wire      [7:0] n2526;
wire      [7:0] n2527;
wire      [7:0] n2528;
wire      [7:0] n2529;
wire            n253;
wire      [7:0] n2530;
wire      [7:0] n2531;
wire      [7:0] n2532;
wire      [7:0] n2533;
wire      [7:0] n2534;
wire      [7:0] n2535;
wire      [7:0] n2536;
wire      [7:0] n2537;
wire      [7:0] n2538;
wire      [7:0] n2539;
wire      [7:0] n2540;
wire      [7:0] n2541;
wire      [7:0] n2542;
wire      [7:0] n2543;
wire      [7:0] n2544;
wire      [7:0] n2545;
wire      [7:0] n2546;
wire      [7:0] n2547;
wire      [7:0] n2548;
wire      [7:0] n2549;
wire      [7:0] n255;
wire      [7:0] n2550;
wire      [7:0] n2551;
wire      [7:0] n2552;
wire      [7:0] n2553;
wire      [7:0] n2554;
wire      [7:0] n2555;
wire      [7:0] n2556;
wire      [7:0] n2557;
wire      [7:0] n2558;
wire      [7:0] n2559;
wire            n256;
wire      [7:0] n2560;
wire      [7:0] n2561;
wire      [7:0] n2562;
wire      [7:0] n2563;
wire      [7:0] n2564;
wire      [7:0] n2565;
wire      [7:0] n2566;
wire      [7:0] n2567;
wire      [7:0] n2568;
wire      [7:0] n2569;
wire     [23:0] n2570;
wire      [7:0] n2571;
wire      [7:0] n2572;
wire            n2573;
wire      [7:0] n2574;
wire            n2575;
wire      [7:0] n2576;
wire            n2577;
wire      [7:0] n2578;
wire            n2579;
wire      [7:0] n258;
wire      [7:0] n2580;
wire            n2581;
wire      [7:0] n2582;
wire            n2583;
wire      [7:0] n2584;
wire            n2585;
wire      [7:0] n2586;
wire            n2587;
wire      [7:0] n2588;
wire            n2589;
wire      [7:0] n2590;
wire            n2591;
wire      [7:0] n2592;
wire            n2593;
wire      [7:0] n2594;
wire            n2595;
wire      [7:0] n2596;
wire            n2597;
wire      [7:0] n2598;
wire            n2599;
wire            n26;
wire            n260;
wire      [7:0] n2600;
wire            n2601;
wire      [7:0] n2602;
wire            n2603;
wire      [7:0] n2604;
wire            n2605;
wire      [7:0] n2606;
wire            n2607;
wire      [7:0] n2608;
wire            n2609;
wire      [7:0] n2610;
wire            n2611;
wire      [7:0] n2612;
wire            n2613;
wire      [7:0] n2614;
wire            n2615;
wire      [7:0] n2616;
wire            n2617;
wire      [7:0] n2618;
wire            n2619;
wire      [7:0] n262;
wire      [7:0] n2620;
wire            n2621;
wire      [7:0] n2622;
wire            n2623;
wire      [7:0] n2624;
wire            n2625;
wire      [7:0] n2626;
wire            n2627;
wire      [7:0] n2628;
wire            n2629;
wire            n263;
wire      [7:0] n2630;
wire            n2631;
wire      [7:0] n2632;
wire            n2633;
wire      [7:0] n2634;
wire            n2635;
wire      [7:0] n2636;
wire            n2637;
wire      [7:0] n2638;
wire            n2639;
wire      [7:0] n264;
wire      [7:0] n2640;
wire            n2641;
wire      [7:0] n2642;
wire            n2643;
wire      [7:0] n2644;
wire            n2645;
wire      [7:0] n2646;
wire            n2647;
wire      [7:0] n2648;
wire            n2649;
wire            n265;
wire      [7:0] n2650;
wire            n2651;
wire      [7:0] n2652;
wire            n2653;
wire      [7:0] n2654;
wire            n2655;
wire      [7:0] n2656;
wire            n2657;
wire      [7:0] n2658;
wire            n2659;
wire      [7:0] n266;
wire      [7:0] n2660;
wire            n2661;
wire      [7:0] n2662;
wire            n2663;
wire      [7:0] n2664;
wire            n2665;
wire      [7:0] n2666;
wire            n2667;
wire      [7:0] n2668;
wire            n2669;
wire            n267;
wire      [7:0] n2670;
wire            n2671;
wire      [7:0] n2672;
wire            n2673;
wire      [7:0] n2674;
wire            n2675;
wire      [7:0] n2676;
wire            n2677;
wire      [7:0] n2678;
wire            n2679;
wire      [7:0] n2680;
wire            n2681;
wire      [7:0] n2682;
wire            n2683;
wire      [7:0] n2684;
wire            n2685;
wire      [7:0] n2686;
wire            n2687;
wire      [7:0] n2688;
wire            n2689;
wire      [7:0] n269;
wire      [7:0] n2690;
wire            n2691;
wire      [7:0] n2692;
wire            n2693;
wire      [7:0] n2694;
wire            n2695;
wire      [7:0] n2696;
wire            n2697;
wire      [7:0] n2698;
wire            n2699;
wire      [7:0] n2700;
wire            n2701;
wire      [7:0] n2702;
wire            n2703;
wire      [7:0] n2704;
wire            n2705;
wire      [7:0] n2706;
wire            n2707;
wire      [7:0] n2708;
wire            n2709;
wire            n271;
wire      [7:0] n2710;
wire            n2711;
wire      [7:0] n2712;
wire            n2713;
wire      [7:0] n2714;
wire            n2715;
wire      [7:0] n2716;
wire            n2717;
wire      [7:0] n2718;
wire            n2719;
wire      [7:0] n2720;
wire            n2721;
wire      [7:0] n2722;
wire            n2723;
wire      [7:0] n2724;
wire            n2725;
wire      [7:0] n2726;
wire            n2727;
wire      [7:0] n2728;
wire            n2729;
wire      [7:0] n273;
wire      [7:0] n2730;
wire            n2731;
wire      [7:0] n2732;
wire            n2733;
wire      [7:0] n2734;
wire            n2735;
wire      [7:0] n2736;
wire            n2737;
wire      [7:0] n2738;
wire            n2739;
wire      [7:0] n2740;
wire            n2741;
wire      [7:0] n2742;
wire            n2743;
wire      [7:0] n2744;
wire            n2745;
wire      [7:0] n2746;
wire            n2747;
wire      [7:0] n2748;
wire            n2749;
wire            n275;
wire      [7:0] n2750;
wire            n2751;
wire      [7:0] n2752;
wire            n2753;
wire      [7:0] n2754;
wire            n2755;
wire      [7:0] n2756;
wire            n2757;
wire      [7:0] n2758;
wire            n2759;
wire      [7:0] n2760;
wire            n2761;
wire      [7:0] n2762;
wire            n2763;
wire      [7:0] n2764;
wire            n2765;
wire      [7:0] n2766;
wire            n2767;
wire      [7:0] n2768;
wire            n2769;
wire      [7:0] n277;
wire      [7:0] n2770;
wire            n2771;
wire      [7:0] n2772;
wire            n2773;
wire      [7:0] n2774;
wire            n2775;
wire      [7:0] n2776;
wire            n2777;
wire      [7:0] n2778;
wire            n2779;
wire      [7:0] n2780;
wire            n2781;
wire      [7:0] n2782;
wire            n2783;
wire      [7:0] n2784;
wire            n2785;
wire      [7:0] n2786;
wire            n2787;
wire      [7:0] n2788;
wire            n2789;
wire            n279;
wire      [7:0] n2790;
wire            n2791;
wire      [7:0] n2792;
wire            n2793;
wire      [7:0] n2794;
wire            n2795;
wire      [7:0] n2796;
wire            n2797;
wire      [7:0] n2798;
wire            n2799;
wire      [7:0] n28;
wire      [7:0] n2800;
wire            n2801;
wire      [7:0] n2802;
wire            n2803;
wire      [7:0] n2804;
wire            n2805;
wire      [7:0] n2806;
wire            n2807;
wire      [7:0] n2808;
wire            n2809;
wire      [7:0] n281;
wire      [7:0] n2810;
wire            n2811;
wire      [7:0] n2812;
wire            n2813;
wire      [7:0] n2814;
wire            n2815;
wire      [7:0] n2816;
wire            n2817;
wire      [7:0] n2818;
wire            n2819;
wire            n282;
wire      [7:0] n2820;
wire            n2821;
wire      [7:0] n2822;
wire            n2823;
wire      [7:0] n2824;
wire            n2825;
wire      [7:0] n2826;
wire            n2827;
wire      [7:0] n2828;
wire            n2829;
wire      [7:0] n283;
wire      [7:0] n2830;
wire            n2831;
wire      [7:0] n2832;
wire            n2833;
wire      [7:0] n2834;
wire            n2835;
wire      [7:0] n2836;
wire            n2837;
wire      [7:0] n2838;
wire            n2839;
wire            n284;
wire      [7:0] n2840;
wire            n2841;
wire      [7:0] n2842;
wire            n2843;
wire      [7:0] n2844;
wire            n2845;
wire      [7:0] n2846;
wire            n2847;
wire      [7:0] n2848;
wire            n2849;
wire      [7:0] n2850;
wire            n2851;
wire      [7:0] n2852;
wire            n2853;
wire      [7:0] n2854;
wire            n2855;
wire      [7:0] n2856;
wire            n2857;
wire      [7:0] n2858;
wire            n2859;
wire      [7:0] n286;
wire      [7:0] n2860;
wire            n2861;
wire      [7:0] n2862;
wire            n2863;
wire      [7:0] n2864;
wire            n2865;
wire      [7:0] n2866;
wire            n2867;
wire      [7:0] n2868;
wire            n2869;
wire      [7:0] n2870;
wire            n2871;
wire      [7:0] n2872;
wire            n2873;
wire      [7:0] n2874;
wire            n2875;
wire      [7:0] n2876;
wire            n2877;
wire      [7:0] n2878;
wire            n2879;
wire            n288;
wire      [7:0] n2880;
wire            n2881;
wire      [7:0] n2882;
wire            n2883;
wire      [7:0] n2884;
wire            n2885;
wire      [7:0] n2886;
wire            n2887;
wire      [7:0] n2888;
wire            n2889;
wire      [7:0] n2890;
wire            n2891;
wire      [7:0] n2892;
wire            n2893;
wire      [7:0] n2894;
wire            n2895;
wire      [7:0] n2896;
wire            n2897;
wire      [7:0] n2898;
wire            n2899;
wire      [7:0] n290;
wire      [7:0] n2900;
wire            n2901;
wire      [7:0] n2902;
wire            n2903;
wire      [7:0] n2904;
wire            n2905;
wire      [7:0] n2906;
wire            n2907;
wire      [7:0] n2908;
wire            n2909;
wire      [7:0] n2910;
wire            n2911;
wire      [7:0] n2912;
wire            n2913;
wire      [7:0] n2914;
wire            n2915;
wire      [7:0] n2916;
wire            n2917;
wire      [7:0] n2918;
wire            n2919;
wire            n292;
wire      [7:0] n2920;
wire            n2921;
wire      [7:0] n2922;
wire            n2923;
wire      [7:0] n2924;
wire            n2925;
wire      [7:0] n2926;
wire            n2927;
wire      [7:0] n2928;
wire            n2929;
wire      [7:0] n2930;
wire            n2931;
wire      [7:0] n2932;
wire            n2933;
wire      [7:0] n2934;
wire            n2935;
wire      [7:0] n2936;
wire            n2937;
wire      [7:0] n2938;
wire            n2939;
wire      [7:0] n294;
wire      [7:0] n2940;
wire            n2941;
wire      [7:0] n2942;
wire            n2943;
wire      [7:0] n2944;
wire            n2945;
wire      [7:0] n2946;
wire            n2947;
wire      [7:0] n2948;
wire            n2949;
wire      [7:0] n2950;
wire            n2951;
wire      [7:0] n2952;
wire            n2953;
wire      [7:0] n2954;
wire            n2955;
wire      [7:0] n2956;
wire            n2957;
wire      [7:0] n2958;
wire            n2959;
wire            n296;
wire      [7:0] n2960;
wire            n2961;
wire      [7:0] n2962;
wire            n2963;
wire      [7:0] n2964;
wire            n2965;
wire      [7:0] n2966;
wire            n2967;
wire      [7:0] n2968;
wire            n2969;
wire      [7:0] n297;
wire      [7:0] n2970;
wire            n2971;
wire      [7:0] n2972;
wire            n2973;
wire      [7:0] n2974;
wire            n2975;
wire      [7:0] n2976;
wire            n2977;
wire      [7:0] n2978;
wire            n2979;
wire            n298;
wire      [7:0] n2980;
wire            n2981;
wire      [7:0] n2982;
wire            n2983;
wire      [7:0] n2984;
wire            n2985;
wire      [7:0] n2986;
wire            n2987;
wire      [7:0] n2988;
wire            n2989;
wire      [7:0] n299;
wire      [7:0] n2990;
wire            n2991;
wire      [7:0] n2992;
wire            n2993;
wire      [7:0] n2994;
wire            n2995;
wire      [7:0] n2996;
wire            n2997;
wire      [7:0] n2998;
wire            n2999;
wire      [7:0] n3;
wire            n30;
wire      [7:0] n3000;
wire            n3001;
wire      [7:0] n3002;
wire            n3003;
wire      [7:0] n3004;
wire            n3005;
wire      [7:0] n3006;
wire            n3007;
wire      [7:0] n3008;
wire            n3009;
wire            n301;
wire      [7:0] n3010;
wire            n3011;
wire      [7:0] n3012;
wire            n3013;
wire      [7:0] n3014;
wire            n3015;
wire      [7:0] n3016;
wire            n3017;
wire      [7:0] n3018;
wire            n3019;
wire      [7:0] n3020;
wire            n3021;
wire      [7:0] n3022;
wire            n3023;
wire      [7:0] n3024;
wire            n3025;
wire      [7:0] n3026;
wire            n3027;
wire      [7:0] n3028;
wire            n3029;
wire      [7:0] n303;
wire      [7:0] n3030;
wire            n3031;
wire      [7:0] n3032;
wire            n3033;
wire      [7:0] n3034;
wire            n3035;
wire      [7:0] n3036;
wire            n3037;
wire      [7:0] n3038;
wire            n3039;
wire            n304;
wire      [7:0] n3040;
wire            n3041;
wire      [7:0] n3042;
wire            n3043;
wire      [7:0] n3044;
wire            n3045;
wire      [7:0] n3046;
wire            n3047;
wire      [7:0] n3048;
wire            n3049;
wire      [7:0] n305;
wire      [7:0] n3050;
wire            n3051;
wire      [7:0] n3052;
wire            n3053;
wire      [7:0] n3054;
wire            n3055;
wire      [7:0] n3056;
wire            n3057;
wire      [7:0] n3058;
wire            n3059;
wire      [7:0] n3060;
wire            n3061;
wire      [7:0] n3062;
wire            n3063;
wire      [7:0] n3064;
wire            n3065;
wire      [7:0] n3066;
wire            n3067;
wire      [7:0] n3068;
wire            n3069;
wire            n307;
wire      [7:0] n3070;
wire            n3071;
wire      [7:0] n3072;
wire            n3073;
wire      [7:0] n3074;
wire            n3075;
wire      [7:0] n3076;
wire            n3077;
wire      [7:0] n3078;
wire            n3079;
wire      [7:0] n3080;
wire            n3081;
wire      [7:0] n3082;
wire            n3083;
wire      [7:0] n3084;
wire      [7:0] n3085;
wire      [7:0] n3086;
wire      [7:0] n3087;
wire      [7:0] n3088;
wire      [7:0] n3089;
wire      [7:0] n309;
wire      [7:0] n3090;
wire      [7:0] n3091;
wire      [7:0] n3092;
wire      [7:0] n3093;
wire      [7:0] n3094;
wire      [7:0] n3095;
wire      [7:0] n3096;
wire      [7:0] n3097;
wire      [7:0] n3098;
wire      [7:0] n3099;
wire      [7:0] n3100;
wire      [7:0] n3101;
wire      [7:0] n3102;
wire      [7:0] n3103;
wire      [7:0] n3104;
wire      [7:0] n3105;
wire      [7:0] n3106;
wire      [7:0] n3107;
wire      [7:0] n3108;
wire      [7:0] n3109;
wire            n311;
wire      [7:0] n3110;
wire      [7:0] n3111;
wire      [7:0] n3112;
wire      [7:0] n3113;
wire      [7:0] n3114;
wire      [7:0] n3115;
wire      [7:0] n3116;
wire      [7:0] n3117;
wire      [7:0] n3118;
wire      [7:0] n3119;
wire      [7:0] n3120;
wire      [7:0] n3121;
wire      [7:0] n3122;
wire      [7:0] n3123;
wire      [7:0] n3124;
wire      [7:0] n3125;
wire      [7:0] n3126;
wire      [7:0] n3127;
wire      [7:0] n3128;
wire      [7:0] n3129;
wire      [7:0] n313;
wire      [7:0] n3130;
wire      [7:0] n3131;
wire      [7:0] n3132;
wire      [7:0] n3133;
wire      [7:0] n3134;
wire      [7:0] n3135;
wire      [7:0] n3136;
wire      [7:0] n3137;
wire      [7:0] n3138;
wire      [7:0] n3139;
wire      [7:0] n3140;
wire      [7:0] n3141;
wire      [7:0] n3142;
wire      [7:0] n3143;
wire      [7:0] n3144;
wire      [7:0] n3145;
wire      [7:0] n3146;
wire      [7:0] n3147;
wire      [7:0] n3148;
wire      [7:0] n3149;
wire            n315;
wire      [7:0] n3150;
wire      [7:0] n3151;
wire      [7:0] n3152;
wire      [7:0] n3153;
wire      [7:0] n3154;
wire      [7:0] n3155;
wire      [7:0] n3156;
wire      [7:0] n3157;
wire      [7:0] n3158;
wire      [7:0] n3159;
wire      [7:0] n3160;
wire      [7:0] n3161;
wire      [7:0] n3162;
wire      [7:0] n3163;
wire      [7:0] n3164;
wire      [7:0] n3165;
wire      [7:0] n3166;
wire      [7:0] n3167;
wire      [7:0] n3168;
wire      [7:0] n3169;
wire      [7:0] n317;
wire      [7:0] n3170;
wire      [7:0] n3171;
wire      [7:0] n3172;
wire      [7:0] n3173;
wire      [7:0] n3174;
wire      [7:0] n3175;
wire      [7:0] n3176;
wire      [7:0] n3177;
wire      [7:0] n3178;
wire      [7:0] n3179;
wire      [7:0] n3180;
wire      [7:0] n3181;
wire      [7:0] n3182;
wire      [7:0] n3183;
wire      [7:0] n3184;
wire      [7:0] n3185;
wire      [7:0] n3186;
wire      [7:0] n3187;
wire      [7:0] n3188;
wire      [7:0] n3189;
wire            n319;
wire      [7:0] n3190;
wire      [7:0] n3191;
wire      [7:0] n3192;
wire      [7:0] n3193;
wire      [7:0] n3194;
wire      [7:0] n3195;
wire      [7:0] n3196;
wire      [7:0] n3197;
wire      [7:0] n3198;
wire      [7:0] n3199;
wire      [7:0] n32;
wire      [7:0] n320;
wire      [7:0] n3200;
wire      [7:0] n3201;
wire      [7:0] n3202;
wire      [7:0] n3203;
wire      [7:0] n3204;
wire      [7:0] n3205;
wire      [7:0] n3206;
wire      [7:0] n3207;
wire      [7:0] n3208;
wire      [7:0] n3209;
wire            n321;
wire      [7:0] n3210;
wire      [7:0] n3211;
wire      [7:0] n3212;
wire      [7:0] n3213;
wire      [7:0] n3214;
wire      [7:0] n3215;
wire      [7:0] n3216;
wire      [7:0] n3217;
wire      [7:0] n3218;
wire      [7:0] n3219;
wire      [7:0] n322;
wire      [7:0] n3220;
wire      [7:0] n3221;
wire      [7:0] n3222;
wire      [7:0] n3223;
wire      [7:0] n3224;
wire      [7:0] n3225;
wire      [7:0] n3226;
wire      [7:0] n3227;
wire      [7:0] n3228;
wire      [7:0] n3229;
wire      [7:0] n3230;
wire      [7:0] n3231;
wire      [7:0] n3232;
wire      [7:0] n3233;
wire      [7:0] n3234;
wire      [7:0] n3235;
wire      [7:0] n3236;
wire      [7:0] n3237;
wire      [7:0] n3238;
wire      [7:0] n3239;
wire            n324;
wire      [7:0] n3240;
wire      [7:0] n3241;
wire      [7:0] n3242;
wire      [7:0] n3243;
wire      [7:0] n3244;
wire      [7:0] n3245;
wire      [7:0] n3246;
wire      [7:0] n3247;
wire      [7:0] n3248;
wire      [7:0] n3249;
wire      [7:0] n325;
wire      [7:0] n3250;
wire      [7:0] n3251;
wire      [7:0] n3252;
wire      [7:0] n3253;
wire      [7:0] n3254;
wire      [7:0] n3255;
wire      [7:0] n3256;
wire      [7:0] n3257;
wire      [7:0] n3258;
wire      [7:0] n3259;
wire      [7:0] n3260;
wire      [7:0] n3261;
wire      [7:0] n3262;
wire      [7:0] n3263;
wire      [7:0] n3264;
wire      [7:0] n3265;
wire      [7:0] n3266;
wire      [7:0] n3267;
wire      [7:0] n3268;
wire      [7:0] n3269;
wire            n327;
wire      [7:0] n3270;
wire      [7:0] n3271;
wire      [7:0] n3272;
wire      [7:0] n3273;
wire      [7:0] n3274;
wire      [7:0] n3275;
wire      [7:0] n3276;
wire      [7:0] n3277;
wire      [7:0] n3278;
wire      [7:0] n3279;
wire      [7:0] n3280;
wire      [7:0] n3281;
wire      [7:0] n3282;
wire      [7:0] n3283;
wire      [7:0] n3284;
wire      [7:0] n3285;
wire      [7:0] n3286;
wire      [7:0] n3287;
wire      [7:0] n3288;
wire      [7:0] n3289;
wire      [7:0] n329;
wire      [7:0] n3290;
wire      [7:0] n3291;
wire      [7:0] n3292;
wire      [7:0] n3293;
wire      [7:0] n3294;
wire      [7:0] n3295;
wire      [7:0] n3296;
wire      [7:0] n3297;
wire      [7:0] n3298;
wire      [7:0] n3299;
wire            n330;
wire      [7:0] n3300;
wire      [7:0] n3301;
wire      [7:0] n3302;
wire      [7:0] n3303;
wire      [7:0] n3304;
wire      [7:0] n3305;
wire      [7:0] n3306;
wire      [7:0] n3307;
wire      [7:0] n3308;
wire      [7:0] n3309;
wire      [7:0] n3310;
wire      [7:0] n3311;
wire      [7:0] n3312;
wire      [7:0] n3313;
wire      [7:0] n3314;
wire      [7:0] n3315;
wire      [7:0] n3316;
wire      [7:0] n3317;
wire      [7:0] n3318;
wire      [7:0] n3319;
wire      [7:0] n332;
wire      [7:0] n3320;
wire      [7:0] n3321;
wire      [7:0] n3322;
wire      [7:0] n3323;
wire      [7:0] n3324;
wire      [7:0] n3325;
wire      [7:0] n3326;
wire      [7:0] n3327;
wire      [7:0] n3328;
wire      [7:0] n3329;
wire      [7:0] n3330;
wire      [7:0] n3331;
wire      [7:0] n3332;
wire      [7:0] n3333;
wire      [7:0] n3334;
wire      [7:0] n3335;
wire      [7:0] n3336;
wire      [7:0] n3337;
wire      [7:0] n3338;
wire      [7:0] n3339;
wire            n334;
wire      [7:0] n3340;
wire     [31:0] n3341;
wire      [7:0] n3342;
wire      [7:0] n3343;
wire      [7:0] n3344;
wire      [7:0] n3345;
wire      [7:0] n3346;
wire     [39:0] n3347;
wire      [7:0] n3348;
wire      [7:0] n3349;
wire      [7:0] n3350;
wire      [7:0] n3351;
wire     [47:0] n3352;
wire      [7:0] n3353;
wire      [7:0] n3354;
wire      [7:0] n3355;
wire      [7:0] n3356;
wire     [55:0] n3357;
wire      [7:0] n3358;
wire      [7:0] n3359;
wire      [7:0] n336;
wire      [7:0] n3360;
wire      [7:0] n3361;
wire     [63:0] n3362;
wire      [7:0] n3363;
wire      [7:0] n3364;
wire      [7:0] n3365;
wire      [7:0] n3366;
wire      [7:0] n3367;
wire      [7:0] n3368;
wire      [7:0] n3369;
wire     [71:0] n3370;
wire      [7:0] n3371;
wire      [7:0] n3372;
wire      [7:0] n3373;
wire      [7:0] n3374;
wire      [7:0] n3375;
wire      [7:0] n3376;
wire     [79:0] n3377;
wire      [7:0] n3378;
wire      [7:0] n3379;
wire            n338;
wire      [7:0] n3380;
wire      [7:0] n3381;
wire      [7:0] n3382;
wire      [7:0] n3383;
wire     [87:0] n3384;
wire      [7:0] n3385;
wire      [7:0] n3386;
wire      [7:0] n3387;
wire      [7:0] n3388;
wire      [7:0] n3389;
wire      [7:0] n3390;
wire     [95:0] n3391;
wire      [7:0] n3392;
wire      [7:0] n3393;
wire      [7:0] n3394;
wire      [7:0] n3395;
wire      [7:0] n3396;
wire      [7:0] n3397;
wire      [7:0] n3398;
wire      [7:0] n3399;
wire            n34;
wire      [7:0] n340;
wire      [7:0] n3400;
wire    [103:0] n3401;
wire      [7:0] n3402;
wire      [7:0] n3403;
wire      [7:0] n3404;
wire      [7:0] n3405;
wire      [7:0] n3406;
wire      [7:0] n3407;
wire      [7:0] n3408;
wire      [7:0] n3409;
wire    [111:0] n3410;
wire      [7:0] n3411;
wire      [7:0] n3412;
wire      [7:0] n3413;
wire      [7:0] n3414;
wire      [7:0] n3415;
wire      [7:0] n3416;
wire      [7:0] n3417;
wire      [7:0] n3418;
wire    [119:0] n3419;
wire            n342;
wire      [7:0] n3420;
wire      [7:0] n3421;
wire      [7:0] n3422;
wire      [7:0] n3423;
wire      [7:0] n3424;
wire      [7:0] n3425;
wire      [7:0] n3426;
wire      [7:0] n3427;
wire    [127:0] n3428;
wire    [127:0] n3429;
wire      [7:0] n344;
wire            n346;
wire      [7:0] n348;
wire            n349;
wire      [7:0] n351;
wire            n353;
wire      [7:0] n354;
wire            n356;
wire      [7:0] n357;
wire            n358;
wire      [7:0] n36;
wire      [7:0] n360;
wire            n362;
wire      [7:0] n364;
wire            n366;
wire      [7:0] n367;
wire            n368;
wire      [7:0] n370;
wire            n372;
wire      [7:0] n373;
wire            n374;
wire      [7:0] n375;
wire            n376;
wire      [7:0] n378;
wire            n38;
wire            n380;
wire      [7:0] n382;
wire            n384;
wire      [7:0] n386;
wire            n387;
wire      [7:0] n389;
wire            n390;
wire      [7:0] n392;
wire            n394;
wire      [7:0] n395;
wire            n397;
wire      [7:0] n399;
wire      [7:0] n4;
wire      [7:0] n40;
wire            n400;
wire      [7:0] n402;
wire            n403;
wire      [7:0] n405;
wire            n407;
wire      [7:0] n409;
wire            n410;
wire      [7:0] n412;
wire            n413;
wire      [7:0] n415;
wire            n416;
wire      [7:0] n418;
wire            n419;
wire            n42;
wire      [7:0] n421;
wire            n422;
wire      [7:0] n424;
wire            n425;
wire      [7:0] n426;
wire            n427;
wire      [7:0] n428;
wire            n429;
wire      [7:0] n431;
wire            n432;
wire      [7:0] n434;
wire            n436;
wire      [7:0] n437;
wire            n439;
wire      [7:0] n44;
wire      [7:0] n441;
wire            n443;
wire      [7:0] n444;
wire            n446;
wire      [7:0] n448;
wire            n449;
wire      [7:0] n451;
wire            n453;
wire      [7:0] n454;
wire            n456;
wire      [7:0] n457;
wire            n458;
wire      [7:0] n459;
wire            n46;
wire            n461;
wire      [7:0] n462;
wire            n464;
wire      [7:0] n466;
wire            n468;
wire      [7:0] n470;
wire            n471;
wire      [7:0] n472;
wire            n473;
wire      [7:0] n474;
wire            n475;
wire      [7:0] n476;
wire            n478;
wire      [7:0] n479;
wire      [7:0] n48;
wire            n481;
wire      [7:0] n483;
wire            n485;
wire      [7:0] n486;
wire            n487;
wire      [7:0] n488;
wire            n489;
wire      [7:0] n490;
wire            n492;
wire      [7:0] n494;
wire            n496;
wire      [7:0] n497;
wire            n498;
wire            n50;
wire      [7:0] n500;
wire            n502;
wire      [7:0] n503;
wire            n505;
wire      [7:0] n506;
wire            n507;
wire      [7:0] n509;
wire            n510;
wire      [7:0] n512;
wire            n514;
wire      [7:0] n515;
wire            n517;
wire      [7:0] n519;
wire      [7:0] n52;
wire            n520;
wire      [7:0] n521;
wire            n522;
wire      [7:0] n524;
wire            n526;
wire      [7:0] n527;
wire            n528;
wire      [7:0] n530;
wire            n531;
wire      [7:0] n533;
wire            n534;
wire      [7:0] n536;
wire            n538;
wire      [7:0] n539;
wire            n54;
wire            n540;
wire      [7:0] n541;
wire            n542;
wire      [7:0] n543;
wire            n544;
wire      [7:0] n545;
wire            n546;
wire      [7:0] n547;
wire            n548;
wire      [7:0] n550;
wire            n551;
wire      [7:0] n553;
wire            n554;
wire      [7:0] n556;
wire            n558;
wire      [7:0] n56;
wire      [7:0] n560;
wire            n562;
wire      [7:0] n563;
wire            n565;
wire      [7:0] n566;
wire            n567;
wire      [7:0] n568;
wire            n569;
wire      [7:0] n570;
wire            n571;
wire      [7:0] n572;
wire            n573;
wire      [7:0] n574;
wire            n575;
wire      [7:0] n577;
wire            n579;
wire            n58;
wire      [7:0] n580;
wire            n582;
wire      [7:0] n584;
wire            n585;
wire      [7:0] n586;
wire            n587;
wire      [7:0] n588;
wire            n589;
wire      [7:0] n590;
wire            n591;
wire      [7:0] n593;
wire            n594;
wire      [7:0] n595;
wire            n596;
wire      [7:0] n598;
wire            n599;
wire            n6;
wire      [7:0] n60;
wire      [7:0] n600;
wire            n601;
wire      [7:0] n602;
wire            n603;
wire      [7:0] n605;
wire            n606;
wire      [7:0] n607;
wire            n609;
wire      [7:0] n610;
wire            n611;
wire      [7:0] n612;
wire            n613;
wire      [7:0] n614;
wire            n615;
wire      [7:0] n617;
wire            n618;
wire            n62;
wire      [7:0] n620;
wire            n621;
wire      [7:0] n623;
wire            n624;
wire      [7:0] n625;
wire            n626;
wire      [7:0] n628;
wire            n630;
wire      [7:0] n631;
wire            n632;
wire      [7:0] n633;
wire            n634;
wire      [7:0] n636;
wire            n637;
wire      [7:0] n638;
wire            n639;
wire      [7:0] n64;
wire      [7:0] n640;
wire            n641;
wire      [7:0] n642;
wire            n643;
wire      [7:0] n645;
wire            n646;
wire      [7:0] n648;
wire            n649;
wire      [7:0] n650;
wire            n652;
wire      [7:0] n654;
wire            n655;
wire      [7:0] n656;
wire            n658;
wire            n66;
wire      [7:0] n660;
wire            n661;
wire      [7:0] n662;
wire            n663;
wire      [7:0] n665;
wire            n667;
wire      [7:0] n668;
wire            n670;
wire      [7:0] n672;
wire            n673;
wire      [7:0] n675;
wire            n676;
wire      [7:0] n677;
wire            n678;
wire      [7:0] n679;
wire      [7:0] n68;
wire            n680;
wire      [7:0] n681;
wire            n683;
wire      [7:0] n684;
wire            n685;
wire      [7:0] n686;
wire            n687;
wire      [7:0] n688;
wire            n689;
wire      [7:0] n690;
wire            n691;
wire      [7:0] n692;
wire            n694;
wire      [7:0] n695;
wire            n696;
wire      [7:0] n697;
wire            n698;
wire      [7:0] n699;
wire            n70;
wire            n700;
wire      [7:0] n701;
wire            n702;
wire      [7:0] n703;
wire            n704;
wire      [7:0] n705;
wire            n706;
wire      [7:0] n707;
wire            n708;
wire      [7:0] n709;
wire            n710;
wire      [7:0] n711;
wire            n712;
wire      [7:0] n713;
wire            n714;
wire      [7:0] n715;
wire            n716;
wire      [7:0] n717;
wire            n718;
wire      [7:0] n719;
wire      [7:0] n72;
wire            n720;
wire      [7:0] n721;
wire            n722;
wire      [7:0] n723;
wire            n724;
wire      [7:0] n725;
wire            n726;
wire      [7:0] n727;
wire            n728;
wire      [7:0] n729;
wire            n730;
wire      [7:0] n731;
wire            n732;
wire      [7:0] n733;
wire            n734;
wire      [7:0] n735;
wire            n736;
wire      [7:0] n737;
wire            n738;
wire      [7:0] n739;
wire            n74;
wire            n740;
wire      [7:0] n741;
wire            n742;
wire      [7:0] n743;
wire            n744;
wire      [7:0] n745;
wire            n746;
wire      [7:0] n747;
wire            n748;
wire      [7:0] n749;
wire            n750;
wire      [7:0] n751;
wire            n752;
wire      [7:0] n754;
wire            n755;
wire      [7:0] n756;
wire            n757;
wire      [7:0] n758;
wire            n759;
wire      [7:0] n76;
wire      [7:0] n760;
wire            n761;
wire      [7:0] n762;
wire            n763;
wire      [7:0] n764;
wire            n765;
wire      [7:0] n766;
wire            n767;
wire      [7:0] n768;
wire            n769;
wire      [7:0] n770;
wire            n771;
wire      [7:0] n772;
wire      [7:0] n773;
wire      [7:0] n774;
wire      [7:0] n775;
wire      [7:0] n776;
wire      [7:0] n777;
wire      [7:0] n778;
wire      [7:0] n779;
wire            n78;
wire      [7:0] n780;
wire      [7:0] n781;
wire      [7:0] n782;
wire      [7:0] n783;
wire      [7:0] n784;
wire      [7:0] n785;
wire      [7:0] n786;
wire      [7:0] n787;
wire      [7:0] n788;
wire      [7:0] n789;
wire      [7:0] n790;
wire      [7:0] n791;
wire      [7:0] n792;
wire      [7:0] n793;
wire      [7:0] n794;
wire      [7:0] n795;
wire      [7:0] n796;
wire      [7:0] n797;
wire      [7:0] n798;
wire      [7:0] n799;
wire      [7:0] n8;
wire      [7:0] n80;
wire      [7:0] n800;
wire      [7:0] n801;
wire      [7:0] n802;
wire      [7:0] n803;
wire      [7:0] n804;
wire      [7:0] n805;
wire      [7:0] n806;
wire      [7:0] n807;
wire      [7:0] n808;
wire      [7:0] n809;
wire      [7:0] n810;
wire      [7:0] n811;
wire      [7:0] n812;
wire      [7:0] n813;
wire      [7:0] n814;
wire      [7:0] n815;
wire      [7:0] n816;
wire      [7:0] n817;
wire      [7:0] n818;
wire      [7:0] n819;
wire            n82;
wire      [7:0] n820;
wire      [7:0] n821;
wire      [7:0] n822;
wire      [7:0] n823;
wire      [7:0] n824;
wire      [7:0] n825;
wire      [7:0] n826;
wire      [7:0] n827;
wire      [7:0] n828;
wire      [7:0] n829;
wire      [7:0] n830;
wire      [7:0] n831;
wire      [7:0] n832;
wire      [7:0] n833;
wire      [7:0] n834;
wire      [7:0] n835;
wire      [7:0] n836;
wire      [7:0] n837;
wire      [7:0] n838;
wire      [7:0] n839;
wire      [7:0] n84;
wire      [7:0] n840;
wire      [7:0] n841;
wire      [7:0] n842;
wire      [7:0] n843;
wire      [7:0] n844;
wire      [7:0] n845;
wire      [7:0] n846;
wire      [7:0] n847;
wire      [7:0] n848;
wire      [7:0] n849;
wire      [7:0] n850;
wire      [7:0] n851;
wire      [7:0] n852;
wire      [7:0] n853;
wire      [7:0] n854;
wire      [7:0] n855;
wire      [7:0] n856;
wire      [7:0] n857;
wire      [7:0] n858;
wire      [7:0] n859;
wire            n86;
wire      [7:0] n860;
wire      [7:0] n861;
wire      [7:0] n862;
wire      [7:0] n863;
wire      [7:0] n864;
wire      [7:0] n865;
wire      [7:0] n866;
wire      [7:0] n867;
wire      [7:0] n868;
wire      [7:0] n869;
wire      [7:0] n870;
wire      [7:0] n871;
wire      [7:0] n872;
wire      [7:0] n873;
wire      [7:0] n874;
wire      [7:0] n875;
wire      [7:0] n876;
wire      [7:0] n877;
wire      [7:0] n878;
wire      [7:0] n879;
wire      [7:0] n88;
wire      [7:0] n880;
wire      [7:0] n881;
wire      [7:0] n882;
wire      [7:0] n883;
wire      [7:0] n884;
wire      [7:0] n885;
wire      [7:0] n886;
wire      [7:0] n887;
wire      [7:0] n888;
wire      [7:0] n889;
wire      [7:0] n890;
wire      [7:0] n891;
wire      [7:0] n892;
wire      [7:0] n893;
wire      [7:0] n894;
wire      [7:0] n895;
wire      [7:0] n896;
wire      [7:0] n897;
wire      [7:0] n898;
wire      [7:0] n899;
wire            n90;
wire      [7:0] n900;
wire      [7:0] n901;
wire      [7:0] n902;
wire      [7:0] n903;
wire      [7:0] n904;
wire      [7:0] n905;
wire      [7:0] n906;
wire      [7:0] n907;
wire      [7:0] n908;
wire      [7:0] n909;
wire      [7:0] n910;
wire      [7:0] n911;
wire      [7:0] n912;
wire      [7:0] n913;
wire      [7:0] n914;
wire      [7:0] n915;
wire      [7:0] n916;
wire      [7:0] n917;
wire      [7:0] n918;
wire      [7:0] n919;
wire      [7:0] n92;
wire      [7:0] n920;
wire      [7:0] n921;
wire      [7:0] n922;
wire      [7:0] n923;
wire      [7:0] n924;
wire      [7:0] n925;
wire      [7:0] n926;
wire      [7:0] n927;
wire      [7:0] n928;
wire      [7:0] n929;
wire            n93;
wire      [7:0] n930;
wire      [7:0] n931;
wire      [7:0] n932;
wire      [7:0] n933;
wire      [7:0] n934;
wire      [7:0] n935;
wire      [7:0] n936;
wire      [7:0] n937;
wire      [7:0] n938;
wire      [7:0] n939;
wire      [7:0] n940;
wire      [7:0] n941;
wire      [7:0] n942;
wire      [7:0] n943;
wire      [7:0] n944;
wire      [7:0] n945;
wire      [7:0] n946;
wire      [7:0] n947;
wire      [7:0] n948;
wire      [7:0] n949;
wire      [7:0] n95;
wire      [7:0] n950;
wire      [7:0] n951;
wire      [7:0] n952;
wire      [7:0] n953;
wire      [7:0] n954;
wire      [7:0] n955;
wire      [7:0] n956;
wire      [7:0] n957;
wire      [7:0] n958;
wire      [7:0] n959;
wire      [7:0] n960;
wire      [7:0] n961;
wire      [7:0] n962;
wire      [7:0] n963;
wire      [7:0] n964;
wire      [7:0] n965;
wire      [7:0] n966;
wire      [7:0] n967;
wire      [7:0] n968;
wire      [7:0] n969;
wire            n97;
wire      [7:0] n970;
wire      [7:0] n971;
wire      [7:0] n972;
wire      [7:0] n973;
wire      [7:0] n974;
wire      [7:0] n975;
wire      [7:0] n976;
wire      [7:0] n977;
wire      [7:0] n978;
wire      [7:0] n979;
wire      [7:0] n980;
wire      [7:0] n981;
wire      [7:0] n982;
wire      [7:0] n983;
wire      [7:0] n984;
wire      [7:0] n985;
wire      [7:0] n986;
wire      [7:0] n987;
wire      [7:0] n988;
wire      [7:0] n989;
wire      [7:0] n99;
wire      [7:0] n990;
wire      [7:0] n991;
wire      [7:0] n992;
wire      [7:0] n993;
wire      [7:0] n994;
wire      [7:0] n995;
wire      [7:0] n996;
wire      [7:0] n997;
wire      [7:0] n998;
wire      [7:0] n999;
wire            rst;
assign __ILA_bar_valid__ = 1'b1 ;
assign __ILA_bar_decode_of_i1__ = 1'b1 ;
assign bv_128_0_n1 = 128'h0 ;
assign n2 = in[127:120] ;
assign n3 =  ( n2 ) ^ ( rcon )  ;
assign n4 = in[23:16] ;
assign bv_8_255_n5 = 8'hff ;
assign n6 =  ( n4 ) == ( bv_8_255_n5 )  ;
assign bv_8_22_n7 = 8'h16 ;
assign n8 = in[23:16] ;
assign bv_8_254_n9 = 8'hfe ;
assign n10 =  ( n8 ) == ( bv_8_254_n9 )  ;
assign bv_8_187_n11 = 8'hbb ;
assign n12 = in[23:16] ;
assign bv_8_253_n13 = 8'hfd ;
assign n14 =  ( n12 ) == ( bv_8_253_n13 )  ;
assign bv_8_84_n15 = 8'h54 ;
assign n16 = in[23:16] ;
assign bv_8_252_n17 = 8'hfc ;
assign n18 =  ( n16 ) == ( bv_8_252_n17 )  ;
assign bv_8_176_n19 = 8'hb0 ;
assign n20 = in[23:16] ;
assign bv_8_251_n21 = 8'hfb ;
assign n22 =  ( n20 ) == ( bv_8_251_n21 )  ;
assign bv_8_15_n23 = 8'hf ;
assign n24 = in[23:16] ;
assign bv_8_250_n25 = 8'hfa ;
assign n26 =  ( n24 ) == ( bv_8_250_n25 )  ;
assign bv_8_45_n27 = 8'h2d ;
assign n28 = in[23:16] ;
assign bv_8_249_n29 = 8'hf9 ;
assign n30 =  ( n28 ) == ( bv_8_249_n29 )  ;
assign bv_8_153_n31 = 8'h99 ;
assign n32 = in[23:16] ;
assign bv_8_248_n33 = 8'hf8 ;
assign n34 =  ( n32 ) == ( bv_8_248_n33 )  ;
assign bv_8_65_n35 = 8'h41 ;
assign n36 = in[23:16] ;
assign bv_8_247_n37 = 8'hf7 ;
assign n38 =  ( n36 ) == ( bv_8_247_n37 )  ;
assign bv_8_104_n39 = 8'h68 ;
assign n40 = in[23:16] ;
assign bv_8_246_n41 = 8'hf6 ;
assign n42 =  ( n40 ) == ( bv_8_246_n41 )  ;
assign bv_8_66_n43 = 8'h42 ;
assign n44 = in[23:16] ;
assign bv_8_245_n45 = 8'hf5 ;
assign n46 =  ( n44 ) == ( bv_8_245_n45 )  ;
assign bv_8_230_n47 = 8'he6 ;
assign n48 = in[23:16] ;
assign bv_8_244_n49 = 8'hf4 ;
assign n50 =  ( n48 ) == ( bv_8_244_n49 )  ;
assign bv_8_191_n51 = 8'hbf ;
assign n52 = in[23:16] ;
assign bv_8_243_n53 = 8'hf3 ;
assign n54 =  ( n52 ) == ( bv_8_243_n53 )  ;
assign bv_8_13_n55 = 8'hd ;
assign n56 = in[23:16] ;
assign bv_8_242_n57 = 8'hf2 ;
assign n58 =  ( n56 ) == ( bv_8_242_n57 )  ;
assign bv_8_137_n59 = 8'h89 ;
assign n60 = in[23:16] ;
assign bv_8_241_n61 = 8'hf1 ;
assign n62 =  ( n60 ) == ( bv_8_241_n61 )  ;
assign bv_8_161_n63 = 8'ha1 ;
assign n64 = in[23:16] ;
assign bv_8_240_n65 = 8'hf0 ;
assign n66 =  ( n64 ) == ( bv_8_240_n65 )  ;
assign bv_8_140_n67 = 8'h8c ;
assign n68 = in[23:16] ;
assign bv_8_239_n69 = 8'hef ;
assign n70 =  ( n68 ) == ( bv_8_239_n69 )  ;
assign bv_8_223_n71 = 8'hdf ;
assign n72 = in[23:16] ;
assign bv_8_238_n73 = 8'hee ;
assign n74 =  ( n72 ) == ( bv_8_238_n73 )  ;
assign bv_8_40_n75 = 8'h28 ;
assign n76 = in[23:16] ;
assign bv_8_237_n77 = 8'hed ;
assign n78 =  ( n76 ) == ( bv_8_237_n77 )  ;
assign bv_8_85_n79 = 8'h55 ;
assign n80 = in[23:16] ;
assign bv_8_236_n81 = 8'hec ;
assign n82 =  ( n80 ) == ( bv_8_236_n81 )  ;
assign bv_8_206_n83 = 8'hce ;
assign n84 = in[23:16] ;
assign bv_8_235_n85 = 8'heb ;
assign n86 =  ( n84 ) == ( bv_8_235_n85 )  ;
assign bv_8_233_n87 = 8'he9 ;
assign n88 = in[23:16] ;
assign bv_8_234_n89 = 8'hea ;
assign n90 =  ( n88 ) == ( bv_8_234_n89 )  ;
assign bv_8_135_n91 = 8'h87 ;
assign n92 = in[23:16] ;
assign n93 =  ( n92 ) == ( bv_8_233_n87 )  ;
assign bv_8_30_n94 = 8'h1e ;
assign n95 = in[23:16] ;
assign bv_8_232_n96 = 8'he8 ;
assign n97 =  ( n95 ) == ( bv_8_232_n96 )  ;
assign bv_8_155_n98 = 8'h9b ;
assign n99 = in[23:16] ;
assign bv_8_231_n100 = 8'he7 ;
assign n101 =  ( n99 ) == ( bv_8_231_n100 )  ;
assign bv_8_148_n102 = 8'h94 ;
assign n103 = in[23:16] ;
assign n104 =  ( n103 ) == ( bv_8_230_n47 )  ;
assign bv_8_142_n105 = 8'h8e ;
assign n106 = in[23:16] ;
assign bv_8_229_n107 = 8'he5 ;
assign n108 =  ( n106 ) == ( bv_8_229_n107 )  ;
assign bv_8_217_n109 = 8'hd9 ;
assign n110 = in[23:16] ;
assign bv_8_228_n111 = 8'he4 ;
assign n112 =  ( n110 ) == ( bv_8_228_n111 )  ;
assign bv_8_105_n113 = 8'h69 ;
assign n114 = in[23:16] ;
assign bv_8_227_n115 = 8'he3 ;
assign n116 =  ( n114 ) == ( bv_8_227_n115 )  ;
assign bv_8_17_n117 = 8'h11 ;
assign n118 = in[23:16] ;
assign bv_8_226_n119 = 8'he2 ;
assign n120 =  ( n118 ) == ( bv_8_226_n119 )  ;
assign bv_8_152_n121 = 8'h98 ;
assign n122 = in[23:16] ;
assign bv_8_225_n123 = 8'he1 ;
assign n124 =  ( n122 ) == ( bv_8_225_n123 )  ;
assign n125 = in[23:16] ;
assign bv_8_224_n126 = 8'he0 ;
assign n127 =  ( n125 ) == ( bv_8_224_n126 )  ;
assign n128 = in[23:16] ;
assign n129 =  ( n128 ) == ( bv_8_223_n71 )  ;
assign bv_8_158_n130 = 8'h9e ;
assign n131 = in[23:16] ;
assign bv_8_222_n132 = 8'hde ;
assign n133 =  ( n131 ) == ( bv_8_222_n132 )  ;
assign bv_8_29_n134 = 8'h1d ;
assign n135 = in[23:16] ;
assign bv_8_221_n136 = 8'hdd ;
assign n137 =  ( n135 ) == ( bv_8_221_n136 )  ;
assign bv_8_193_n138 = 8'hc1 ;
assign n139 = in[23:16] ;
assign bv_8_220_n140 = 8'hdc ;
assign n141 =  ( n139 ) == ( bv_8_220_n140 )  ;
assign bv_8_134_n142 = 8'h86 ;
assign n143 = in[23:16] ;
assign bv_8_219_n144 = 8'hdb ;
assign n145 =  ( n143 ) == ( bv_8_219_n144 )  ;
assign bv_8_185_n146 = 8'hb9 ;
assign n147 = in[23:16] ;
assign bv_8_218_n148 = 8'hda ;
assign n149 =  ( n147 ) == ( bv_8_218_n148 )  ;
assign bv_8_87_n150 = 8'h57 ;
assign n151 = in[23:16] ;
assign n152 =  ( n151 ) == ( bv_8_217_n109 )  ;
assign bv_8_53_n153 = 8'h35 ;
assign n154 = in[23:16] ;
assign bv_8_216_n155 = 8'hd8 ;
assign n156 =  ( n154 ) == ( bv_8_216_n155 )  ;
assign bv_8_97_n157 = 8'h61 ;
assign n158 = in[23:16] ;
assign bv_8_215_n159 = 8'hd7 ;
assign n160 =  ( n158 ) == ( bv_8_215_n159 )  ;
assign bv_8_14_n161 = 8'he ;
assign n162 = in[23:16] ;
assign bv_8_214_n163 = 8'hd6 ;
assign n164 =  ( n162 ) == ( bv_8_214_n163 )  ;
assign n165 = in[23:16] ;
assign bv_8_213_n166 = 8'hd5 ;
assign n167 =  ( n165 ) == ( bv_8_213_n166 )  ;
assign bv_8_3_n168 = 8'h3 ;
assign n169 = in[23:16] ;
assign bv_8_212_n170 = 8'hd4 ;
assign n171 =  ( n169 ) == ( bv_8_212_n170 )  ;
assign bv_8_72_n172 = 8'h48 ;
assign n173 = in[23:16] ;
assign bv_8_211_n174 = 8'hd3 ;
assign n175 =  ( n173 ) == ( bv_8_211_n174 )  ;
assign bv_8_102_n176 = 8'h66 ;
assign n177 = in[23:16] ;
assign bv_8_210_n178 = 8'hd2 ;
assign n179 =  ( n177 ) == ( bv_8_210_n178 )  ;
assign bv_8_181_n180 = 8'hb5 ;
assign n181 = in[23:16] ;
assign bv_8_209_n182 = 8'hd1 ;
assign n183 =  ( n181 ) == ( bv_8_209_n182 )  ;
assign bv_8_62_n184 = 8'h3e ;
assign n185 = in[23:16] ;
assign bv_8_208_n186 = 8'hd0 ;
assign n187 =  ( n185 ) == ( bv_8_208_n186 )  ;
assign bv_8_112_n188 = 8'h70 ;
assign n189 = in[23:16] ;
assign bv_8_207_n190 = 8'hcf ;
assign n191 =  ( n189 ) == ( bv_8_207_n190 )  ;
assign bv_8_138_n192 = 8'h8a ;
assign n193 = in[23:16] ;
assign n194 =  ( n193 ) == ( bv_8_206_n83 )  ;
assign bv_8_139_n195 = 8'h8b ;
assign n196 = in[23:16] ;
assign bv_8_205_n197 = 8'hcd ;
assign n198 =  ( n196 ) == ( bv_8_205_n197 )  ;
assign bv_8_189_n199 = 8'hbd ;
assign n200 = in[23:16] ;
assign bv_8_204_n201 = 8'hcc ;
assign n202 =  ( n200 ) == ( bv_8_204_n201 )  ;
assign bv_8_75_n203 = 8'h4b ;
assign n204 = in[23:16] ;
assign bv_8_203_n205 = 8'hcb ;
assign n206 =  ( n204 ) == ( bv_8_203_n205 )  ;
assign bv_8_31_n207 = 8'h1f ;
assign n208 = in[23:16] ;
assign bv_8_202_n209 = 8'hca ;
assign n210 =  ( n208 ) == ( bv_8_202_n209 )  ;
assign bv_8_116_n211 = 8'h74 ;
assign n212 = in[23:16] ;
assign bv_8_201_n213 = 8'hc9 ;
assign n214 =  ( n212 ) == ( bv_8_201_n213 )  ;
assign n215 = in[23:16] ;
assign bv_8_200_n216 = 8'hc8 ;
assign n217 =  ( n215 ) == ( bv_8_200_n216 )  ;
assign n218 = in[23:16] ;
assign bv_8_199_n219 = 8'hc7 ;
assign n220 =  ( n218 ) == ( bv_8_199_n219 )  ;
assign bv_8_198_n221 = 8'hc6 ;
assign n222 = in[23:16] ;
assign n223 =  ( n222 ) == ( bv_8_198_n221 )  ;
assign bv_8_180_n224 = 8'hb4 ;
assign n225 = in[23:16] ;
assign bv_8_197_n226 = 8'hc5 ;
assign n227 =  ( n225 ) == ( bv_8_197_n226 )  ;
assign bv_8_166_n228 = 8'ha6 ;
assign n229 = in[23:16] ;
assign bv_8_196_n230 = 8'hc4 ;
assign n231 =  ( n229 ) == ( bv_8_196_n230 )  ;
assign bv_8_28_n232 = 8'h1c ;
assign n233 = in[23:16] ;
assign bv_8_195_n234 = 8'hc3 ;
assign n235 =  ( n233 ) == ( bv_8_195_n234 )  ;
assign bv_8_46_n236 = 8'h2e ;
assign n237 = in[23:16] ;
assign bv_8_194_n238 = 8'hc2 ;
assign n239 =  ( n237 ) == ( bv_8_194_n238 )  ;
assign bv_8_37_n240 = 8'h25 ;
assign n241 = in[23:16] ;
assign n242 =  ( n241 ) == ( bv_8_193_n138 )  ;
assign bv_8_120_n243 = 8'h78 ;
assign n244 = in[23:16] ;
assign bv_8_192_n245 = 8'hc0 ;
assign n246 =  ( n244 ) == ( bv_8_192_n245 )  ;
assign bv_8_186_n247 = 8'hba ;
assign n248 = in[23:16] ;
assign n249 =  ( n248 ) == ( bv_8_191_n51 )  ;
assign bv_8_8_n250 = 8'h8 ;
assign n251 = in[23:16] ;
assign bv_8_190_n252 = 8'hbe ;
assign n253 =  ( n251 ) == ( bv_8_190_n252 )  ;
assign bv_8_174_n254 = 8'hae ;
assign n255 = in[23:16] ;
assign n256 =  ( n255 ) == ( bv_8_189_n199 )  ;
assign bv_8_122_n257 = 8'h7a ;
assign n258 = in[23:16] ;
assign bv_8_188_n259 = 8'hbc ;
assign n260 =  ( n258 ) == ( bv_8_188_n259 )  ;
assign bv_8_101_n261 = 8'h65 ;
assign n262 = in[23:16] ;
assign n263 =  ( n262 ) == ( bv_8_187_n11 )  ;
assign n264 = in[23:16] ;
assign n265 =  ( n264 ) == ( bv_8_186_n247 )  ;
assign n266 = in[23:16] ;
assign n267 =  ( n266 ) == ( bv_8_185_n146 )  ;
assign bv_8_86_n268 = 8'h56 ;
assign n269 = in[23:16] ;
assign bv_8_184_n270 = 8'hb8 ;
assign n271 =  ( n269 ) == ( bv_8_184_n270 )  ;
assign bv_8_108_n272 = 8'h6c ;
assign n273 = in[23:16] ;
assign bv_8_183_n274 = 8'hb7 ;
assign n275 =  ( n273 ) == ( bv_8_183_n274 )  ;
assign bv_8_169_n276 = 8'ha9 ;
assign n277 = in[23:16] ;
assign bv_8_182_n278 = 8'hb6 ;
assign n279 =  ( n277 ) == ( bv_8_182_n278 )  ;
assign bv_8_78_n280 = 8'h4e ;
assign n281 = in[23:16] ;
assign n282 =  ( n281 ) == ( bv_8_181_n180 )  ;
assign n283 = in[23:16] ;
assign n284 =  ( n283 ) == ( bv_8_180_n224 )  ;
assign bv_8_141_n285 = 8'h8d ;
assign n286 = in[23:16] ;
assign bv_8_179_n287 = 8'hb3 ;
assign n288 =  ( n286 ) == ( bv_8_179_n287 )  ;
assign bv_8_109_n289 = 8'h6d ;
assign n290 = in[23:16] ;
assign bv_8_178_n291 = 8'hb2 ;
assign n292 =  ( n290 ) == ( bv_8_178_n291 )  ;
assign bv_8_55_n293 = 8'h37 ;
assign n294 = in[23:16] ;
assign bv_8_177_n295 = 8'hb1 ;
assign n296 =  ( n294 ) == ( bv_8_177_n295 )  ;
assign n297 = in[23:16] ;
assign n298 =  ( n297 ) == ( bv_8_176_n19 )  ;
assign n299 = in[23:16] ;
assign bv_8_175_n300 = 8'haf ;
assign n301 =  ( n299 ) == ( bv_8_175_n300 )  ;
assign bv_8_121_n302 = 8'h79 ;
assign n303 = in[23:16] ;
assign n304 =  ( n303 ) == ( bv_8_174_n254 )  ;
assign n305 = in[23:16] ;
assign bv_8_173_n306 = 8'had ;
assign n307 =  ( n305 ) == ( bv_8_173_n306 )  ;
assign bv_8_149_n308 = 8'h95 ;
assign n309 = in[23:16] ;
assign bv_8_172_n310 = 8'hac ;
assign n311 =  ( n309 ) == ( bv_8_172_n310 )  ;
assign bv_8_145_n312 = 8'h91 ;
assign n313 = in[23:16] ;
assign bv_8_171_n314 = 8'hab ;
assign n315 =  ( n313 ) == ( bv_8_171_n314 )  ;
assign bv_8_98_n316 = 8'h62 ;
assign n317 = in[23:16] ;
assign bv_8_170_n318 = 8'haa ;
assign n319 =  ( n317 ) == ( bv_8_170_n318 )  ;
assign n320 = in[23:16] ;
assign n321 =  ( n320 ) == ( bv_8_169_n276 )  ;
assign n322 = in[23:16] ;
assign bv_8_168_n323 = 8'ha8 ;
assign n324 =  ( n322 ) == ( bv_8_168_n323 )  ;
assign n325 = in[23:16] ;
assign bv_8_167_n326 = 8'ha7 ;
assign n327 =  ( n325 ) == ( bv_8_167_n326 )  ;
assign bv_8_92_n328 = 8'h5c ;
assign n329 = in[23:16] ;
assign n330 =  ( n329 ) == ( bv_8_166_n228 )  ;
assign bv_8_36_n331 = 8'h24 ;
assign n332 = in[23:16] ;
assign bv_8_165_n333 = 8'ha5 ;
assign n334 =  ( n332 ) == ( bv_8_165_n333 )  ;
assign bv_8_6_n335 = 8'h6 ;
assign n336 = in[23:16] ;
assign bv_8_164_n337 = 8'ha4 ;
assign n338 =  ( n336 ) == ( bv_8_164_n337 )  ;
assign bv_8_73_n339 = 8'h49 ;
assign n340 = in[23:16] ;
assign bv_8_163_n341 = 8'ha3 ;
assign n342 =  ( n340 ) == ( bv_8_163_n341 )  ;
assign bv_8_10_n343 = 8'ha ;
assign n344 = in[23:16] ;
assign bv_8_162_n345 = 8'ha2 ;
assign n346 =  ( n344 ) == ( bv_8_162_n345 )  ;
assign bv_8_58_n347 = 8'h3a ;
assign n348 = in[23:16] ;
assign n349 =  ( n348 ) == ( bv_8_161_n63 )  ;
assign bv_8_50_n350 = 8'h32 ;
assign n351 = in[23:16] ;
assign bv_8_160_n352 = 8'ha0 ;
assign n353 =  ( n351 ) == ( bv_8_160_n352 )  ;
assign n354 = in[23:16] ;
assign bv_8_159_n355 = 8'h9f ;
assign n356 =  ( n354 ) == ( bv_8_159_n355 )  ;
assign n357 = in[23:16] ;
assign n358 =  ( n357 ) == ( bv_8_158_n130 )  ;
assign bv_8_11_n359 = 8'hb ;
assign n360 = in[23:16] ;
assign bv_8_157_n361 = 8'h9d ;
assign n362 =  ( n360 ) == ( bv_8_157_n361 )  ;
assign bv_8_94_n363 = 8'h5e ;
assign n364 = in[23:16] ;
assign bv_8_156_n365 = 8'h9c ;
assign n366 =  ( n364 ) == ( bv_8_156_n365 )  ;
assign n367 = in[23:16] ;
assign n368 =  ( n367 ) == ( bv_8_155_n98 )  ;
assign bv_8_20_n369 = 8'h14 ;
assign n370 = in[23:16] ;
assign bv_8_154_n371 = 8'h9a ;
assign n372 =  ( n370 ) == ( bv_8_154_n371 )  ;
assign n373 = in[23:16] ;
assign n374 =  ( n373 ) == ( bv_8_153_n31 )  ;
assign n375 = in[23:16] ;
assign n376 =  ( n375 ) == ( bv_8_152_n121 )  ;
assign bv_8_70_n377 = 8'h46 ;
assign n378 = in[23:16] ;
assign bv_8_151_n379 = 8'h97 ;
assign n380 =  ( n378 ) == ( bv_8_151_n379 )  ;
assign bv_8_136_n381 = 8'h88 ;
assign n382 = in[23:16] ;
assign bv_8_150_n383 = 8'h96 ;
assign n384 =  ( n382 ) == ( bv_8_150_n383 )  ;
assign bv_8_144_n385 = 8'h90 ;
assign n386 = in[23:16] ;
assign n387 =  ( n386 ) == ( bv_8_149_n308 )  ;
assign bv_8_42_n388 = 8'h2a ;
assign n389 = in[23:16] ;
assign n390 =  ( n389 ) == ( bv_8_148_n102 )  ;
assign bv_8_34_n391 = 8'h22 ;
assign n392 = in[23:16] ;
assign bv_8_147_n393 = 8'h93 ;
assign n394 =  ( n392 ) == ( bv_8_147_n393 )  ;
assign n395 = in[23:16] ;
assign bv_8_146_n396 = 8'h92 ;
assign n397 =  ( n395 ) == ( bv_8_146_n396 )  ;
assign bv_8_79_n398 = 8'h4f ;
assign n399 = in[23:16] ;
assign n400 =  ( n399 ) == ( bv_8_145_n312 )  ;
assign bv_8_129_n401 = 8'h81 ;
assign n402 = in[23:16] ;
assign n403 =  ( n402 ) == ( bv_8_144_n385 )  ;
assign bv_8_96_n404 = 8'h60 ;
assign n405 = in[23:16] ;
assign bv_8_143_n406 = 8'h8f ;
assign n407 =  ( n405 ) == ( bv_8_143_n406 )  ;
assign bv_8_115_n408 = 8'h73 ;
assign n409 = in[23:16] ;
assign n410 =  ( n409 ) == ( bv_8_142_n105 )  ;
assign bv_8_25_n411 = 8'h19 ;
assign n412 = in[23:16] ;
assign n413 =  ( n412 ) == ( bv_8_141_n285 )  ;
assign bv_8_93_n414 = 8'h5d ;
assign n415 = in[23:16] ;
assign n416 =  ( n415 ) == ( bv_8_140_n67 )  ;
assign bv_8_100_n417 = 8'h64 ;
assign n418 = in[23:16] ;
assign n419 =  ( n418 ) == ( bv_8_139_n195 )  ;
assign bv_8_61_n420 = 8'h3d ;
assign n421 = in[23:16] ;
assign n422 =  ( n421 ) == ( bv_8_138_n192 )  ;
assign bv_8_126_n423 = 8'h7e ;
assign n424 = in[23:16] ;
assign n425 =  ( n424 ) == ( bv_8_137_n59 )  ;
assign n426 = in[23:16] ;
assign n427 =  ( n426 ) == ( bv_8_136_n381 )  ;
assign n428 = in[23:16] ;
assign n429 =  ( n428 ) == ( bv_8_135_n91 )  ;
assign bv_8_23_n430 = 8'h17 ;
assign n431 = in[23:16] ;
assign n432 =  ( n431 ) == ( bv_8_134_n142 )  ;
assign bv_8_68_n433 = 8'h44 ;
assign n434 = in[23:16] ;
assign bv_8_133_n435 = 8'h85 ;
assign n436 =  ( n434 ) == ( bv_8_133_n435 )  ;
assign n437 = in[23:16] ;
assign bv_8_132_n438 = 8'h84 ;
assign n439 =  ( n437 ) == ( bv_8_132_n438 )  ;
assign bv_8_95_n440 = 8'h5f ;
assign n441 = in[23:16] ;
assign bv_8_131_n442 = 8'h83 ;
assign n443 =  ( n441 ) == ( bv_8_131_n442 )  ;
assign n444 = in[23:16] ;
assign bv_8_130_n445 = 8'h82 ;
assign n446 =  ( n444 ) == ( bv_8_130_n445 )  ;
assign bv_8_19_n447 = 8'h13 ;
assign n448 = in[23:16] ;
assign n449 =  ( n448 ) == ( bv_8_129_n401 )  ;
assign bv_8_12_n450 = 8'hc ;
assign n451 = in[23:16] ;
assign bv_8_128_n452 = 8'h80 ;
assign n453 =  ( n451 ) == ( bv_8_128_n452 )  ;
assign n454 = in[23:16] ;
assign bv_8_127_n455 = 8'h7f ;
assign n456 =  ( n454 ) == ( bv_8_127_n455 )  ;
assign n457 = in[23:16] ;
assign n458 =  ( n457 ) == ( bv_8_126_n423 )  ;
assign n459 = in[23:16] ;
assign bv_8_125_n460 = 8'h7d ;
assign n461 =  ( n459 ) == ( bv_8_125_n460 )  ;
assign n462 = in[23:16] ;
assign bv_8_124_n463 = 8'h7c ;
assign n464 =  ( n462 ) == ( bv_8_124_n463 )  ;
assign bv_8_16_n465 = 8'h10 ;
assign n466 = in[23:16] ;
assign bv_8_123_n467 = 8'h7b ;
assign n468 =  ( n466 ) == ( bv_8_123_n467 )  ;
assign bv_8_33_n469 = 8'h21 ;
assign n470 = in[23:16] ;
assign n471 =  ( n470 ) == ( bv_8_122_n257 )  ;
assign n472 = in[23:16] ;
assign n473 =  ( n472 ) == ( bv_8_121_n302 )  ;
assign n474 = in[23:16] ;
assign n475 =  ( n474 ) == ( bv_8_120_n243 )  ;
assign n476 = in[23:16] ;
assign bv_8_119_n477 = 8'h77 ;
assign n478 =  ( n476 ) == ( bv_8_119_n477 )  ;
assign n479 = in[23:16] ;
assign bv_8_118_n480 = 8'h76 ;
assign n481 =  ( n479 ) == ( bv_8_118_n480 )  ;
assign bv_8_56_n482 = 8'h38 ;
assign n483 = in[23:16] ;
assign bv_8_117_n484 = 8'h75 ;
assign n485 =  ( n483 ) == ( bv_8_117_n484 )  ;
assign n486 = in[23:16] ;
assign n487 =  ( n486 ) == ( bv_8_116_n211 )  ;
assign n488 = in[23:16] ;
assign n489 =  ( n488 ) == ( bv_8_115_n408 )  ;
assign n490 = in[23:16] ;
assign bv_8_114_n491 = 8'h72 ;
assign n492 =  ( n490 ) == ( bv_8_114_n491 )  ;
assign bv_8_64_n493 = 8'h40 ;
assign n494 = in[23:16] ;
assign bv_8_113_n495 = 8'h71 ;
assign n496 =  ( n494 ) == ( bv_8_113_n495 )  ;
assign n497 = in[23:16] ;
assign n498 =  ( n497 ) == ( bv_8_112_n188 )  ;
assign bv_8_81_n499 = 8'h51 ;
assign n500 = in[23:16] ;
assign bv_8_111_n501 = 8'h6f ;
assign n502 =  ( n500 ) == ( bv_8_111_n501 )  ;
assign n503 = in[23:16] ;
assign bv_8_110_n504 = 8'h6e ;
assign n505 =  ( n503 ) == ( bv_8_110_n504 )  ;
assign n506 = in[23:16] ;
assign n507 =  ( n506 ) == ( bv_8_109_n289 )  ;
assign bv_8_60_n508 = 8'h3c ;
assign n509 = in[23:16] ;
assign n510 =  ( n509 ) == ( bv_8_108_n272 )  ;
assign bv_8_80_n511 = 8'h50 ;
assign n512 = in[23:16] ;
assign bv_8_107_n513 = 8'h6b ;
assign n514 =  ( n512 ) == ( bv_8_107_n513 )  ;
assign n515 = in[23:16] ;
assign bv_8_106_n516 = 8'h6a ;
assign n517 =  ( n515 ) == ( bv_8_106_n516 )  ;
assign bv_8_2_n518 = 8'h2 ;
assign n519 = in[23:16] ;
assign n520 =  ( n519 ) == ( bv_8_105_n113 )  ;
assign n521 = in[23:16] ;
assign n522 =  ( n521 ) == ( bv_8_104_n39 )  ;
assign bv_8_69_n523 = 8'h45 ;
assign n524 = in[23:16] ;
assign bv_8_103_n525 = 8'h67 ;
assign n526 =  ( n524 ) == ( bv_8_103_n525 )  ;
assign n527 = in[23:16] ;
assign n528 =  ( n527 ) == ( bv_8_102_n176 )  ;
assign bv_8_51_n529 = 8'h33 ;
assign n530 = in[23:16] ;
assign n531 =  ( n530 ) == ( bv_8_101_n261 )  ;
assign bv_8_77_n532 = 8'h4d ;
assign n533 = in[23:16] ;
assign n534 =  ( n533 ) == ( bv_8_100_n417 )  ;
assign bv_8_67_n535 = 8'h43 ;
assign n536 = in[23:16] ;
assign bv_8_99_n537 = 8'h63 ;
assign n538 =  ( n536 ) == ( bv_8_99_n537 )  ;
assign n539 = in[23:16] ;
assign n540 =  ( n539 ) == ( bv_8_98_n316 )  ;
assign n541 = in[23:16] ;
assign n542 =  ( n541 ) == ( bv_8_97_n157 )  ;
assign n543 = in[23:16] ;
assign n544 =  ( n543 ) == ( bv_8_96_n404 )  ;
assign n545 = in[23:16] ;
assign n546 =  ( n545 ) == ( bv_8_95_n440 )  ;
assign n547 = in[23:16] ;
assign n548 =  ( n547 ) == ( bv_8_94_n363 )  ;
assign bv_8_88_n549 = 8'h58 ;
assign n550 = in[23:16] ;
assign n551 =  ( n550 ) == ( bv_8_93_n414 )  ;
assign bv_8_76_n552 = 8'h4c ;
assign n553 = in[23:16] ;
assign n554 =  ( n553 ) == ( bv_8_92_n328 )  ;
assign bv_8_74_n555 = 8'h4a ;
assign n556 = in[23:16] ;
assign bv_8_91_n557 = 8'h5b ;
assign n558 =  ( n556 ) == ( bv_8_91_n557 )  ;
assign bv_8_57_n559 = 8'h39 ;
assign n560 = in[23:16] ;
assign bv_8_90_n561 = 8'h5a ;
assign n562 =  ( n560 ) == ( bv_8_90_n561 )  ;
assign n563 = in[23:16] ;
assign bv_8_89_n564 = 8'h59 ;
assign n565 =  ( n563 ) == ( bv_8_89_n564 )  ;
assign n566 = in[23:16] ;
assign n567 =  ( n566 ) == ( bv_8_88_n549 )  ;
assign n568 = in[23:16] ;
assign n569 =  ( n568 ) == ( bv_8_87_n150 )  ;
assign n570 = in[23:16] ;
assign n571 =  ( n570 ) == ( bv_8_86_n268 )  ;
assign n572 = in[23:16] ;
assign n573 =  ( n572 ) == ( bv_8_85_n79 )  ;
assign n574 = in[23:16] ;
assign n575 =  ( n574 ) == ( bv_8_84_n15 )  ;
assign bv_8_32_n576 = 8'h20 ;
assign n577 = in[23:16] ;
assign bv_8_83_n578 = 8'h53 ;
assign n579 =  ( n577 ) == ( bv_8_83_n578 )  ;
assign n580 = in[23:16] ;
assign bv_8_82_n581 = 8'h52 ;
assign n582 =  ( n580 ) == ( bv_8_82_n581 )  ;
assign bv_8_0_n583 = 8'h0 ;
assign n584 = in[23:16] ;
assign n585 =  ( n584 ) == ( bv_8_81_n499 )  ;
assign n586 = in[23:16] ;
assign n587 =  ( n586 ) == ( bv_8_80_n511 )  ;
assign n588 = in[23:16] ;
assign n589 =  ( n588 ) == ( bv_8_79_n398 )  ;
assign n590 = in[23:16] ;
assign n591 =  ( n590 ) == ( bv_8_78_n280 )  ;
assign bv_8_47_n592 = 8'h2f ;
assign n593 = in[23:16] ;
assign n594 =  ( n593 ) == ( bv_8_77_n532 )  ;
assign n595 = in[23:16] ;
assign n596 =  ( n595 ) == ( bv_8_76_n552 )  ;
assign bv_8_41_n597 = 8'h29 ;
assign n598 = in[23:16] ;
assign n599 =  ( n598 ) == ( bv_8_75_n203 )  ;
assign n600 = in[23:16] ;
assign n601 =  ( n600 ) == ( bv_8_74_n555 )  ;
assign n602 = in[23:16] ;
assign n603 =  ( n602 ) == ( bv_8_73_n339 )  ;
assign bv_8_59_n604 = 8'h3b ;
assign n605 = in[23:16] ;
assign n606 =  ( n605 ) == ( bv_8_72_n172 )  ;
assign n607 = in[23:16] ;
assign bv_8_71_n608 = 8'h47 ;
assign n609 =  ( n607 ) == ( bv_8_71_n608 )  ;
assign n610 = in[23:16] ;
assign n611 =  ( n610 ) == ( bv_8_70_n377 )  ;
assign n612 = in[23:16] ;
assign n613 =  ( n612 ) == ( bv_8_69_n523 )  ;
assign n614 = in[23:16] ;
assign n615 =  ( n614 ) == ( bv_8_68_n433 )  ;
assign bv_8_27_n616 = 8'h1b ;
assign n617 = in[23:16] ;
assign n618 =  ( n617 ) == ( bv_8_67_n535 )  ;
assign bv_8_26_n619 = 8'h1a ;
assign n620 = in[23:16] ;
assign n621 =  ( n620 ) == ( bv_8_66_n43 )  ;
assign bv_8_44_n622 = 8'h2c ;
assign n623 = in[23:16] ;
assign n624 =  ( n623 ) == ( bv_8_65_n35 )  ;
assign n625 = in[23:16] ;
assign n626 =  ( n625 ) == ( bv_8_64_n493 )  ;
assign bv_8_9_n627 = 8'h9 ;
assign n628 = in[23:16] ;
assign bv_8_63_n629 = 8'h3f ;
assign n630 =  ( n628 ) == ( bv_8_63_n629 )  ;
assign n631 = in[23:16] ;
assign n632 =  ( n631 ) == ( bv_8_62_n184 )  ;
assign n633 = in[23:16] ;
assign n634 =  ( n633 ) == ( bv_8_61_n420 )  ;
assign bv_8_39_n635 = 8'h27 ;
assign n636 = in[23:16] ;
assign n637 =  ( n636 ) == ( bv_8_60_n508 )  ;
assign n638 = in[23:16] ;
assign n639 =  ( n638 ) == ( bv_8_59_n604 )  ;
assign n640 = in[23:16] ;
assign n641 =  ( n640 ) == ( bv_8_58_n347 )  ;
assign n642 = in[23:16] ;
assign n643 =  ( n642 ) == ( bv_8_57_n559 )  ;
assign bv_8_18_n644 = 8'h12 ;
assign n645 = in[23:16] ;
assign n646 =  ( n645 ) == ( bv_8_56_n482 )  ;
assign bv_8_7_n647 = 8'h7 ;
assign n648 = in[23:16] ;
assign n649 =  ( n648 ) == ( bv_8_55_n293 )  ;
assign n650 = in[23:16] ;
assign bv_8_54_n651 = 8'h36 ;
assign n652 =  ( n650 ) == ( bv_8_54_n651 )  ;
assign bv_8_5_n653 = 8'h5 ;
assign n654 = in[23:16] ;
assign n655 =  ( n654 ) == ( bv_8_53_n153 )  ;
assign n656 = in[23:16] ;
assign bv_8_52_n657 = 8'h34 ;
assign n658 =  ( n656 ) == ( bv_8_52_n657 )  ;
assign bv_8_24_n659 = 8'h18 ;
assign n660 = in[23:16] ;
assign n661 =  ( n660 ) == ( bv_8_51_n529 )  ;
assign n662 = in[23:16] ;
assign n663 =  ( n662 ) == ( bv_8_50_n350 )  ;
assign bv_8_35_n664 = 8'h23 ;
assign n665 = in[23:16] ;
assign bv_8_49_n666 = 8'h31 ;
assign n667 =  ( n665 ) == ( bv_8_49_n666 )  ;
assign n668 = in[23:16] ;
assign bv_8_48_n669 = 8'h30 ;
assign n670 =  ( n668 ) == ( bv_8_48_n669 )  ;
assign bv_8_4_n671 = 8'h4 ;
assign n672 = in[23:16] ;
assign n673 =  ( n672 ) == ( bv_8_47_n592 )  ;
assign bv_8_21_n674 = 8'h15 ;
assign n675 = in[23:16] ;
assign n676 =  ( n675 ) == ( bv_8_46_n236 )  ;
assign n677 = in[23:16] ;
assign n678 =  ( n677 ) == ( bv_8_45_n27 )  ;
assign n679 = in[23:16] ;
assign n680 =  ( n679 ) == ( bv_8_44_n622 )  ;
assign n681 = in[23:16] ;
assign bv_8_43_n682 = 8'h2b ;
assign n683 =  ( n681 ) == ( bv_8_43_n682 )  ;
assign n684 = in[23:16] ;
assign n685 =  ( n684 ) == ( bv_8_42_n388 )  ;
assign n686 = in[23:16] ;
assign n687 =  ( n686 ) == ( bv_8_41_n597 )  ;
assign n688 = in[23:16] ;
assign n689 =  ( n688 ) == ( bv_8_40_n75 )  ;
assign n690 = in[23:16] ;
assign n691 =  ( n690 ) == ( bv_8_39_n635 )  ;
assign n692 = in[23:16] ;
assign bv_8_38_n693 = 8'h26 ;
assign n694 =  ( n692 ) == ( bv_8_38_n693 )  ;
assign n695 = in[23:16] ;
assign n696 =  ( n695 ) == ( bv_8_37_n240 )  ;
assign n697 = in[23:16] ;
assign n698 =  ( n697 ) == ( bv_8_36_n331 )  ;
assign n699 = in[23:16] ;
assign n700 =  ( n699 ) == ( bv_8_35_n664 )  ;
assign n701 = in[23:16] ;
assign n702 =  ( n701 ) == ( bv_8_34_n391 )  ;
assign n703 = in[23:16] ;
assign n704 =  ( n703 ) == ( bv_8_33_n469 )  ;
assign n705 = in[23:16] ;
assign n706 =  ( n705 ) == ( bv_8_32_n576 )  ;
assign n707 = in[23:16] ;
assign n708 =  ( n707 ) == ( bv_8_31_n207 )  ;
assign n709 = in[23:16] ;
assign n710 =  ( n709 ) == ( bv_8_30_n94 )  ;
assign n711 = in[23:16] ;
assign n712 =  ( n711 ) == ( bv_8_29_n134 )  ;
assign n713 = in[23:16] ;
assign n714 =  ( n713 ) == ( bv_8_28_n232 )  ;
assign n715 = in[23:16] ;
assign n716 =  ( n715 ) == ( bv_8_27_n616 )  ;
assign n717 = in[23:16] ;
assign n718 =  ( n717 ) == ( bv_8_26_n619 )  ;
assign n719 = in[23:16] ;
assign n720 =  ( n719 ) == ( bv_8_25_n411 )  ;
assign n721 = in[23:16] ;
assign n722 =  ( n721 ) == ( bv_8_24_n659 )  ;
assign n723 = in[23:16] ;
assign n724 =  ( n723 ) == ( bv_8_23_n430 )  ;
assign n725 = in[23:16] ;
assign n726 =  ( n725 ) == ( bv_8_22_n7 )  ;
assign n727 = in[23:16] ;
assign n728 =  ( n727 ) == ( bv_8_21_n674 )  ;
assign n729 = in[23:16] ;
assign n730 =  ( n729 ) == ( bv_8_20_n369 )  ;
assign n731 = in[23:16] ;
assign n732 =  ( n731 ) == ( bv_8_19_n447 )  ;
assign n733 = in[23:16] ;
assign n734 =  ( n733 ) == ( bv_8_18_n644 )  ;
assign n735 = in[23:16] ;
assign n736 =  ( n735 ) == ( bv_8_17_n117 )  ;
assign n737 = in[23:16] ;
assign n738 =  ( n737 ) == ( bv_8_16_n465 )  ;
assign n739 = in[23:16] ;
assign n740 =  ( n739 ) == ( bv_8_15_n23 )  ;
assign n741 = in[23:16] ;
assign n742 =  ( n741 ) == ( bv_8_14_n161 )  ;
assign n743 = in[23:16] ;
assign n744 =  ( n743 ) == ( bv_8_13_n55 )  ;
assign n745 = in[23:16] ;
assign n746 =  ( n745 ) == ( bv_8_12_n450 )  ;
assign n747 = in[23:16] ;
assign n748 =  ( n747 ) == ( bv_8_11_n359 )  ;
assign n749 = in[23:16] ;
assign n750 =  ( n749 ) == ( bv_8_10_n343 )  ;
assign n751 = in[23:16] ;
assign n752 =  ( n751 ) == ( bv_8_9_n627 )  ;
assign bv_8_1_n753 = 8'h1 ;
assign n754 = in[23:16] ;
assign n755 =  ( n754 ) == ( bv_8_8_n250 )  ;
assign n756 = in[23:16] ;
assign n757 =  ( n756 ) == ( bv_8_7_n647 )  ;
assign n758 = in[23:16] ;
assign n759 =  ( n758 ) == ( bv_8_6_n335 )  ;
assign n760 = in[23:16] ;
assign n761 =  ( n760 ) == ( bv_8_5_n653 )  ;
assign n762 = in[23:16] ;
assign n763 =  ( n762 ) == ( bv_8_4_n671 )  ;
assign n764 = in[23:16] ;
assign n765 =  ( n764 ) == ( bv_8_3_n168 )  ;
assign n766 = in[23:16] ;
assign n767 =  ( n766 ) == ( bv_8_2_n518 )  ;
assign n768 = in[23:16] ;
assign n769 =  ( n768 ) == ( bv_8_1_n753 )  ;
assign n770 = in[23:16] ;
assign n771 =  ( n770 ) == ( bv_8_0_n583 )  ;
assign n772 =  ( n771 ) ? ( bv_8_99_n537 ) : ( bv_8_0_n583 ) ;
assign n773 =  ( n769 ) ? ( bv_8_124_n463 ) : ( n772 ) ;
assign n774 =  ( n767 ) ? ( bv_8_119_n477 ) : ( n773 ) ;
assign n775 =  ( n765 ) ? ( bv_8_123_n467 ) : ( n774 ) ;
assign n776 =  ( n763 ) ? ( bv_8_242_n57 ) : ( n775 ) ;
assign n777 =  ( n761 ) ? ( bv_8_107_n513 ) : ( n776 ) ;
assign n778 =  ( n759 ) ? ( bv_8_111_n501 ) : ( n777 ) ;
assign n779 =  ( n757 ) ? ( bv_8_197_n226 ) : ( n778 ) ;
assign n780 =  ( n755 ) ? ( bv_8_48_n669 ) : ( n779 ) ;
assign n781 =  ( n752 ) ? ( bv_8_1_n753 ) : ( n780 ) ;
assign n782 =  ( n750 ) ? ( bv_8_103_n525 ) : ( n781 ) ;
assign n783 =  ( n748 ) ? ( bv_8_43_n682 ) : ( n782 ) ;
assign n784 =  ( n746 ) ? ( bv_8_254_n9 ) : ( n783 ) ;
assign n785 =  ( n744 ) ? ( bv_8_215_n159 ) : ( n784 ) ;
assign n786 =  ( n742 ) ? ( bv_8_171_n314 ) : ( n785 ) ;
assign n787 =  ( n740 ) ? ( bv_8_118_n480 ) : ( n786 ) ;
assign n788 =  ( n738 ) ? ( bv_8_202_n209 ) : ( n787 ) ;
assign n789 =  ( n736 ) ? ( bv_8_130_n445 ) : ( n788 ) ;
assign n790 =  ( n734 ) ? ( bv_8_201_n213 ) : ( n789 ) ;
assign n791 =  ( n732 ) ? ( bv_8_125_n460 ) : ( n790 ) ;
assign n792 =  ( n730 ) ? ( bv_8_250_n25 ) : ( n791 ) ;
assign n793 =  ( n728 ) ? ( bv_8_89_n564 ) : ( n792 ) ;
assign n794 =  ( n726 ) ? ( bv_8_71_n608 ) : ( n793 ) ;
assign n795 =  ( n724 ) ? ( bv_8_240_n65 ) : ( n794 ) ;
assign n796 =  ( n722 ) ? ( bv_8_173_n306 ) : ( n795 ) ;
assign n797 =  ( n720 ) ? ( bv_8_212_n170 ) : ( n796 ) ;
assign n798 =  ( n718 ) ? ( bv_8_162_n345 ) : ( n797 ) ;
assign n799 =  ( n716 ) ? ( bv_8_175_n300 ) : ( n798 ) ;
assign n800 =  ( n714 ) ? ( bv_8_156_n365 ) : ( n799 ) ;
assign n801 =  ( n712 ) ? ( bv_8_164_n337 ) : ( n800 ) ;
assign n802 =  ( n710 ) ? ( bv_8_114_n491 ) : ( n801 ) ;
assign n803 =  ( n708 ) ? ( bv_8_192_n245 ) : ( n802 ) ;
assign n804 =  ( n706 ) ? ( bv_8_183_n274 ) : ( n803 ) ;
assign n805 =  ( n704 ) ? ( bv_8_253_n13 ) : ( n804 ) ;
assign n806 =  ( n702 ) ? ( bv_8_147_n393 ) : ( n805 ) ;
assign n807 =  ( n700 ) ? ( bv_8_38_n693 ) : ( n806 ) ;
assign n808 =  ( n698 ) ? ( bv_8_54_n651 ) : ( n807 ) ;
assign n809 =  ( n696 ) ? ( bv_8_63_n629 ) : ( n808 ) ;
assign n810 =  ( n694 ) ? ( bv_8_247_n37 ) : ( n809 ) ;
assign n811 =  ( n691 ) ? ( bv_8_204_n201 ) : ( n810 ) ;
assign n812 =  ( n689 ) ? ( bv_8_52_n657 ) : ( n811 ) ;
assign n813 =  ( n687 ) ? ( bv_8_165_n333 ) : ( n812 ) ;
assign n814 =  ( n685 ) ? ( bv_8_229_n107 ) : ( n813 ) ;
assign n815 =  ( n683 ) ? ( bv_8_241_n61 ) : ( n814 ) ;
assign n816 =  ( n680 ) ? ( bv_8_113_n495 ) : ( n815 ) ;
assign n817 =  ( n678 ) ? ( bv_8_216_n155 ) : ( n816 ) ;
assign n818 =  ( n676 ) ? ( bv_8_49_n666 ) : ( n817 ) ;
assign n819 =  ( n673 ) ? ( bv_8_21_n674 ) : ( n818 ) ;
assign n820 =  ( n670 ) ? ( bv_8_4_n671 ) : ( n819 ) ;
assign n821 =  ( n667 ) ? ( bv_8_199_n219 ) : ( n820 ) ;
assign n822 =  ( n663 ) ? ( bv_8_35_n664 ) : ( n821 ) ;
assign n823 =  ( n661 ) ? ( bv_8_195_n234 ) : ( n822 ) ;
assign n824 =  ( n658 ) ? ( bv_8_24_n659 ) : ( n823 ) ;
assign n825 =  ( n655 ) ? ( bv_8_150_n383 ) : ( n824 ) ;
assign n826 =  ( n652 ) ? ( bv_8_5_n653 ) : ( n825 ) ;
assign n827 =  ( n649 ) ? ( bv_8_154_n371 ) : ( n826 ) ;
assign n828 =  ( n646 ) ? ( bv_8_7_n647 ) : ( n827 ) ;
assign n829 =  ( n643 ) ? ( bv_8_18_n644 ) : ( n828 ) ;
assign n830 =  ( n641 ) ? ( bv_8_128_n452 ) : ( n829 ) ;
assign n831 =  ( n639 ) ? ( bv_8_226_n119 ) : ( n830 ) ;
assign n832 =  ( n637 ) ? ( bv_8_235_n85 ) : ( n831 ) ;
assign n833 =  ( n634 ) ? ( bv_8_39_n635 ) : ( n832 ) ;
assign n834 =  ( n632 ) ? ( bv_8_178_n291 ) : ( n833 ) ;
assign n835 =  ( n630 ) ? ( bv_8_117_n484 ) : ( n834 ) ;
assign n836 =  ( n626 ) ? ( bv_8_9_n627 ) : ( n835 ) ;
assign n837 =  ( n624 ) ? ( bv_8_131_n442 ) : ( n836 ) ;
assign n838 =  ( n621 ) ? ( bv_8_44_n622 ) : ( n837 ) ;
assign n839 =  ( n618 ) ? ( bv_8_26_n619 ) : ( n838 ) ;
assign n840 =  ( n615 ) ? ( bv_8_27_n616 ) : ( n839 ) ;
assign n841 =  ( n613 ) ? ( bv_8_110_n504 ) : ( n840 ) ;
assign n842 =  ( n611 ) ? ( bv_8_90_n561 ) : ( n841 ) ;
assign n843 =  ( n609 ) ? ( bv_8_160_n352 ) : ( n842 ) ;
assign n844 =  ( n606 ) ? ( bv_8_82_n581 ) : ( n843 ) ;
assign n845 =  ( n603 ) ? ( bv_8_59_n604 ) : ( n844 ) ;
assign n846 =  ( n601 ) ? ( bv_8_214_n163 ) : ( n845 ) ;
assign n847 =  ( n599 ) ? ( bv_8_179_n287 ) : ( n846 ) ;
assign n848 =  ( n596 ) ? ( bv_8_41_n597 ) : ( n847 ) ;
assign n849 =  ( n594 ) ? ( bv_8_227_n115 ) : ( n848 ) ;
assign n850 =  ( n591 ) ? ( bv_8_47_n592 ) : ( n849 ) ;
assign n851 =  ( n589 ) ? ( bv_8_132_n438 ) : ( n850 ) ;
assign n852 =  ( n587 ) ? ( bv_8_83_n578 ) : ( n851 ) ;
assign n853 =  ( n585 ) ? ( bv_8_209_n182 ) : ( n852 ) ;
assign n854 =  ( n582 ) ? ( bv_8_0_n583 ) : ( n853 ) ;
assign n855 =  ( n579 ) ? ( bv_8_237_n77 ) : ( n854 ) ;
assign n856 =  ( n575 ) ? ( bv_8_32_n576 ) : ( n855 ) ;
assign n857 =  ( n573 ) ? ( bv_8_252_n17 ) : ( n856 ) ;
assign n858 =  ( n571 ) ? ( bv_8_177_n295 ) : ( n857 ) ;
assign n859 =  ( n569 ) ? ( bv_8_91_n557 ) : ( n858 ) ;
assign n860 =  ( n567 ) ? ( bv_8_106_n516 ) : ( n859 ) ;
assign n861 =  ( n565 ) ? ( bv_8_203_n205 ) : ( n860 ) ;
assign n862 =  ( n562 ) ? ( bv_8_190_n252 ) : ( n861 ) ;
assign n863 =  ( n558 ) ? ( bv_8_57_n559 ) : ( n862 ) ;
assign n864 =  ( n554 ) ? ( bv_8_74_n555 ) : ( n863 ) ;
assign n865 =  ( n551 ) ? ( bv_8_76_n552 ) : ( n864 ) ;
assign n866 =  ( n548 ) ? ( bv_8_88_n549 ) : ( n865 ) ;
assign n867 =  ( n546 ) ? ( bv_8_207_n190 ) : ( n866 ) ;
assign n868 =  ( n544 ) ? ( bv_8_208_n186 ) : ( n867 ) ;
assign n869 =  ( n542 ) ? ( bv_8_239_n69 ) : ( n868 ) ;
assign n870 =  ( n540 ) ? ( bv_8_170_n318 ) : ( n869 ) ;
assign n871 =  ( n538 ) ? ( bv_8_251_n21 ) : ( n870 ) ;
assign n872 =  ( n534 ) ? ( bv_8_67_n535 ) : ( n871 ) ;
assign n873 =  ( n531 ) ? ( bv_8_77_n532 ) : ( n872 ) ;
assign n874 =  ( n528 ) ? ( bv_8_51_n529 ) : ( n873 ) ;
assign n875 =  ( n526 ) ? ( bv_8_133_n435 ) : ( n874 ) ;
assign n876 =  ( n522 ) ? ( bv_8_69_n523 ) : ( n875 ) ;
assign n877 =  ( n520 ) ? ( bv_8_249_n29 ) : ( n876 ) ;
assign n878 =  ( n517 ) ? ( bv_8_2_n518 ) : ( n877 ) ;
assign n879 =  ( n514 ) ? ( bv_8_127_n455 ) : ( n878 ) ;
assign n880 =  ( n510 ) ? ( bv_8_80_n511 ) : ( n879 ) ;
assign n881 =  ( n507 ) ? ( bv_8_60_n508 ) : ( n880 ) ;
assign n882 =  ( n505 ) ? ( bv_8_159_n355 ) : ( n881 ) ;
assign n883 =  ( n502 ) ? ( bv_8_168_n323 ) : ( n882 ) ;
assign n884 =  ( n498 ) ? ( bv_8_81_n499 ) : ( n883 ) ;
assign n885 =  ( n496 ) ? ( bv_8_163_n341 ) : ( n884 ) ;
assign n886 =  ( n492 ) ? ( bv_8_64_n493 ) : ( n885 ) ;
assign n887 =  ( n489 ) ? ( bv_8_143_n406 ) : ( n886 ) ;
assign n888 =  ( n487 ) ? ( bv_8_146_n396 ) : ( n887 ) ;
assign n889 =  ( n485 ) ? ( bv_8_157_n361 ) : ( n888 ) ;
assign n890 =  ( n481 ) ? ( bv_8_56_n482 ) : ( n889 ) ;
assign n891 =  ( n478 ) ? ( bv_8_245_n45 ) : ( n890 ) ;
assign n892 =  ( n475 ) ? ( bv_8_188_n259 ) : ( n891 ) ;
assign n893 =  ( n473 ) ? ( bv_8_182_n278 ) : ( n892 ) ;
assign n894 =  ( n471 ) ? ( bv_8_218_n148 ) : ( n893 ) ;
assign n895 =  ( n468 ) ? ( bv_8_33_n469 ) : ( n894 ) ;
assign n896 =  ( n464 ) ? ( bv_8_16_n465 ) : ( n895 ) ;
assign n897 =  ( n461 ) ? ( bv_8_255_n5 ) : ( n896 ) ;
assign n898 =  ( n458 ) ? ( bv_8_243_n53 ) : ( n897 ) ;
assign n899 =  ( n456 ) ? ( bv_8_210_n178 ) : ( n898 ) ;
assign n900 =  ( n453 ) ? ( bv_8_205_n197 ) : ( n899 ) ;
assign n901 =  ( n449 ) ? ( bv_8_12_n450 ) : ( n900 ) ;
assign n902 =  ( n446 ) ? ( bv_8_19_n447 ) : ( n901 ) ;
assign n903 =  ( n443 ) ? ( bv_8_236_n81 ) : ( n902 ) ;
assign n904 =  ( n439 ) ? ( bv_8_95_n440 ) : ( n903 ) ;
assign n905 =  ( n436 ) ? ( bv_8_151_n379 ) : ( n904 ) ;
assign n906 =  ( n432 ) ? ( bv_8_68_n433 ) : ( n905 ) ;
assign n907 =  ( n429 ) ? ( bv_8_23_n430 ) : ( n906 ) ;
assign n908 =  ( n427 ) ? ( bv_8_196_n230 ) : ( n907 ) ;
assign n909 =  ( n425 ) ? ( bv_8_167_n326 ) : ( n908 ) ;
assign n910 =  ( n422 ) ? ( bv_8_126_n423 ) : ( n909 ) ;
assign n911 =  ( n419 ) ? ( bv_8_61_n420 ) : ( n910 ) ;
assign n912 =  ( n416 ) ? ( bv_8_100_n417 ) : ( n911 ) ;
assign n913 =  ( n413 ) ? ( bv_8_93_n414 ) : ( n912 ) ;
assign n914 =  ( n410 ) ? ( bv_8_25_n411 ) : ( n913 ) ;
assign n915 =  ( n407 ) ? ( bv_8_115_n408 ) : ( n914 ) ;
assign n916 =  ( n403 ) ? ( bv_8_96_n404 ) : ( n915 ) ;
assign n917 =  ( n400 ) ? ( bv_8_129_n401 ) : ( n916 ) ;
assign n918 =  ( n397 ) ? ( bv_8_79_n398 ) : ( n917 ) ;
assign n919 =  ( n394 ) ? ( bv_8_220_n140 ) : ( n918 ) ;
assign n920 =  ( n390 ) ? ( bv_8_34_n391 ) : ( n919 ) ;
assign n921 =  ( n387 ) ? ( bv_8_42_n388 ) : ( n920 ) ;
assign n922 =  ( n384 ) ? ( bv_8_144_n385 ) : ( n921 ) ;
assign n923 =  ( n380 ) ? ( bv_8_136_n381 ) : ( n922 ) ;
assign n924 =  ( n376 ) ? ( bv_8_70_n377 ) : ( n923 ) ;
assign n925 =  ( n374 ) ? ( bv_8_238_n73 ) : ( n924 ) ;
assign n926 =  ( n372 ) ? ( bv_8_184_n270 ) : ( n925 ) ;
assign n927 =  ( n368 ) ? ( bv_8_20_n369 ) : ( n926 ) ;
assign n928 =  ( n366 ) ? ( bv_8_222_n132 ) : ( n927 ) ;
assign n929 =  ( n362 ) ? ( bv_8_94_n363 ) : ( n928 ) ;
assign n930 =  ( n358 ) ? ( bv_8_11_n359 ) : ( n929 ) ;
assign n931 =  ( n356 ) ? ( bv_8_219_n144 ) : ( n930 ) ;
assign n932 =  ( n353 ) ? ( bv_8_224_n126 ) : ( n931 ) ;
assign n933 =  ( n349 ) ? ( bv_8_50_n350 ) : ( n932 ) ;
assign n934 =  ( n346 ) ? ( bv_8_58_n347 ) : ( n933 ) ;
assign n935 =  ( n342 ) ? ( bv_8_10_n343 ) : ( n934 ) ;
assign n936 =  ( n338 ) ? ( bv_8_73_n339 ) : ( n935 ) ;
assign n937 =  ( n334 ) ? ( bv_8_6_n335 ) : ( n936 ) ;
assign n938 =  ( n330 ) ? ( bv_8_36_n331 ) : ( n937 ) ;
assign n939 =  ( n327 ) ? ( bv_8_92_n328 ) : ( n938 ) ;
assign n940 =  ( n324 ) ? ( bv_8_194_n238 ) : ( n939 ) ;
assign n941 =  ( n321 ) ? ( bv_8_211_n174 ) : ( n940 ) ;
assign n942 =  ( n319 ) ? ( bv_8_172_n310 ) : ( n941 ) ;
assign n943 =  ( n315 ) ? ( bv_8_98_n316 ) : ( n942 ) ;
assign n944 =  ( n311 ) ? ( bv_8_145_n312 ) : ( n943 ) ;
assign n945 =  ( n307 ) ? ( bv_8_149_n308 ) : ( n944 ) ;
assign n946 =  ( n304 ) ? ( bv_8_228_n111 ) : ( n945 ) ;
assign n947 =  ( n301 ) ? ( bv_8_121_n302 ) : ( n946 ) ;
assign n948 =  ( n298 ) ? ( bv_8_231_n100 ) : ( n947 ) ;
assign n949 =  ( n296 ) ? ( bv_8_200_n216 ) : ( n948 ) ;
assign n950 =  ( n292 ) ? ( bv_8_55_n293 ) : ( n949 ) ;
assign n951 =  ( n288 ) ? ( bv_8_109_n289 ) : ( n950 ) ;
assign n952 =  ( n284 ) ? ( bv_8_141_n285 ) : ( n951 ) ;
assign n953 =  ( n282 ) ? ( bv_8_213_n166 ) : ( n952 ) ;
assign n954 =  ( n279 ) ? ( bv_8_78_n280 ) : ( n953 ) ;
assign n955 =  ( n275 ) ? ( bv_8_169_n276 ) : ( n954 ) ;
assign n956 =  ( n271 ) ? ( bv_8_108_n272 ) : ( n955 ) ;
assign n957 =  ( n267 ) ? ( bv_8_86_n268 ) : ( n956 ) ;
assign n958 =  ( n265 ) ? ( bv_8_244_n49 ) : ( n957 ) ;
assign n959 =  ( n263 ) ? ( bv_8_234_n89 ) : ( n958 ) ;
assign n960 =  ( n260 ) ? ( bv_8_101_n261 ) : ( n959 ) ;
assign n961 =  ( n256 ) ? ( bv_8_122_n257 ) : ( n960 ) ;
assign n962 =  ( n253 ) ? ( bv_8_174_n254 ) : ( n961 ) ;
assign n963 =  ( n249 ) ? ( bv_8_8_n250 ) : ( n962 ) ;
assign n964 =  ( n246 ) ? ( bv_8_186_n247 ) : ( n963 ) ;
assign n965 =  ( n242 ) ? ( bv_8_120_n243 ) : ( n964 ) ;
assign n966 =  ( n239 ) ? ( bv_8_37_n240 ) : ( n965 ) ;
assign n967 =  ( n235 ) ? ( bv_8_46_n236 ) : ( n966 ) ;
assign n968 =  ( n231 ) ? ( bv_8_28_n232 ) : ( n967 ) ;
assign n969 =  ( n227 ) ? ( bv_8_166_n228 ) : ( n968 ) ;
assign n970 =  ( n223 ) ? ( bv_8_180_n224 ) : ( n969 ) ;
assign n971 =  ( n220 ) ? ( bv_8_198_n221 ) : ( n970 ) ;
assign n972 =  ( n217 ) ? ( bv_8_232_n96 ) : ( n971 ) ;
assign n973 =  ( n214 ) ? ( bv_8_221_n136 ) : ( n972 ) ;
assign n974 =  ( n210 ) ? ( bv_8_116_n211 ) : ( n973 ) ;
assign n975 =  ( n206 ) ? ( bv_8_31_n207 ) : ( n974 ) ;
assign n976 =  ( n202 ) ? ( bv_8_75_n203 ) : ( n975 ) ;
assign n977 =  ( n198 ) ? ( bv_8_189_n199 ) : ( n976 ) ;
assign n978 =  ( n194 ) ? ( bv_8_139_n195 ) : ( n977 ) ;
assign n979 =  ( n191 ) ? ( bv_8_138_n192 ) : ( n978 ) ;
assign n980 =  ( n187 ) ? ( bv_8_112_n188 ) : ( n979 ) ;
assign n981 =  ( n183 ) ? ( bv_8_62_n184 ) : ( n980 ) ;
assign n982 =  ( n179 ) ? ( bv_8_181_n180 ) : ( n981 ) ;
assign n983 =  ( n175 ) ? ( bv_8_102_n176 ) : ( n982 ) ;
assign n984 =  ( n171 ) ? ( bv_8_72_n172 ) : ( n983 ) ;
assign n985 =  ( n167 ) ? ( bv_8_3_n168 ) : ( n984 ) ;
assign n986 =  ( n164 ) ? ( bv_8_246_n41 ) : ( n985 ) ;
assign n987 =  ( n160 ) ? ( bv_8_14_n161 ) : ( n986 ) ;
assign n988 =  ( n156 ) ? ( bv_8_97_n157 ) : ( n987 ) ;
assign n989 =  ( n152 ) ? ( bv_8_53_n153 ) : ( n988 ) ;
assign n990 =  ( n149 ) ? ( bv_8_87_n150 ) : ( n989 ) ;
assign n991 =  ( n145 ) ? ( bv_8_185_n146 ) : ( n990 ) ;
assign n992 =  ( n141 ) ? ( bv_8_134_n142 ) : ( n991 ) ;
assign n993 =  ( n137 ) ? ( bv_8_193_n138 ) : ( n992 ) ;
assign n994 =  ( n133 ) ? ( bv_8_29_n134 ) : ( n993 ) ;
assign n995 =  ( n129 ) ? ( bv_8_158_n130 ) : ( n994 ) ;
assign n996 =  ( n127 ) ? ( bv_8_225_n123 ) : ( n995 ) ;
assign n997 =  ( n124 ) ? ( bv_8_248_n33 ) : ( n996 ) ;
assign n998 =  ( n120 ) ? ( bv_8_152_n121 ) : ( n997 ) ;
assign n999 =  ( n116 ) ? ( bv_8_17_n117 ) : ( n998 ) ;
assign n1000 =  ( n112 ) ? ( bv_8_105_n113 ) : ( n999 ) ;
assign n1001 =  ( n108 ) ? ( bv_8_217_n109 ) : ( n1000 ) ;
assign n1002 =  ( n104 ) ? ( bv_8_142_n105 ) : ( n1001 ) ;
assign n1003 =  ( n101 ) ? ( bv_8_148_n102 ) : ( n1002 ) ;
assign n1004 =  ( n97 ) ? ( bv_8_155_n98 ) : ( n1003 ) ;
assign n1005 =  ( n93 ) ? ( bv_8_30_n94 ) : ( n1004 ) ;
assign n1006 =  ( n90 ) ? ( bv_8_135_n91 ) : ( n1005 ) ;
assign n1007 =  ( n86 ) ? ( bv_8_233_n87 ) : ( n1006 ) ;
assign n1008 =  ( n82 ) ? ( bv_8_206_n83 ) : ( n1007 ) ;
assign n1009 =  ( n78 ) ? ( bv_8_85_n79 ) : ( n1008 ) ;
assign n1010 =  ( n74 ) ? ( bv_8_40_n75 ) : ( n1009 ) ;
assign n1011 =  ( n70 ) ? ( bv_8_223_n71 ) : ( n1010 ) ;
assign n1012 =  ( n66 ) ? ( bv_8_140_n67 ) : ( n1011 ) ;
assign n1013 =  ( n62 ) ? ( bv_8_161_n63 ) : ( n1012 ) ;
assign n1014 =  ( n58 ) ? ( bv_8_137_n59 ) : ( n1013 ) ;
assign n1015 =  ( n54 ) ? ( bv_8_13_n55 ) : ( n1014 ) ;
assign n1016 =  ( n50 ) ? ( bv_8_191_n51 ) : ( n1015 ) ;
assign n1017 =  ( n46 ) ? ( bv_8_230_n47 ) : ( n1016 ) ;
assign n1018 =  ( n42 ) ? ( bv_8_66_n43 ) : ( n1017 ) ;
assign n1019 =  ( n38 ) ? ( bv_8_104_n39 ) : ( n1018 ) ;
assign n1020 =  ( n34 ) ? ( bv_8_65_n35 ) : ( n1019 ) ;
assign n1021 =  ( n30 ) ? ( bv_8_153_n31 ) : ( n1020 ) ;
assign n1022 =  ( n26 ) ? ( bv_8_45_n27 ) : ( n1021 ) ;
assign n1023 =  ( n22 ) ? ( bv_8_15_n23 ) : ( n1022 ) ;
assign n1024 =  ( n18 ) ? ( bv_8_176_n19 ) : ( n1023 ) ;
assign n1025 =  ( n14 ) ? ( bv_8_84_n15 ) : ( n1024 ) ;
assign n1026 =  ( n10 ) ? ( bv_8_187_n11 ) : ( n1025 ) ;
assign n1027 =  ( n6 ) ? ( bv_8_22_n7 ) : ( n1026 ) ;
assign n1028 =  ( n3 ) ^ ( n1027 )  ;
assign n1029 = in[119:112] ;
assign n1030 = in[15:8] ;
assign n1031 =  ( n1030 ) == ( bv_8_255_n5 )  ;
assign n1032 = in[15:8] ;
assign n1033 =  ( n1032 ) == ( bv_8_254_n9 )  ;
assign n1034 = in[15:8] ;
assign n1035 =  ( n1034 ) == ( bv_8_253_n13 )  ;
assign n1036 = in[15:8] ;
assign n1037 =  ( n1036 ) == ( bv_8_252_n17 )  ;
assign n1038 = in[15:8] ;
assign n1039 =  ( n1038 ) == ( bv_8_251_n21 )  ;
assign n1040 = in[15:8] ;
assign n1041 =  ( n1040 ) == ( bv_8_250_n25 )  ;
assign n1042 = in[15:8] ;
assign n1043 =  ( n1042 ) == ( bv_8_249_n29 )  ;
assign n1044 = in[15:8] ;
assign n1045 =  ( n1044 ) == ( bv_8_248_n33 )  ;
assign n1046 = in[15:8] ;
assign n1047 =  ( n1046 ) == ( bv_8_247_n37 )  ;
assign n1048 = in[15:8] ;
assign n1049 =  ( n1048 ) == ( bv_8_246_n41 )  ;
assign n1050 = in[15:8] ;
assign n1051 =  ( n1050 ) == ( bv_8_245_n45 )  ;
assign n1052 = in[15:8] ;
assign n1053 =  ( n1052 ) == ( bv_8_244_n49 )  ;
assign n1054 = in[15:8] ;
assign n1055 =  ( n1054 ) == ( bv_8_243_n53 )  ;
assign n1056 = in[15:8] ;
assign n1057 =  ( n1056 ) == ( bv_8_242_n57 )  ;
assign n1058 = in[15:8] ;
assign n1059 =  ( n1058 ) == ( bv_8_241_n61 )  ;
assign n1060 = in[15:8] ;
assign n1061 =  ( n1060 ) == ( bv_8_240_n65 )  ;
assign n1062 = in[15:8] ;
assign n1063 =  ( n1062 ) == ( bv_8_239_n69 )  ;
assign n1064 = in[15:8] ;
assign n1065 =  ( n1064 ) == ( bv_8_238_n73 )  ;
assign n1066 = in[15:8] ;
assign n1067 =  ( n1066 ) == ( bv_8_237_n77 )  ;
assign n1068 = in[15:8] ;
assign n1069 =  ( n1068 ) == ( bv_8_236_n81 )  ;
assign n1070 = in[15:8] ;
assign n1071 =  ( n1070 ) == ( bv_8_235_n85 )  ;
assign n1072 = in[15:8] ;
assign n1073 =  ( n1072 ) == ( bv_8_234_n89 )  ;
assign n1074 = in[15:8] ;
assign n1075 =  ( n1074 ) == ( bv_8_233_n87 )  ;
assign n1076 = in[15:8] ;
assign n1077 =  ( n1076 ) == ( bv_8_232_n96 )  ;
assign n1078 = in[15:8] ;
assign n1079 =  ( n1078 ) == ( bv_8_231_n100 )  ;
assign n1080 = in[15:8] ;
assign n1081 =  ( n1080 ) == ( bv_8_230_n47 )  ;
assign n1082 = in[15:8] ;
assign n1083 =  ( n1082 ) == ( bv_8_229_n107 )  ;
assign n1084 = in[15:8] ;
assign n1085 =  ( n1084 ) == ( bv_8_228_n111 )  ;
assign n1086 = in[15:8] ;
assign n1087 =  ( n1086 ) == ( bv_8_227_n115 )  ;
assign n1088 = in[15:8] ;
assign n1089 =  ( n1088 ) == ( bv_8_226_n119 )  ;
assign n1090 = in[15:8] ;
assign n1091 =  ( n1090 ) == ( bv_8_225_n123 )  ;
assign n1092 = in[15:8] ;
assign n1093 =  ( n1092 ) == ( bv_8_224_n126 )  ;
assign n1094 = in[15:8] ;
assign n1095 =  ( n1094 ) == ( bv_8_223_n71 )  ;
assign n1096 = in[15:8] ;
assign n1097 =  ( n1096 ) == ( bv_8_222_n132 )  ;
assign n1098 = in[15:8] ;
assign n1099 =  ( n1098 ) == ( bv_8_221_n136 )  ;
assign n1100 = in[15:8] ;
assign n1101 =  ( n1100 ) == ( bv_8_220_n140 )  ;
assign n1102 = in[15:8] ;
assign n1103 =  ( n1102 ) == ( bv_8_219_n144 )  ;
assign n1104 = in[15:8] ;
assign n1105 =  ( n1104 ) == ( bv_8_218_n148 )  ;
assign n1106 = in[15:8] ;
assign n1107 =  ( n1106 ) == ( bv_8_217_n109 )  ;
assign n1108 = in[15:8] ;
assign n1109 =  ( n1108 ) == ( bv_8_216_n155 )  ;
assign n1110 = in[15:8] ;
assign n1111 =  ( n1110 ) == ( bv_8_215_n159 )  ;
assign n1112 = in[15:8] ;
assign n1113 =  ( n1112 ) == ( bv_8_214_n163 )  ;
assign n1114 = in[15:8] ;
assign n1115 =  ( n1114 ) == ( bv_8_213_n166 )  ;
assign n1116 = in[15:8] ;
assign n1117 =  ( n1116 ) == ( bv_8_212_n170 )  ;
assign n1118 = in[15:8] ;
assign n1119 =  ( n1118 ) == ( bv_8_211_n174 )  ;
assign n1120 = in[15:8] ;
assign n1121 =  ( n1120 ) == ( bv_8_210_n178 )  ;
assign n1122 = in[15:8] ;
assign n1123 =  ( n1122 ) == ( bv_8_209_n182 )  ;
assign n1124 = in[15:8] ;
assign n1125 =  ( n1124 ) == ( bv_8_208_n186 )  ;
assign n1126 = in[15:8] ;
assign n1127 =  ( n1126 ) == ( bv_8_207_n190 )  ;
assign n1128 = in[15:8] ;
assign n1129 =  ( n1128 ) == ( bv_8_206_n83 )  ;
assign n1130 = in[15:8] ;
assign n1131 =  ( n1130 ) == ( bv_8_205_n197 )  ;
assign n1132 = in[15:8] ;
assign n1133 =  ( n1132 ) == ( bv_8_204_n201 )  ;
assign n1134 = in[15:8] ;
assign n1135 =  ( n1134 ) == ( bv_8_203_n205 )  ;
assign n1136 = in[15:8] ;
assign n1137 =  ( n1136 ) == ( bv_8_202_n209 )  ;
assign n1138 = in[15:8] ;
assign n1139 =  ( n1138 ) == ( bv_8_201_n213 )  ;
assign n1140 = in[15:8] ;
assign n1141 =  ( n1140 ) == ( bv_8_200_n216 )  ;
assign n1142 = in[15:8] ;
assign n1143 =  ( n1142 ) == ( bv_8_199_n219 )  ;
assign n1144 = in[15:8] ;
assign n1145 =  ( n1144 ) == ( bv_8_198_n221 )  ;
assign n1146 = in[15:8] ;
assign n1147 =  ( n1146 ) == ( bv_8_197_n226 )  ;
assign n1148 = in[15:8] ;
assign n1149 =  ( n1148 ) == ( bv_8_196_n230 )  ;
assign n1150 = in[15:8] ;
assign n1151 =  ( n1150 ) == ( bv_8_195_n234 )  ;
assign n1152 = in[15:8] ;
assign n1153 =  ( n1152 ) == ( bv_8_194_n238 )  ;
assign n1154 = in[15:8] ;
assign n1155 =  ( n1154 ) == ( bv_8_193_n138 )  ;
assign n1156 = in[15:8] ;
assign n1157 =  ( n1156 ) == ( bv_8_192_n245 )  ;
assign n1158 = in[15:8] ;
assign n1159 =  ( n1158 ) == ( bv_8_191_n51 )  ;
assign n1160 = in[15:8] ;
assign n1161 =  ( n1160 ) == ( bv_8_190_n252 )  ;
assign n1162 = in[15:8] ;
assign n1163 =  ( n1162 ) == ( bv_8_189_n199 )  ;
assign n1164 = in[15:8] ;
assign n1165 =  ( n1164 ) == ( bv_8_188_n259 )  ;
assign n1166 = in[15:8] ;
assign n1167 =  ( n1166 ) == ( bv_8_187_n11 )  ;
assign n1168 = in[15:8] ;
assign n1169 =  ( n1168 ) == ( bv_8_186_n247 )  ;
assign n1170 = in[15:8] ;
assign n1171 =  ( n1170 ) == ( bv_8_185_n146 )  ;
assign n1172 = in[15:8] ;
assign n1173 =  ( n1172 ) == ( bv_8_184_n270 )  ;
assign n1174 = in[15:8] ;
assign n1175 =  ( n1174 ) == ( bv_8_183_n274 )  ;
assign n1176 = in[15:8] ;
assign n1177 =  ( n1176 ) == ( bv_8_182_n278 )  ;
assign n1178 = in[15:8] ;
assign n1179 =  ( n1178 ) == ( bv_8_181_n180 )  ;
assign n1180 = in[15:8] ;
assign n1181 =  ( n1180 ) == ( bv_8_180_n224 )  ;
assign n1182 = in[15:8] ;
assign n1183 =  ( n1182 ) == ( bv_8_179_n287 )  ;
assign n1184 = in[15:8] ;
assign n1185 =  ( n1184 ) == ( bv_8_178_n291 )  ;
assign n1186 = in[15:8] ;
assign n1187 =  ( n1186 ) == ( bv_8_177_n295 )  ;
assign n1188 = in[15:8] ;
assign n1189 =  ( n1188 ) == ( bv_8_176_n19 )  ;
assign n1190 = in[15:8] ;
assign n1191 =  ( n1190 ) == ( bv_8_175_n300 )  ;
assign n1192 = in[15:8] ;
assign n1193 =  ( n1192 ) == ( bv_8_174_n254 )  ;
assign n1194 = in[15:8] ;
assign n1195 =  ( n1194 ) == ( bv_8_173_n306 )  ;
assign n1196 = in[15:8] ;
assign n1197 =  ( n1196 ) == ( bv_8_172_n310 )  ;
assign n1198 = in[15:8] ;
assign n1199 =  ( n1198 ) == ( bv_8_171_n314 )  ;
assign n1200 = in[15:8] ;
assign n1201 =  ( n1200 ) == ( bv_8_170_n318 )  ;
assign n1202 = in[15:8] ;
assign n1203 =  ( n1202 ) == ( bv_8_169_n276 )  ;
assign n1204 = in[15:8] ;
assign n1205 =  ( n1204 ) == ( bv_8_168_n323 )  ;
assign n1206 = in[15:8] ;
assign n1207 =  ( n1206 ) == ( bv_8_167_n326 )  ;
assign n1208 = in[15:8] ;
assign n1209 =  ( n1208 ) == ( bv_8_166_n228 )  ;
assign n1210 = in[15:8] ;
assign n1211 =  ( n1210 ) == ( bv_8_165_n333 )  ;
assign n1212 = in[15:8] ;
assign n1213 =  ( n1212 ) == ( bv_8_164_n337 )  ;
assign n1214 = in[15:8] ;
assign n1215 =  ( n1214 ) == ( bv_8_163_n341 )  ;
assign n1216 = in[15:8] ;
assign n1217 =  ( n1216 ) == ( bv_8_162_n345 )  ;
assign n1218 = in[15:8] ;
assign n1219 =  ( n1218 ) == ( bv_8_161_n63 )  ;
assign n1220 = in[15:8] ;
assign n1221 =  ( n1220 ) == ( bv_8_160_n352 )  ;
assign n1222 = in[15:8] ;
assign n1223 =  ( n1222 ) == ( bv_8_159_n355 )  ;
assign n1224 = in[15:8] ;
assign n1225 =  ( n1224 ) == ( bv_8_158_n130 )  ;
assign n1226 = in[15:8] ;
assign n1227 =  ( n1226 ) == ( bv_8_157_n361 )  ;
assign n1228 = in[15:8] ;
assign n1229 =  ( n1228 ) == ( bv_8_156_n365 )  ;
assign n1230 = in[15:8] ;
assign n1231 =  ( n1230 ) == ( bv_8_155_n98 )  ;
assign n1232 = in[15:8] ;
assign n1233 =  ( n1232 ) == ( bv_8_154_n371 )  ;
assign n1234 = in[15:8] ;
assign n1235 =  ( n1234 ) == ( bv_8_153_n31 )  ;
assign n1236 = in[15:8] ;
assign n1237 =  ( n1236 ) == ( bv_8_152_n121 )  ;
assign n1238 = in[15:8] ;
assign n1239 =  ( n1238 ) == ( bv_8_151_n379 )  ;
assign n1240 = in[15:8] ;
assign n1241 =  ( n1240 ) == ( bv_8_150_n383 )  ;
assign n1242 = in[15:8] ;
assign n1243 =  ( n1242 ) == ( bv_8_149_n308 )  ;
assign n1244 = in[15:8] ;
assign n1245 =  ( n1244 ) == ( bv_8_148_n102 )  ;
assign n1246 = in[15:8] ;
assign n1247 =  ( n1246 ) == ( bv_8_147_n393 )  ;
assign n1248 = in[15:8] ;
assign n1249 =  ( n1248 ) == ( bv_8_146_n396 )  ;
assign n1250 = in[15:8] ;
assign n1251 =  ( n1250 ) == ( bv_8_145_n312 )  ;
assign n1252 = in[15:8] ;
assign n1253 =  ( n1252 ) == ( bv_8_144_n385 )  ;
assign n1254 = in[15:8] ;
assign n1255 =  ( n1254 ) == ( bv_8_143_n406 )  ;
assign n1256 = in[15:8] ;
assign n1257 =  ( n1256 ) == ( bv_8_142_n105 )  ;
assign n1258 = in[15:8] ;
assign n1259 =  ( n1258 ) == ( bv_8_141_n285 )  ;
assign n1260 = in[15:8] ;
assign n1261 =  ( n1260 ) == ( bv_8_140_n67 )  ;
assign n1262 = in[15:8] ;
assign n1263 =  ( n1262 ) == ( bv_8_139_n195 )  ;
assign n1264 = in[15:8] ;
assign n1265 =  ( n1264 ) == ( bv_8_138_n192 )  ;
assign n1266 = in[15:8] ;
assign n1267 =  ( n1266 ) == ( bv_8_137_n59 )  ;
assign n1268 = in[15:8] ;
assign n1269 =  ( n1268 ) == ( bv_8_136_n381 )  ;
assign n1270 = in[15:8] ;
assign n1271 =  ( n1270 ) == ( bv_8_135_n91 )  ;
assign n1272 = in[15:8] ;
assign n1273 =  ( n1272 ) == ( bv_8_134_n142 )  ;
assign n1274 = in[15:8] ;
assign n1275 =  ( n1274 ) == ( bv_8_133_n435 )  ;
assign n1276 = in[15:8] ;
assign n1277 =  ( n1276 ) == ( bv_8_132_n438 )  ;
assign n1278 = in[15:8] ;
assign n1279 =  ( n1278 ) == ( bv_8_131_n442 )  ;
assign n1280 = in[15:8] ;
assign n1281 =  ( n1280 ) == ( bv_8_130_n445 )  ;
assign n1282 = in[15:8] ;
assign n1283 =  ( n1282 ) == ( bv_8_129_n401 )  ;
assign n1284 = in[15:8] ;
assign n1285 =  ( n1284 ) == ( bv_8_128_n452 )  ;
assign n1286 = in[15:8] ;
assign n1287 =  ( n1286 ) == ( bv_8_127_n455 )  ;
assign n1288 = in[15:8] ;
assign n1289 =  ( n1288 ) == ( bv_8_126_n423 )  ;
assign n1290 = in[15:8] ;
assign n1291 =  ( n1290 ) == ( bv_8_125_n460 )  ;
assign n1292 = in[15:8] ;
assign n1293 =  ( n1292 ) == ( bv_8_124_n463 )  ;
assign n1294 = in[15:8] ;
assign n1295 =  ( n1294 ) == ( bv_8_123_n467 )  ;
assign n1296 = in[15:8] ;
assign n1297 =  ( n1296 ) == ( bv_8_122_n257 )  ;
assign n1298 = in[15:8] ;
assign n1299 =  ( n1298 ) == ( bv_8_121_n302 )  ;
assign n1300 = in[15:8] ;
assign n1301 =  ( n1300 ) == ( bv_8_120_n243 )  ;
assign n1302 = in[15:8] ;
assign n1303 =  ( n1302 ) == ( bv_8_119_n477 )  ;
assign n1304 = in[15:8] ;
assign n1305 =  ( n1304 ) == ( bv_8_118_n480 )  ;
assign n1306 = in[15:8] ;
assign n1307 =  ( n1306 ) == ( bv_8_117_n484 )  ;
assign n1308 = in[15:8] ;
assign n1309 =  ( n1308 ) == ( bv_8_116_n211 )  ;
assign n1310 = in[15:8] ;
assign n1311 =  ( n1310 ) == ( bv_8_115_n408 )  ;
assign n1312 = in[15:8] ;
assign n1313 =  ( n1312 ) == ( bv_8_114_n491 )  ;
assign n1314 = in[15:8] ;
assign n1315 =  ( n1314 ) == ( bv_8_113_n495 )  ;
assign n1316 = in[15:8] ;
assign n1317 =  ( n1316 ) == ( bv_8_112_n188 )  ;
assign n1318 = in[15:8] ;
assign n1319 =  ( n1318 ) == ( bv_8_111_n501 )  ;
assign n1320 = in[15:8] ;
assign n1321 =  ( n1320 ) == ( bv_8_110_n504 )  ;
assign n1322 = in[15:8] ;
assign n1323 =  ( n1322 ) == ( bv_8_109_n289 )  ;
assign n1324 = in[15:8] ;
assign n1325 =  ( n1324 ) == ( bv_8_108_n272 )  ;
assign n1326 = in[15:8] ;
assign n1327 =  ( n1326 ) == ( bv_8_107_n513 )  ;
assign n1328 = in[15:8] ;
assign n1329 =  ( n1328 ) == ( bv_8_106_n516 )  ;
assign n1330 = in[15:8] ;
assign n1331 =  ( n1330 ) == ( bv_8_105_n113 )  ;
assign n1332 = in[15:8] ;
assign n1333 =  ( n1332 ) == ( bv_8_104_n39 )  ;
assign n1334 = in[15:8] ;
assign n1335 =  ( n1334 ) == ( bv_8_103_n525 )  ;
assign n1336 = in[15:8] ;
assign n1337 =  ( n1336 ) == ( bv_8_102_n176 )  ;
assign n1338 = in[15:8] ;
assign n1339 =  ( n1338 ) == ( bv_8_101_n261 )  ;
assign n1340 = in[15:8] ;
assign n1341 =  ( n1340 ) == ( bv_8_100_n417 )  ;
assign n1342 = in[15:8] ;
assign n1343 =  ( n1342 ) == ( bv_8_99_n537 )  ;
assign n1344 = in[15:8] ;
assign n1345 =  ( n1344 ) == ( bv_8_98_n316 )  ;
assign n1346 = in[15:8] ;
assign n1347 =  ( n1346 ) == ( bv_8_97_n157 )  ;
assign n1348 = in[15:8] ;
assign n1349 =  ( n1348 ) == ( bv_8_96_n404 )  ;
assign n1350 = in[15:8] ;
assign n1351 =  ( n1350 ) == ( bv_8_95_n440 )  ;
assign n1352 = in[15:8] ;
assign n1353 =  ( n1352 ) == ( bv_8_94_n363 )  ;
assign n1354 = in[15:8] ;
assign n1355 =  ( n1354 ) == ( bv_8_93_n414 )  ;
assign n1356 = in[15:8] ;
assign n1357 =  ( n1356 ) == ( bv_8_92_n328 )  ;
assign n1358 = in[15:8] ;
assign n1359 =  ( n1358 ) == ( bv_8_91_n557 )  ;
assign n1360 = in[15:8] ;
assign n1361 =  ( n1360 ) == ( bv_8_90_n561 )  ;
assign n1362 = in[15:8] ;
assign n1363 =  ( n1362 ) == ( bv_8_89_n564 )  ;
assign n1364 = in[15:8] ;
assign n1365 =  ( n1364 ) == ( bv_8_88_n549 )  ;
assign n1366 = in[15:8] ;
assign n1367 =  ( n1366 ) == ( bv_8_87_n150 )  ;
assign n1368 = in[15:8] ;
assign n1369 =  ( n1368 ) == ( bv_8_86_n268 )  ;
assign n1370 = in[15:8] ;
assign n1371 =  ( n1370 ) == ( bv_8_85_n79 )  ;
assign n1372 = in[15:8] ;
assign n1373 =  ( n1372 ) == ( bv_8_84_n15 )  ;
assign n1374 = in[15:8] ;
assign n1375 =  ( n1374 ) == ( bv_8_83_n578 )  ;
assign n1376 = in[15:8] ;
assign n1377 =  ( n1376 ) == ( bv_8_82_n581 )  ;
assign n1378 = in[15:8] ;
assign n1379 =  ( n1378 ) == ( bv_8_81_n499 )  ;
assign n1380 = in[15:8] ;
assign n1381 =  ( n1380 ) == ( bv_8_80_n511 )  ;
assign n1382 = in[15:8] ;
assign n1383 =  ( n1382 ) == ( bv_8_79_n398 )  ;
assign n1384 = in[15:8] ;
assign n1385 =  ( n1384 ) == ( bv_8_78_n280 )  ;
assign n1386 = in[15:8] ;
assign n1387 =  ( n1386 ) == ( bv_8_77_n532 )  ;
assign n1388 = in[15:8] ;
assign n1389 =  ( n1388 ) == ( bv_8_76_n552 )  ;
assign n1390 = in[15:8] ;
assign n1391 =  ( n1390 ) == ( bv_8_75_n203 )  ;
assign n1392 = in[15:8] ;
assign n1393 =  ( n1392 ) == ( bv_8_74_n555 )  ;
assign n1394 = in[15:8] ;
assign n1395 =  ( n1394 ) == ( bv_8_73_n339 )  ;
assign n1396 = in[15:8] ;
assign n1397 =  ( n1396 ) == ( bv_8_72_n172 )  ;
assign n1398 = in[15:8] ;
assign n1399 =  ( n1398 ) == ( bv_8_71_n608 )  ;
assign n1400 = in[15:8] ;
assign n1401 =  ( n1400 ) == ( bv_8_70_n377 )  ;
assign n1402 = in[15:8] ;
assign n1403 =  ( n1402 ) == ( bv_8_69_n523 )  ;
assign n1404 = in[15:8] ;
assign n1405 =  ( n1404 ) == ( bv_8_68_n433 )  ;
assign n1406 = in[15:8] ;
assign n1407 =  ( n1406 ) == ( bv_8_67_n535 )  ;
assign n1408 = in[15:8] ;
assign n1409 =  ( n1408 ) == ( bv_8_66_n43 )  ;
assign n1410 = in[15:8] ;
assign n1411 =  ( n1410 ) == ( bv_8_65_n35 )  ;
assign n1412 = in[15:8] ;
assign n1413 =  ( n1412 ) == ( bv_8_64_n493 )  ;
assign n1414 = in[15:8] ;
assign n1415 =  ( n1414 ) == ( bv_8_63_n629 )  ;
assign n1416 = in[15:8] ;
assign n1417 =  ( n1416 ) == ( bv_8_62_n184 )  ;
assign n1418 = in[15:8] ;
assign n1419 =  ( n1418 ) == ( bv_8_61_n420 )  ;
assign n1420 = in[15:8] ;
assign n1421 =  ( n1420 ) == ( bv_8_60_n508 )  ;
assign n1422 = in[15:8] ;
assign n1423 =  ( n1422 ) == ( bv_8_59_n604 )  ;
assign n1424 = in[15:8] ;
assign n1425 =  ( n1424 ) == ( bv_8_58_n347 )  ;
assign n1426 = in[15:8] ;
assign n1427 =  ( n1426 ) == ( bv_8_57_n559 )  ;
assign n1428 = in[15:8] ;
assign n1429 =  ( n1428 ) == ( bv_8_56_n482 )  ;
assign n1430 = in[15:8] ;
assign n1431 =  ( n1430 ) == ( bv_8_55_n293 )  ;
assign n1432 = in[15:8] ;
assign n1433 =  ( n1432 ) == ( bv_8_54_n651 )  ;
assign n1434 = in[15:8] ;
assign n1435 =  ( n1434 ) == ( bv_8_53_n153 )  ;
assign n1436 = in[15:8] ;
assign n1437 =  ( n1436 ) == ( bv_8_52_n657 )  ;
assign n1438 = in[15:8] ;
assign n1439 =  ( n1438 ) == ( bv_8_51_n529 )  ;
assign n1440 = in[15:8] ;
assign n1441 =  ( n1440 ) == ( bv_8_50_n350 )  ;
assign n1442 = in[15:8] ;
assign n1443 =  ( n1442 ) == ( bv_8_49_n666 )  ;
assign n1444 = in[15:8] ;
assign n1445 =  ( n1444 ) == ( bv_8_48_n669 )  ;
assign n1446 = in[15:8] ;
assign n1447 =  ( n1446 ) == ( bv_8_47_n592 )  ;
assign n1448 = in[15:8] ;
assign n1449 =  ( n1448 ) == ( bv_8_46_n236 )  ;
assign n1450 = in[15:8] ;
assign n1451 =  ( n1450 ) == ( bv_8_45_n27 )  ;
assign n1452 = in[15:8] ;
assign n1453 =  ( n1452 ) == ( bv_8_44_n622 )  ;
assign n1454 = in[15:8] ;
assign n1455 =  ( n1454 ) == ( bv_8_43_n682 )  ;
assign n1456 = in[15:8] ;
assign n1457 =  ( n1456 ) == ( bv_8_42_n388 )  ;
assign n1458 = in[15:8] ;
assign n1459 =  ( n1458 ) == ( bv_8_41_n597 )  ;
assign n1460 = in[15:8] ;
assign n1461 =  ( n1460 ) == ( bv_8_40_n75 )  ;
assign n1462 = in[15:8] ;
assign n1463 =  ( n1462 ) == ( bv_8_39_n635 )  ;
assign n1464 = in[15:8] ;
assign n1465 =  ( n1464 ) == ( bv_8_38_n693 )  ;
assign n1466 = in[15:8] ;
assign n1467 =  ( n1466 ) == ( bv_8_37_n240 )  ;
assign n1468 = in[15:8] ;
assign n1469 =  ( n1468 ) == ( bv_8_36_n331 )  ;
assign n1470 = in[15:8] ;
assign n1471 =  ( n1470 ) == ( bv_8_35_n664 )  ;
assign n1472 = in[15:8] ;
assign n1473 =  ( n1472 ) == ( bv_8_34_n391 )  ;
assign n1474 = in[15:8] ;
assign n1475 =  ( n1474 ) == ( bv_8_33_n469 )  ;
assign n1476 = in[15:8] ;
assign n1477 =  ( n1476 ) == ( bv_8_32_n576 )  ;
assign n1478 = in[15:8] ;
assign n1479 =  ( n1478 ) == ( bv_8_31_n207 )  ;
assign n1480 = in[15:8] ;
assign n1481 =  ( n1480 ) == ( bv_8_30_n94 )  ;
assign n1482 = in[15:8] ;
assign n1483 =  ( n1482 ) == ( bv_8_29_n134 )  ;
assign n1484 = in[15:8] ;
assign n1485 =  ( n1484 ) == ( bv_8_28_n232 )  ;
assign n1486 = in[15:8] ;
assign n1487 =  ( n1486 ) == ( bv_8_27_n616 )  ;
assign n1488 = in[15:8] ;
assign n1489 =  ( n1488 ) == ( bv_8_26_n619 )  ;
assign n1490 = in[15:8] ;
assign n1491 =  ( n1490 ) == ( bv_8_25_n411 )  ;
assign n1492 = in[15:8] ;
assign n1493 =  ( n1492 ) == ( bv_8_24_n659 )  ;
assign n1494 = in[15:8] ;
assign n1495 =  ( n1494 ) == ( bv_8_23_n430 )  ;
assign n1496 = in[15:8] ;
assign n1497 =  ( n1496 ) == ( bv_8_22_n7 )  ;
assign n1498 = in[15:8] ;
assign n1499 =  ( n1498 ) == ( bv_8_21_n674 )  ;
assign n1500 = in[15:8] ;
assign n1501 =  ( n1500 ) == ( bv_8_20_n369 )  ;
assign n1502 = in[15:8] ;
assign n1503 =  ( n1502 ) == ( bv_8_19_n447 )  ;
assign n1504 = in[15:8] ;
assign n1505 =  ( n1504 ) == ( bv_8_18_n644 )  ;
assign n1506 = in[15:8] ;
assign n1507 =  ( n1506 ) == ( bv_8_17_n117 )  ;
assign n1508 = in[15:8] ;
assign n1509 =  ( n1508 ) == ( bv_8_16_n465 )  ;
assign n1510 = in[15:8] ;
assign n1511 =  ( n1510 ) == ( bv_8_15_n23 )  ;
assign n1512 = in[15:8] ;
assign n1513 =  ( n1512 ) == ( bv_8_14_n161 )  ;
assign n1514 = in[15:8] ;
assign n1515 =  ( n1514 ) == ( bv_8_13_n55 )  ;
assign n1516 = in[15:8] ;
assign n1517 =  ( n1516 ) == ( bv_8_12_n450 )  ;
assign n1518 = in[15:8] ;
assign n1519 =  ( n1518 ) == ( bv_8_11_n359 )  ;
assign n1520 = in[15:8] ;
assign n1521 =  ( n1520 ) == ( bv_8_10_n343 )  ;
assign n1522 = in[15:8] ;
assign n1523 =  ( n1522 ) == ( bv_8_9_n627 )  ;
assign n1524 = in[15:8] ;
assign n1525 =  ( n1524 ) == ( bv_8_8_n250 )  ;
assign n1526 = in[15:8] ;
assign n1527 =  ( n1526 ) == ( bv_8_7_n647 )  ;
assign n1528 = in[15:8] ;
assign n1529 =  ( n1528 ) == ( bv_8_6_n335 )  ;
assign n1530 = in[15:8] ;
assign n1531 =  ( n1530 ) == ( bv_8_5_n653 )  ;
assign n1532 = in[15:8] ;
assign n1533 =  ( n1532 ) == ( bv_8_4_n671 )  ;
assign n1534 = in[15:8] ;
assign n1535 =  ( n1534 ) == ( bv_8_3_n168 )  ;
assign n1536 = in[15:8] ;
assign n1537 =  ( n1536 ) == ( bv_8_2_n518 )  ;
assign n1538 = in[15:8] ;
assign n1539 =  ( n1538 ) == ( bv_8_1_n753 )  ;
assign n1540 = in[15:8] ;
assign n1541 =  ( n1540 ) == ( bv_8_0_n583 )  ;
assign n1542 =  ( n1541 ) ? ( bv_8_99_n537 ) : ( bv_8_0_n583 ) ;
assign n1543 =  ( n1539 ) ? ( bv_8_124_n463 ) : ( n1542 ) ;
assign n1544 =  ( n1537 ) ? ( bv_8_119_n477 ) : ( n1543 ) ;
assign n1545 =  ( n1535 ) ? ( bv_8_123_n467 ) : ( n1544 ) ;
assign n1546 =  ( n1533 ) ? ( bv_8_242_n57 ) : ( n1545 ) ;
assign n1547 =  ( n1531 ) ? ( bv_8_107_n513 ) : ( n1546 ) ;
assign n1548 =  ( n1529 ) ? ( bv_8_111_n501 ) : ( n1547 ) ;
assign n1549 =  ( n1527 ) ? ( bv_8_197_n226 ) : ( n1548 ) ;
assign n1550 =  ( n1525 ) ? ( bv_8_48_n669 ) : ( n1549 ) ;
assign n1551 =  ( n1523 ) ? ( bv_8_1_n753 ) : ( n1550 ) ;
assign n1552 =  ( n1521 ) ? ( bv_8_103_n525 ) : ( n1551 ) ;
assign n1553 =  ( n1519 ) ? ( bv_8_43_n682 ) : ( n1552 ) ;
assign n1554 =  ( n1517 ) ? ( bv_8_254_n9 ) : ( n1553 ) ;
assign n1555 =  ( n1515 ) ? ( bv_8_215_n159 ) : ( n1554 ) ;
assign n1556 =  ( n1513 ) ? ( bv_8_171_n314 ) : ( n1555 ) ;
assign n1557 =  ( n1511 ) ? ( bv_8_118_n480 ) : ( n1556 ) ;
assign n1558 =  ( n1509 ) ? ( bv_8_202_n209 ) : ( n1557 ) ;
assign n1559 =  ( n1507 ) ? ( bv_8_130_n445 ) : ( n1558 ) ;
assign n1560 =  ( n1505 ) ? ( bv_8_201_n213 ) : ( n1559 ) ;
assign n1561 =  ( n1503 ) ? ( bv_8_125_n460 ) : ( n1560 ) ;
assign n1562 =  ( n1501 ) ? ( bv_8_250_n25 ) : ( n1561 ) ;
assign n1563 =  ( n1499 ) ? ( bv_8_89_n564 ) : ( n1562 ) ;
assign n1564 =  ( n1497 ) ? ( bv_8_71_n608 ) : ( n1563 ) ;
assign n1565 =  ( n1495 ) ? ( bv_8_240_n65 ) : ( n1564 ) ;
assign n1566 =  ( n1493 ) ? ( bv_8_173_n306 ) : ( n1565 ) ;
assign n1567 =  ( n1491 ) ? ( bv_8_212_n170 ) : ( n1566 ) ;
assign n1568 =  ( n1489 ) ? ( bv_8_162_n345 ) : ( n1567 ) ;
assign n1569 =  ( n1487 ) ? ( bv_8_175_n300 ) : ( n1568 ) ;
assign n1570 =  ( n1485 ) ? ( bv_8_156_n365 ) : ( n1569 ) ;
assign n1571 =  ( n1483 ) ? ( bv_8_164_n337 ) : ( n1570 ) ;
assign n1572 =  ( n1481 ) ? ( bv_8_114_n491 ) : ( n1571 ) ;
assign n1573 =  ( n1479 ) ? ( bv_8_192_n245 ) : ( n1572 ) ;
assign n1574 =  ( n1477 ) ? ( bv_8_183_n274 ) : ( n1573 ) ;
assign n1575 =  ( n1475 ) ? ( bv_8_253_n13 ) : ( n1574 ) ;
assign n1576 =  ( n1473 ) ? ( bv_8_147_n393 ) : ( n1575 ) ;
assign n1577 =  ( n1471 ) ? ( bv_8_38_n693 ) : ( n1576 ) ;
assign n1578 =  ( n1469 ) ? ( bv_8_54_n651 ) : ( n1577 ) ;
assign n1579 =  ( n1467 ) ? ( bv_8_63_n629 ) : ( n1578 ) ;
assign n1580 =  ( n1465 ) ? ( bv_8_247_n37 ) : ( n1579 ) ;
assign n1581 =  ( n1463 ) ? ( bv_8_204_n201 ) : ( n1580 ) ;
assign n1582 =  ( n1461 ) ? ( bv_8_52_n657 ) : ( n1581 ) ;
assign n1583 =  ( n1459 ) ? ( bv_8_165_n333 ) : ( n1582 ) ;
assign n1584 =  ( n1457 ) ? ( bv_8_229_n107 ) : ( n1583 ) ;
assign n1585 =  ( n1455 ) ? ( bv_8_241_n61 ) : ( n1584 ) ;
assign n1586 =  ( n1453 ) ? ( bv_8_113_n495 ) : ( n1585 ) ;
assign n1587 =  ( n1451 ) ? ( bv_8_216_n155 ) : ( n1586 ) ;
assign n1588 =  ( n1449 ) ? ( bv_8_49_n666 ) : ( n1587 ) ;
assign n1589 =  ( n1447 ) ? ( bv_8_21_n674 ) : ( n1588 ) ;
assign n1590 =  ( n1445 ) ? ( bv_8_4_n671 ) : ( n1589 ) ;
assign n1591 =  ( n1443 ) ? ( bv_8_199_n219 ) : ( n1590 ) ;
assign n1592 =  ( n1441 ) ? ( bv_8_35_n664 ) : ( n1591 ) ;
assign n1593 =  ( n1439 ) ? ( bv_8_195_n234 ) : ( n1592 ) ;
assign n1594 =  ( n1437 ) ? ( bv_8_24_n659 ) : ( n1593 ) ;
assign n1595 =  ( n1435 ) ? ( bv_8_150_n383 ) : ( n1594 ) ;
assign n1596 =  ( n1433 ) ? ( bv_8_5_n653 ) : ( n1595 ) ;
assign n1597 =  ( n1431 ) ? ( bv_8_154_n371 ) : ( n1596 ) ;
assign n1598 =  ( n1429 ) ? ( bv_8_7_n647 ) : ( n1597 ) ;
assign n1599 =  ( n1427 ) ? ( bv_8_18_n644 ) : ( n1598 ) ;
assign n1600 =  ( n1425 ) ? ( bv_8_128_n452 ) : ( n1599 ) ;
assign n1601 =  ( n1423 ) ? ( bv_8_226_n119 ) : ( n1600 ) ;
assign n1602 =  ( n1421 ) ? ( bv_8_235_n85 ) : ( n1601 ) ;
assign n1603 =  ( n1419 ) ? ( bv_8_39_n635 ) : ( n1602 ) ;
assign n1604 =  ( n1417 ) ? ( bv_8_178_n291 ) : ( n1603 ) ;
assign n1605 =  ( n1415 ) ? ( bv_8_117_n484 ) : ( n1604 ) ;
assign n1606 =  ( n1413 ) ? ( bv_8_9_n627 ) : ( n1605 ) ;
assign n1607 =  ( n1411 ) ? ( bv_8_131_n442 ) : ( n1606 ) ;
assign n1608 =  ( n1409 ) ? ( bv_8_44_n622 ) : ( n1607 ) ;
assign n1609 =  ( n1407 ) ? ( bv_8_26_n619 ) : ( n1608 ) ;
assign n1610 =  ( n1405 ) ? ( bv_8_27_n616 ) : ( n1609 ) ;
assign n1611 =  ( n1403 ) ? ( bv_8_110_n504 ) : ( n1610 ) ;
assign n1612 =  ( n1401 ) ? ( bv_8_90_n561 ) : ( n1611 ) ;
assign n1613 =  ( n1399 ) ? ( bv_8_160_n352 ) : ( n1612 ) ;
assign n1614 =  ( n1397 ) ? ( bv_8_82_n581 ) : ( n1613 ) ;
assign n1615 =  ( n1395 ) ? ( bv_8_59_n604 ) : ( n1614 ) ;
assign n1616 =  ( n1393 ) ? ( bv_8_214_n163 ) : ( n1615 ) ;
assign n1617 =  ( n1391 ) ? ( bv_8_179_n287 ) : ( n1616 ) ;
assign n1618 =  ( n1389 ) ? ( bv_8_41_n597 ) : ( n1617 ) ;
assign n1619 =  ( n1387 ) ? ( bv_8_227_n115 ) : ( n1618 ) ;
assign n1620 =  ( n1385 ) ? ( bv_8_47_n592 ) : ( n1619 ) ;
assign n1621 =  ( n1383 ) ? ( bv_8_132_n438 ) : ( n1620 ) ;
assign n1622 =  ( n1381 ) ? ( bv_8_83_n578 ) : ( n1621 ) ;
assign n1623 =  ( n1379 ) ? ( bv_8_209_n182 ) : ( n1622 ) ;
assign n1624 =  ( n1377 ) ? ( bv_8_0_n583 ) : ( n1623 ) ;
assign n1625 =  ( n1375 ) ? ( bv_8_237_n77 ) : ( n1624 ) ;
assign n1626 =  ( n1373 ) ? ( bv_8_32_n576 ) : ( n1625 ) ;
assign n1627 =  ( n1371 ) ? ( bv_8_252_n17 ) : ( n1626 ) ;
assign n1628 =  ( n1369 ) ? ( bv_8_177_n295 ) : ( n1627 ) ;
assign n1629 =  ( n1367 ) ? ( bv_8_91_n557 ) : ( n1628 ) ;
assign n1630 =  ( n1365 ) ? ( bv_8_106_n516 ) : ( n1629 ) ;
assign n1631 =  ( n1363 ) ? ( bv_8_203_n205 ) : ( n1630 ) ;
assign n1632 =  ( n1361 ) ? ( bv_8_190_n252 ) : ( n1631 ) ;
assign n1633 =  ( n1359 ) ? ( bv_8_57_n559 ) : ( n1632 ) ;
assign n1634 =  ( n1357 ) ? ( bv_8_74_n555 ) : ( n1633 ) ;
assign n1635 =  ( n1355 ) ? ( bv_8_76_n552 ) : ( n1634 ) ;
assign n1636 =  ( n1353 ) ? ( bv_8_88_n549 ) : ( n1635 ) ;
assign n1637 =  ( n1351 ) ? ( bv_8_207_n190 ) : ( n1636 ) ;
assign n1638 =  ( n1349 ) ? ( bv_8_208_n186 ) : ( n1637 ) ;
assign n1639 =  ( n1347 ) ? ( bv_8_239_n69 ) : ( n1638 ) ;
assign n1640 =  ( n1345 ) ? ( bv_8_170_n318 ) : ( n1639 ) ;
assign n1641 =  ( n1343 ) ? ( bv_8_251_n21 ) : ( n1640 ) ;
assign n1642 =  ( n1341 ) ? ( bv_8_67_n535 ) : ( n1641 ) ;
assign n1643 =  ( n1339 ) ? ( bv_8_77_n532 ) : ( n1642 ) ;
assign n1644 =  ( n1337 ) ? ( bv_8_51_n529 ) : ( n1643 ) ;
assign n1645 =  ( n1335 ) ? ( bv_8_133_n435 ) : ( n1644 ) ;
assign n1646 =  ( n1333 ) ? ( bv_8_69_n523 ) : ( n1645 ) ;
assign n1647 =  ( n1331 ) ? ( bv_8_249_n29 ) : ( n1646 ) ;
assign n1648 =  ( n1329 ) ? ( bv_8_2_n518 ) : ( n1647 ) ;
assign n1649 =  ( n1327 ) ? ( bv_8_127_n455 ) : ( n1648 ) ;
assign n1650 =  ( n1325 ) ? ( bv_8_80_n511 ) : ( n1649 ) ;
assign n1651 =  ( n1323 ) ? ( bv_8_60_n508 ) : ( n1650 ) ;
assign n1652 =  ( n1321 ) ? ( bv_8_159_n355 ) : ( n1651 ) ;
assign n1653 =  ( n1319 ) ? ( bv_8_168_n323 ) : ( n1652 ) ;
assign n1654 =  ( n1317 ) ? ( bv_8_81_n499 ) : ( n1653 ) ;
assign n1655 =  ( n1315 ) ? ( bv_8_163_n341 ) : ( n1654 ) ;
assign n1656 =  ( n1313 ) ? ( bv_8_64_n493 ) : ( n1655 ) ;
assign n1657 =  ( n1311 ) ? ( bv_8_143_n406 ) : ( n1656 ) ;
assign n1658 =  ( n1309 ) ? ( bv_8_146_n396 ) : ( n1657 ) ;
assign n1659 =  ( n1307 ) ? ( bv_8_157_n361 ) : ( n1658 ) ;
assign n1660 =  ( n1305 ) ? ( bv_8_56_n482 ) : ( n1659 ) ;
assign n1661 =  ( n1303 ) ? ( bv_8_245_n45 ) : ( n1660 ) ;
assign n1662 =  ( n1301 ) ? ( bv_8_188_n259 ) : ( n1661 ) ;
assign n1663 =  ( n1299 ) ? ( bv_8_182_n278 ) : ( n1662 ) ;
assign n1664 =  ( n1297 ) ? ( bv_8_218_n148 ) : ( n1663 ) ;
assign n1665 =  ( n1295 ) ? ( bv_8_33_n469 ) : ( n1664 ) ;
assign n1666 =  ( n1293 ) ? ( bv_8_16_n465 ) : ( n1665 ) ;
assign n1667 =  ( n1291 ) ? ( bv_8_255_n5 ) : ( n1666 ) ;
assign n1668 =  ( n1289 ) ? ( bv_8_243_n53 ) : ( n1667 ) ;
assign n1669 =  ( n1287 ) ? ( bv_8_210_n178 ) : ( n1668 ) ;
assign n1670 =  ( n1285 ) ? ( bv_8_205_n197 ) : ( n1669 ) ;
assign n1671 =  ( n1283 ) ? ( bv_8_12_n450 ) : ( n1670 ) ;
assign n1672 =  ( n1281 ) ? ( bv_8_19_n447 ) : ( n1671 ) ;
assign n1673 =  ( n1279 ) ? ( bv_8_236_n81 ) : ( n1672 ) ;
assign n1674 =  ( n1277 ) ? ( bv_8_95_n440 ) : ( n1673 ) ;
assign n1675 =  ( n1275 ) ? ( bv_8_151_n379 ) : ( n1674 ) ;
assign n1676 =  ( n1273 ) ? ( bv_8_68_n433 ) : ( n1675 ) ;
assign n1677 =  ( n1271 ) ? ( bv_8_23_n430 ) : ( n1676 ) ;
assign n1678 =  ( n1269 ) ? ( bv_8_196_n230 ) : ( n1677 ) ;
assign n1679 =  ( n1267 ) ? ( bv_8_167_n326 ) : ( n1678 ) ;
assign n1680 =  ( n1265 ) ? ( bv_8_126_n423 ) : ( n1679 ) ;
assign n1681 =  ( n1263 ) ? ( bv_8_61_n420 ) : ( n1680 ) ;
assign n1682 =  ( n1261 ) ? ( bv_8_100_n417 ) : ( n1681 ) ;
assign n1683 =  ( n1259 ) ? ( bv_8_93_n414 ) : ( n1682 ) ;
assign n1684 =  ( n1257 ) ? ( bv_8_25_n411 ) : ( n1683 ) ;
assign n1685 =  ( n1255 ) ? ( bv_8_115_n408 ) : ( n1684 ) ;
assign n1686 =  ( n1253 ) ? ( bv_8_96_n404 ) : ( n1685 ) ;
assign n1687 =  ( n1251 ) ? ( bv_8_129_n401 ) : ( n1686 ) ;
assign n1688 =  ( n1249 ) ? ( bv_8_79_n398 ) : ( n1687 ) ;
assign n1689 =  ( n1247 ) ? ( bv_8_220_n140 ) : ( n1688 ) ;
assign n1690 =  ( n1245 ) ? ( bv_8_34_n391 ) : ( n1689 ) ;
assign n1691 =  ( n1243 ) ? ( bv_8_42_n388 ) : ( n1690 ) ;
assign n1692 =  ( n1241 ) ? ( bv_8_144_n385 ) : ( n1691 ) ;
assign n1693 =  ( n1239 ) ? ( bv_8_136_n381 ) : ( n1692 ) ;
assign n1694 =  ( n1237 ) ? ( bv_8_70_n377 ) : ( n1693 ) ;
assign n1695 =  ( n1235 ) ? ( bv_8_238_n73 ) : ( n1694 ) ;
assign n1696 =  ( n1233 ) ? ( bv_8_184_n270 ) : ( n1695 ) ;
assign n1697 =  ( n1231 ) ? ( bv_8_20_n369 ) : ( n1696 ) ;
assign n1698 =  ( n1229 ) ? ( bv_8_222_n132 ) : ( n1697 ) ;
assign n1699 =  ( n1227 ) ? ( bv_8_94_n363 ) : ( n1698 ) ;
assign n1700 =  ( n1225 ) ? ( bv_8_11_n359 ) : ( n1699 ) ;
assign n1701 =  ( n1223 ) ? ( bv_8_219_n144 ) : ( n1700 ) ;
assign n1702 =  ( n1221 ) ? ( bv_8_224_n126 ) : ( n1701 ) ;
assign n1703 =  ( n1219 ) ? ( bv_8_50_n350 ) : ( n1702 ) ;
assign n1704 =  ( n1217 ) ? ( bv_8_58_n347 ) : ( n1703 ) ;
assign n1705 =  ( n1215 ) ? ( bv_8_10_n343 ) : ( n1704 ) ;
assign n1706 =  ( n1213 ) ? ( bv_8_73_n339 ) : ( n1705 ) ;
assign n1707 =  ( n1211 ) ? ( bv_8_6_n335 ) : ( n1706 ) ;
assign n1708 =  ( n1209 ) ? ( bv_8_36_n331 ) : ( n1707 ) ;
assign n1709 =  ( n1207 ) ? ( bv_8_92_n328 ) : ( n1708 ) ;
assign n1710 =  ( n1205 ) ? ( bv_8_194_n238 ) : ( n1709 ) ;
assign n1711 =  ( n1203 ) ? ( bv_8_211_n174 ) : ( n1710 ) ;
assign n1712 =  ( n1201 ) ? ( bv_8_172_n310 ) : ( n1711 ) ;
assign n1713 =  ( n1199 ) ? ( bv_8_98_n316 ) : ( n1712 ) ;
assign n1714 =  ( n1197 ) ? ( bv_8_145_n312 ) : ( n1713 ) ;
assign n1715 =  ( n1195 ) ? ( bv_8_149_n308 ) : ( n1714 ) ;
assign n1716 =  ( n1193 ) ? ( bv_8_228_n111 ) : ( n1715 ) ;
assign n1717 =  ( n1191 ) ? ( bv_8_121_n302 ) : ( n1716 ) ;
assign n1718 =  ( n1189 ) ? ( bv_8_231_n100 ) : ( n1717 ) ;
assign n1719 =  ( n1187 ) ? ( bv_8_200_n216 ) : ( n1718 ) ;
assign n1720 =  ( n1185 ) ? ( bv_8_55_n293 ) : ( n1719 ) ;
assign n1721 =  ( n1183 ) ? ( bv_8_109_n289 ) : ( n1720 ) ;
assign n1722 =  ( n1181 ) ? ( bv_8_141_n285 ) : ( n1721 ) ;
assign n1723 =  ( n1179 ) ? ( bv_8_213_n166 ) : ( n1722 ) ;
assign n1724 =  ( n1177 ) ? ( bv_8_78_n280 ) : ( n1723 ) ;
assign n1725 =  ( n1175 ) ? ( bv_8_169_n276 ) : ( n1724 ) ;
assign n1726 =  ( n1173 ) ? ( bv_8_108_n272 ) : ( n1725 ) ;
assign n1727 =  ( n1171 ) ? ( bv_8_86_n268 ) : ( n1726 ) ;
assign n1728 =  ( n1169 ) ? ( bv_8_244_n49 ) : ( n1727 ) ;
assign n1729 =  ( n1167 ) ? ( bv_8_234_n89 ) : ( n1728 ) ;
assign n1730 =  ( n1165 ) ? ( bv_8_101_n261 ) : ( n1729 ) ;
assign n1731 =  ( n1163 ) ? ( bv_8_122_n257 ) : ( n1730 ) ;
assign n1732 =  ( n1161 ) ? ( bv_8_174_n254 ) : ( n1731 ) ;
assign n1733 =  ( n1159 ) ? ( bv_8_8_n250 ) : ( n1732 ) ;
assign n1734 =  ( n1157 ) ? ( bv_8_186_n247 ) : ( n1733 ) ;
assign n1735 =  ( n1155 ) ? ( bv_8_120_n243 ) : ( n1734 ) ;
assign n1736 =  ( n1153 ) ? ( bv_8_37_n240 ) : ( n1735 ) ;
assign n1737 =  ( n1151 ) ? ( bv_8_46_n236 ) : ( n1736 ) ;
assign n1738 =  ( n1149 ) ? ( bv_8_28_n232 ) : ( n1737 ) ;
assign n1739 =  ( n1147 ) ? ( bv_8_166_n228 ) : ( n1738 ) ;
assign n1740 =  ( n1145 ) ? ( bv_8_180_n224 ) : ( n1739 ) ;
assign n1741 =  ( n1143 ) ? ( bv_8_198_n221 ) : ( n1740 ) ;
assign n1742 =  ( n1141 ) ? ( bv_8_232_n96 ) : ( n1741 ) ;
assign n1743 =  ( n1139 ) ? ( bv_8_221_n136 ) : ( n1742 ) ;
assign n1744 =  ( n1137 ) ? ( bv_8_116_n211 ) : ( n1743 ) ;
assign n1745 =  ( n1135 ) ? ( bv_8_31_n207 ) : ( n1744 ) ;
assign n1746 =  ( n1133 ) ? ( bv_8_75_n203 ) : ( n1745 ) ;
assign n1747 =  ( n1131 ) ? ( bv_8_189_n199 ) : ( n1746 ) ;
assign n1748 =  ( n1129 ) ? ( bv_8_139_n195 ) : ( n1747 ) ;
assign n1749 =  ( n1127 ) ? ( bv_8_138_n192 ) : ( n1748 ) ;
assign n1750 =  ( n1125 ) ? ( bv_8_112_n188 ) : ( n1749 ) ;
assign n1751 =  ( n1123 ) ? ( bv_8_62_n184 ) : ( n1750 ) ;
assign n1752 =  ( n1121 ) ? ( bv_8_181_n180 ) : ( n1751 ) ;
assign n1753 =  ( n1119 ) ? ( bv_8_102_n176 ) : ( n1752 ) ;
assign n1754 =  ( n1117 ) ? ( bv_8_72_n172 ) : ( n1753 ) ;
assign n1755 =  ( n1115 ) ? ( bv_8_3_n168 ) : ( n1754 ) ;
assign n1756 =  ( n1113 ) ? ( bv_8_246_n41 ) : ( n1755 ) ;
assign n1757 =  ( n1111 ) ? ( bv_8_14_n161 ) : ( n1756 ) ;
assign n1758 =  ( n1109 ) ? ( bv_8_97_n157 ) : ( n1757 ) ;
assign n1759 =  ( n1107 ) ? ( bv_8_53_n153 ) : ( n1758 ) ;
assign n1760 =  ( n1105 ) ? ( bv_8_87_n150 ) : ( n1759 ) ;
assign n1761 =  ( n1103 ) ? ( bv_8_185_n146 ) : ( n1760 ) ;
assign n1762 =  ( n1101 ) ? ( bv_8_134_n142 ) : ( n1761 ) ;
assign n1763 =  ( n1099 ) ? ( bv_8_193_n138 ) : ( n1762 ) ;
assign n1764 =  ( n1097 ) ? ( bv_8_29_n134 ) : ( n1763 ) ;
assign n1765 =  ( n1095 ) ? ( bv_8_158_n130 ) : ( n1764 ) ;
assign n1766 =  ( n1093 ) ? ( bv_8_225_n123 ) : ( n1765 ) ;
assign n1767 =  ( n1091 ) ? ( bv_8_248_n33 ) : ( n1766 ) ;
assign n1768 =  ( n1089 ) ? ( bv_8_152_n121 ) : ( n1767 ) ;
assign n1769 =  ( n1087 ) ? ( bv_8_17_n117 ) : ( n1768 ) ;
assign n1770 =  ( n1085 ) ? ( bv_8_105_n113 ) : ( n1769 ) ;
assign n1771 =  ( n1083 ) ? ( bv_8_217_n109 ) : ( n1770 ) ;
assign n1772 =  ( n1081 ) ? ( bv_8_142_n105 ) : ( n1771 ) ;
assign n1773 =  ( n1079 ) ? ( bv_8_148_n102 ) : ( n1772 ) ;
assign n1774 =  ( n1077 ) ? ( bv_8_155_n98 ) : ( n1773 ) ;
assign n1775 =  ( n1075 ) ? ( bv_8_30_n94 ) : ( n1774 ) ;
assign n1776 =  ( n1073 ) ? ( bv_8_135_n91 ) : ( n1775 ) ;
assign n1777 =  ( n1071 ) ? ( bv_8_233_n87 ) : ( n1776 ) ;
assign n1778 =  ( n1069 ) ? ( bv_8_206_n83 ) : ( n1777 ) ;
assign n1779 =  ( n1067 ) ? ( bv_8_85_n79 ) : ( n1778 ) ;
assign n1780 =  ( n1065 ) ? ( bv_8_40_n75 ) : ( n1779 ) ;
assign n1781 =  ( n1063 ) ? ( bv_8_223_n71 ) : ( n1780 ) ;
assign n1782 =  ( n1061 ) ? ( bv_8_140_n67 ) : ( n1781 ) ;
assign n1783 =  ( n1059 ) ? ( bv_8_161_n63 ) : ( n1782 ) ;
assign n1784 =  ( n1057 ) ? ( bv_8_137_n59 ) : ( n1783 ) ;
assign n1785 =  ( n1055 ) ? ( bv_8_13_n55 ) : ( n1784 ) ;
assign n1786 =  ( n1053 ) ? ( bv_8_191_n51 ) : ( n1785 ) ;
assign n1787 =  ( n1051 ) ? ( bv_8_230_n47 ) : ( n1786 ) ;
assign n1788 =  ( n1049 ) ? ( bv_8_66_n43 ) : ( n1787 ) ;
assign n1789 =  ( n1047 ) ? ( bv_8_104_n39 ) : ( n1788 ) ;
assign n1790 =  ( n1045 ) ? ( bv_8_65_n35 ) : ( n1789 ) ;
assign n1791 =  ( n1043 ) ? ( bv_8_153_n31 ) : ( n1790 ) ;
assign n1792 =  ( n1041 ) ? ( bv_8_45_n27 ) : ( n1791 ) ;
assign n1793 =  ( n1039 ) ? ( bv_8_15_n23 ) : ( n1792 ) ;
assign n1794 =  ( n1037 ) ? ( bv_8_176_n19 ) : ( n1793 ) ;
assign n1795 =  ( n1035 ) ? ( bv_8_84_n15 ) : ( n1794 ) ;
assign n1796 =  ( n1033 ) ? ( bv_8_187_n11 ) : ( n1795 ) ;
assign n1797 =  ( n1031 ) ? ( bv_8_22_n7 ) : ( n1796 ) ;
assign n1798 =  ( n1029 ) ^ ( n1797 )  ;
assign n1799 =  { ( n1028 ) , ( n1798 ) }  ;
assign n1800 = in[111:104] ;
assign n1801 = in[7:0] ;
assign n1802 =  ( n1801 ) == ( bv_8_255_n5 )  ;
assign n1803 = in[7:0] ;
assign n1804 =  ( n1803 ) == ( bv_8_254_n9 )  ;
assign n1805 = in[7:0] ;
assign n1806 =  ( n1805 ) == ( bv_8_253_n13 )  ;
assign n1807 = in[7:0] ;
assign n1808 =  ( n1807 ) == ( bv_8_252_n17 )  ;
assign n1809 = in[7:0] ;
assign n1810 =  ( n1809 ) == ( bv_8_251_n21 )  ;
assign n1811 = in[7:0] ;
assign n1812 =  ( n1811 ) == ( bv_8_250_n25 )  ;
assign n1813 = in[7:0] ;
assign n1814 =  ( n1813 ) == ( bv_8_249_n29 )  ;
assign n1815 = in[7:0] ;
assign n1816 =  ( n1815 ) == ( bv_8_248_n33 )  ;
assign n1817 = in[7:0] ;
assign n1818 =  ( n1817 ) == ( bv_8_247_n37 )  ;
assign n1819 = in[7:0] ;
assign n1820 =  ( n1819 ) == ( bv_8_246_n41 )  ;
assign n1821 = in[7:0] ;
assign n1822 =  ( n1821 ) == ( bv_8_245_n45 )  ;
assign n1823 = in[7:0] ;
assign n1824 =  ( n1823 ) == ( bv_8_244_n49 )  ;
assign n1825 = in[7:0] ;
assign n1826 =  ( n1825 ) == ( bv_8_243_n53 )  ;
assign n1827 = in[7:0] ;
assign n1828 =  ( n1827 ) == ( bv_8_242_n57 )  ;
assign n1829 = in[7:0] ;
assign n1830 =  ( n1829 ) == ( bv_8_241_n61 )  ;
assign n1831 = in[7:0] ;
assign n1832 =  ( n1831 ) == ( bv_8_240_n65 )  ;
assign n1833 = in[7:0] ;
assign n1834 =  ( n1833 ) == ( bv_8_239_n69 )  ;
assign n1835 = in[7:0] ;
assign n1836 =  ( n1835 ) == ( bv_8_238_n73 )  ;
assign n1837 = in[7:0] ;
assign n1838 =  ( n1837 ) == ( bv_8_237_n77 )  ;
assign n1839 = in[7:0] ;
assign n1840 =  ( n1839 ) == ( bv_8_236_n81 )  ;
assign n1841 = in[7:0] ;
assign n1842 =  ( n1841 ) == ( bv_8_235_n85 )  ;
assign n1843 = in[7:0] ;
assign n1844 =  ( n1843 ) == ( bv_8_234_n89 )  ;
assign n1845 = in[7:0] ;
assign n1846 =  ( n1845 ) == ( bv_8_233_n87 )  ;
assign n1847 = in[7:0] ;
assign n1848 =  ( n1847 ) == ( bv_8_232_n96 )  ;
assign n1849 = in[7:0] ;
assign n1850 =  ( n1849 ) == ( bv_8_231_n100 )  ;
assign n1851 = in[7:0] ;
assign n1852 =  ( n1851 ) == ( bv_8_230_n47 )  ;
assign n1853 = in[7:0] ;
assign n1854 =  ( n1853 ) == ( bv_8_229_n107 )  ;
assign n1855 = in[7:0] ;
assign n1856 =  ( n1855 ) == ( bv_8_228_n111 )  ;
assign n1857 = in[7:0] ;
assign n1858 =  ( n1857 ) == ( bv_8_227_n115 )  ;
assign n1859 = in[7:0] ;
assign n1860 =  ( n1859 ) == ( bv_8_226_n119 )  ;
assign n1861 = in[7:0] ;
assign n1862 =  ( n1861 ) == ( bv_8_225_n123 )  ;
assign n1863 = in[7:0] ;
assign n1864 =  ( n1863 ) == ( bv_8_224_n126 )  ;
assign n1865 = in[7:0] ;
assign n1866 =  ( n1865 ) == ( bv_8_223_n71 )  ;
assign n1867 = in[7:0] ;
assign n1868 =  ( n1867 ) == ( bv_8_222_n132 )  ;
assign n1869 = in[7:0] ;
assign n1870 =  ( n1869 ) == ( bv_8_221_n136 )  ;
assign n1871 = in[7:0] ;
assign n1872 =  ( n1871 ) == ( bv_8_220_n140 )  ;
assign n1873 = in[7:0] ;
assign n1874 =  ( n1873 ) == ( bv_8_219_n144 )  ;
assign n1875 = in[7:0] ;
assign n1876 =  ( n1875 ) == ( bv_8_218_n148 )  ;
assign n1877 = in[7:0] ;
assign n1878 =  ( n1877 ) == ( bv_8_217_n109 )  ;
assign n1879 = in[7:0] ;
assign n1880 =  ( n1879 ) == ( bv_8_216_n155 )  ;
assign n1881 = in[7:0] ;
assign n1882 =  ( n1881 ) == ( bv_8_215_n159 )  ;
assign n1883 = in[7:0] ;
assign n1884 =  ( n1883 ) == ( bv_8_214_n163 )  ;
assign n1885 = in[7:0] ;
assign n1886 =  ( n1885 ) == ( bv_8_213_n166 )  ;
assign n1887 = in[7:0] ;
assign n1888 =  ( n1887 ) == ( bv_8_212_n170 )  ;
assign n1889 = in[7:0] ;
assign n1890 =  ( n1889 ) == ( bv_8_211_n174 )  ;
assign n1891 = in[7:0] ;
assign n1892 =  ( n1891 ) == ( bv_8_210_n178 )  ;
assign n1893 = in[7:0] ;
assign n1894 =  ( n1893 ) == ( bv_8_209_n182 )  ;
assign n1895 = in[7:0] ;
assign n1896 =  ( n1895 ) == ( bv_8_208_n186 )  ;
assign n1897 = in[7:0] ;
assign n1898 =  ( n1897 ) == ( bv_8_207_n190 )  ;
assign n1899 = in[7:0] ;
assign n1900 =  ( n1899 ) == ( bv_8_206_n83 )  ;
assign n1901 = in[7:0] ;
assign n1902 =  ( n1901 ) == ( bv_8_205_n197 )  ;
assign n1903 = in[7:0] ;
assign n1904 =  ( n1903 ) == ( bv_8_204_n201 )  ;
assign n1905 = in[7:0] ;
assign n1906 =  ( n1905 ) == ( bv_8_203_n205 )  ;
assign n1907 = in[7:0] ;
assign n1908 =  ( n1907 ) == ( bv_8_202_n209 )  ;
assign n1909 = in[7:0] ;
assign n1910 =  ( n1909 ) == ( bv_8_201_n213 )  ;
assign n1911 = in[7:0] ;
assign n1912 =  ( n1911 ) == ( bv_8_200_n216 )  ;
assign n1913 = in[7:0] ;
assign n1914 =  ( n1913 ) == ( bv_8_199_n219 )  ;
assign n1915 = in[7:0] ;
assign n1916 =  ( n1915 ) == ( bv_8_198_n221 )  ;
assign n1917 = in[7:0] ;
assign n1918 =  ( n1917 ) == ( bv_8_197_n226 )  ;
assign n1919 = in[7:0] ;
assign n1920 =  ( n1919 ) == ( bv_8_196_n230 )  ;
assign n1921 = in[7:0] ;
assign n1922 =  ( n1921 ) == ( bv_8_195_n234 )  ;
assign n1923 = in[7:0] ;
assign n1924 =  ( n1923 ) == ( bv_8_194_n238 )  ;
assign n1925 = in[7:0] ;
assign n1926 =  ( n1925 ) == ( bv_8_193_n138 )  ;
assign n1927 = in[7:0] ;
assign n1928 =  ( n1927 ) == ( bv_8_192_n245 )  ;
assign n1929 = in[7:0] ;
assign n1930 =  ( n1929 ) == ( bv_8_191_n51 )  ;
assign n1931 = in[7:0] ;
assign n1932 =  ( n1931 ) == ( bv_8_190_n252 )  ;
assign n1933 = in[7:0] ;
assign n1934 =  ( n1933 ) == ( bv_8_189_n199 )  ;
assign n1935 = in[7:0] ;
assign n1936 =  ( n1935 ) == ( bv_8_188_n259 )  ;
assign n1937 = in[7:0] ;
assign n1938 =  ( n1937 ) == ( bv_8_187_n11 )  ;
assign n1939 = in[7:0] ;
assign n1940 =  ( n1939 ) == ( bv_8_186_n247 )  ;
assign n1941 = in[7:0] ;
assign n1942 =  ( n1941 ) == ( bv_8_185_n146 )  ;
assign n1943 = in[7:0] ;
assign n1944 =  ( n1943 ) == ( bv_8_184_n270 )  ;
assign n1945 = in[7:0] ;
assign n1946 =  ( n1945 ) == ( bv_8_183_n274 )  ;
assign n1947 = in[7:0] ;
assign n1948 =  ( n1947 ) == ( bv_8_182_n278 )  ;
assign n1949 = in[7:0] ;
assign n1950 =  ( n1949 ) == ( bv_8_181_n180 )  ;
assign n1951 = in[7:0] ;
assign n1952 =  ( n1951 ) == ( bv_8_180_n224 )  ;
assign n1953 = in[7:0] ;
assign n1954 =  ( n1953 ) == ( bv_8_179_n287 )  ;
assign n1955 = in[7:0] ;
assign n1956 =  ( n1955 ) == ( bv_8_178_n291 )  ;
assign n1957 = in[7:0] ;
assign n1958 =  ( n1957 ) == ( bv_8_177_n295 )  ;
assign n1959 = in[7:0] ;
assign n1960 =  ( n1959 ) == ( bv_8_176_n19 )  ;
assign n1961 = in[7:0] ;
assign n1962 =  ( n1961 ) == ( bv_8_175_n300 )  ;
assign n1963 = in[7:0] ;
assign n1964 =  ( n1963 ) == ( bv_8_174_n254 )  ;
assign n1965 = in[7:0] ;
assign n1966 =  ( n1965 ) == ( bv_8_173_n306 )  ;
assign n1967 = in[7:0] ;
assign n1968 =  ( n1967 ) == ( bv_8_172_n310 )  ;
assign n1969 = in[7:0] ;
assign n1970 =  ( n1969 ) == ( bv_8_171_n314 )  ;
assign n1971 = in[7:0] ;
assign n1972 =  ( n1971 ) == ( bv_8_170_n318 )  ;
assign n1973 = in[7:0] ;
assign n1974 =  ( n1973 ) == ( bv_8_169_n276 )  ;
assign n1975 = in[7:0] ;
assign n1976 =  ( n1975 ) == ( bv_8_168_n323 )  ;
assign n1977 = in[7:0] ;
assign n1978 =  ( n1977 ) == ( bv_8_167_n326 )  ;
assign n1979 = in[7:0] ;
assign n1980 =  ( n1979 ) == ( bv_8_166_n228 )  ;
assign n1981 = in[7:0] ;
assign n1982 =  ( n1981 ) == ( bv_8_165_n333 )  ;
assign n1983 = in[7:0] ;
assign n1984 =  ( n1983 ) == ( bv_8_164_n337 )  ;
assign n1985 = in[7:0] ;
assign n1986 =  ( n1985 ) == ( bv_8_163_n341 )  ;
assign n1987 = in[7:0] ;
assign n1988 =  ( n1987 ) == ( bv_8_162_n345 )  ;
assign n1989 = in[7:0] ;
assign n1990 =  ( n1989 ) == ( bv_8_161_n63 )  ;
assign n1991 = in[7:0] ;
assign n1992 =  ( n1991 ) == ( bv_8_160_n352 )  ;
assign n1993 = in[7:0] ;
assign n1994 =  ( n1993 ) == ( bv_8_159_n355 )  ;
assign n1995 = in[7:0] ;
assign n1996 =  ( n1995 ) == ( bv_8_158_n130 )  ;
assign n1997 = in[7:0] ;
assign n1998 =  ( n1997 ) == ( bv_8_157_n361 )  ;
assign n1999 = in[7:0] ;
assign n2000 =  ( n1999 ) == ( bv_8_156_n365 )  ;
assign n2001 = in[7:0] ;
assign n2002 =  ( n2001 ) == ( bv_8_155_n98 )  ;
assign n2003 = in[7:0] ;
assign n2004 =  ( n2003 ) == ( bv_8_154_n371 )  ;
assign n2005 = in[7:0] ;
assign n2006 =  ( n2005 ) == ( bv_8_153_n31 )  ;
assign n2007 = in[7:0] ;
assign n2008 =  ( n2007 ) == ( bv_8_152_n121 )  ;
assign n2009 = in[7:0] ;
assign n2010 =  ( n2009 ) == ( bv_8_151_n379 )  ;
assign n2011 = in[7:0] ;
assign n2012 =  ( n2011 ) == ( bv_8_150_n383 )  ;
assign n2013 = in[7:0] ;
assign n2014 =  ( n2013 ) == ( bv_8_149_n308 )  ;
assign n2015 = in[7:0] ;
assign n2016 =  ( n2015 ) == ( bv_8_148_n102 )  ;
assign n2017 = in[7:0] ;
assign n2018 =  ( n2017 ) == ( bv_8_147_n393 )  ;
assign n2019 = in[7:0] ;
assign n2020 =  ( n2019 ) == ( bv_8_146_n396 )  ;
assign n2021 = in[7:0] ;
assign n2022 =  ( n2021 ) == ( bv_8_145_n312 )  ;
assign n2023 = in[7:0] ;
assign n2024 =  ( n2023 ) == ( bv_8_144_n385 )  ;
assign n2025 = in[7:0] ;
assign n2026 =  ( n2025 ) == ( bv_8_143_n406 )  ;
assign n2027 = in[7:0] ;
assign n2028 =  ( n2027 ) == ( bv_8_142_n105 )  ;
assign n2029 = in[7:0] ;
assign n2030 =  ( n2029 ) == ( bv_8_141_n285 )  ;
assign n2031 = in[7:0] ;
assign n2032 =  ( n2031 ) == ( bv_8_140_n67 )  ;
assign n2033 = in[7:0] ;
assign n2034 =  ( n2033 ) == ( bv_8_139_n195 )  ;
assign n2035 = in[7:0] ;
assign n2036 =  ( n2035 ) == ( bv_8_138_n192 )  ;
assign n2037 = in[7:0] ;
assign n2038 =  ( n2037 ) == ( bv_8_137_n59 )  ;
assign n2039 = in[7:0] ;
assign n2040 =  ( n2039 ) == ( bv_8_136_n381 )  ;
assign n2041 = in[7:0] ;
assign n2042 =  ( n2041 ) == ( bv_8_135_n91 )  ;
assign n2043 = in[7:0] ;
assign n2044 =  ( n2043 ) == ( bv_8_134_n142 )  ;
assign n2045 = in[7:0] ;
assign n2046 =  ( n2045 ) == ( bv_8_133_n435 )  ;
assign n2047 = in[7:0] ;
assign n2048 =  ( n2047 ) == ( bv_8_132_n438 )  ;
assign n2049 = in[7:0] ;
assign n2050 =  ( n2049 ) == ( bv_8_131_n442 )  ;
assign n2051 = in[7:0] ;
assign n2052 =  ( n2051 ) == ( bv_8_130_n445 )  ;
assign n2053 = in[7:0] ;
assign n2054 =  ( n2053 ) == ( bv_8_129_n401 )  ;
assign n2055 = in[7:0] ;
assign n2056 =  ( n2055 ) == ( bv_8_128_n452 )  ;
assign n2057 = in[7:0] ;
assign n2058 =  ( n2057 ) == ( bv_8_127_n455 )  ;
assign n2059 = in[7:0] ;
assign n2060 =  ( n2059 ) == ( bv_8_126_n423 )  ;
assign n2061 = in[7:0] ;
assign n2062 =  ( n2061 ) == ( bv_8_125_n460 )  ;
assign n2063 = in[7:0] ;
assign n2064 =  ( n2063 ) == ( bv_8_124_n463 )  ;
assign n2065 = in[7:0] ;
assign n2066 =  ( n2065 ) == ( bv_8_123_n467 )  ;
assign n2067 = in[7:0] ;
assign n2068 =  ( n2067 ) == ( bv_8_122_n257 )  ;
assign n2069 = in[7:0] ;
assign n2070 =  ( n2069 ) == ( bv_8_121_n302 )  ;
assign n2071 = in[7:0] ;
assign n2072 =  ( n2071 ) == ( bv_8_120_n243 )  ;
assign n2073 = in[7:0] ;
assign n2074 =  ( n2073 ) == ( bv_8_119_n477 )  ;
assign n2075 = in[7:0] ;
assign n2076 =  ( n2075 ) == ( bv_8_118_n480 )  ;
assign n2077 = in[7:0] ;
assign n2078 =  ( n2077 ) == ( bv_8_117_n484 )  ;
assign n2079 = in[7:0] ;
assign n2080 =  ( n2079 ) == ( bv_8_116_n211 )  ;
assign n2081 = in[7:0] ;
assign n2082 =  ( n2081 ) == ( bv_8_115_n408 )  ;
assign n2083 = in[7:0] ;
assign n2084 =  ( n2083 ) == ( bv_8_114_n491 )  ;
assign n2085 = in[7:0] ;
assign n2086 =  ( n2085 ) == ( bv_8_113_n495 )  ;
assign n2087 = in[7:0] ;
assign n2088 =  ( n2087 ) == ( bv_8_112_n188 )  ;
assign n2089 = in[7:0] ;
assign n2090 =  ( n2089 ) == ( bv_8_111_n501 )  ;
assign n2091 = in[7:0] ;
assign n2092 =  ( n2091 ) == ( bv_8_110_n504 )  ;
assign n2093 = in[7:0] ;
assign n2094 =  ( n2093 ) == ( bv_8_109_n289 )  ;
assign n2095 = in[7:0] ;
assign n2096 =  ( n2095 ) == ( bv_8_108_n272 )  ;
assign n2097 = in[7:0] ;
assign n2098 =  ( n2097 ) == ( bv_8_107_n513 )  ;
assign n2099 = in[7:0] ;
assign n2100 =  ( n2099 ) == ( bv_8_106_n516 )  ;
assign n2101 = in[7:0] ;
assign n2102 =  ( n2101 ) == ( bv_8_105_n113 )  ;
assign n2103 = in[7:0] ;
assign n2104 =  ( n2103 ) == ( bv_8_104_n39 )  ;
assign n2105 = in[7:0] ;
assign n2106 =  ( n2105 ) == ( bv_8_103_n525 )  ;
assign n2107 = in[7:0] ;
assign n2108 =  ( n2107 ) == ( bv_8_102_n176 )  ;
assign n2109 = in[7:0] ;
assign n2110 =  ( n2109 ) == ( bv_8_101_n261 )  ;
assign n2111 = in[7:0] ;
assign n2112 =  ( n2111 ) == ( bv_8_100_n417 )  ;
assign n2113 = in[7:0] ;
assign n2114 =  ( n2113 ) == ( bv_8_99_n537 )  ;
assign n2115 = in[7:0] ;
assign n2116 =  ( n2115 ) == ( bv_8_98_n316 )  ;
assign n2117 = in[7:0] ;
assign n2118 =  ( n2117 ) == ( bv_8_97_n157 )  ;
assign n2119 = in[7:0] ;
assign n2120 =  ( n2119 ) == ( bv_8_96_n404 )  ;
assign n2121 = in[7:0] ;
assign n2122 =  ( n2121 ) == ( bv_8_95_n440 )  ;
assign n2123 = in[7:0] ;
assign n2124 =  ( n2123 ) == ( bv_8_94_n363 )  ;
assign n2125 = in[7:0] ;
assign n2126 =  ( n2125 ) == ( bv_8_93_n414 )  ;
assign n2127 = in[7:0] ;
assign n2128 =  ( n2127 ) == ( bv_8_92_n328 )  ;
assign n2129 = in[7:0] ;
assign n2130 =  ( n2129 ) == ( bv_8_91_n557 )  ;
assign n2131 = in[7:0] ;
assign n2132 =  ( n2131 ) == ( bv_8_90_n561 )  ;
assign n2133 = in[7:0] ;
assign n2134 =  ( n2133 ) == ( bv_8_89_n564 )  ;
assign n2135 = in[7:0] ;
assign n2136 =  ( n2135 ) == ( bv_8_88_n549 )  ;
assign n2137 = in[7:0] ;
assign n2138 =  ( n2137 ) == ( bv_8_87_n150 )  ;
assign n2139 = in[7:0] ;
assign n2140 =  ( n2139 ) == ( bv_8_86_n268 )  ;
assign n2141 = in[7:0] ;
assign n2142 =  ( n2141 ) == ( bv_8_85_n79 )  ;
assign n2143 = in[7:0] ;
assign n2144 =  ( n2143 ) == ( bv_8_84_n15 )  ;
assign n2145 = in[7:0] ;
assign n2146 =  ( n2145 ) == ( bv_8_83_n578 )  ;
assign n2147 = in[7:0] ;
assign n2148 =  ( n2147 ) == ( bv_8_82_n581 )  ;
assign n2149 = in[7:0] ;
assign n2150 =  ( n2149 ) == ( bv_8_81_n499 )  ;
assign n2151 = in[7:0] ;
assign n2152 =  ( n2151 ) == ( bv_8_80_n511 )  ;
assign n2153 = in[7:0] ;
assign n2154 =  ( n2153 ) == ( bv_8_79_n398 )  ;
assign n2155 = in[7:0] ;
assign n2156 =  ( n2155 ) == ( bv_8_78_n280 )  ;
assign n2157 = in[7:0] ;
assign n2158 =  ( n2157 ) == ( bv_8_77_n532 )  ;
assign n2159 = in[7:0] ;
assign n2160 =  ( n2159 ) == ( bv_8_76_n552 )  ;
assign n2161 = in[7:0] ;
assign n2162 =  ( n2161 ) == ( bv_8_75_n203 )  ;
assign n2163 = in[7:0] ;
assign n2164 =  ( n2163 ) == ( bv_8_74_n555 )  ;
assign n2165 = in[7:0] ;
assign n2166 =  ( n2165 ) == ( bv_8_73_n339 )  ;
assign n2167 = in[7:0] ;
assign n2168 =  ( n2167 ) == ( bv_8_72_n172 )  ;
assign n2169 = in[7:0] ;
assign n2170 =  ( n2169 ) == ( bv_8_71_n608 )  ;
assign n2171 = in[7:0] ;
assign n2172 =  ( n2171 ) == ( bv_8_70_n377 )  ;
assign n2173 = in[7:0] ;
assign n2174 =  ( n2173 ) == ( bv_8_69_n523 )  ;
assign n2175 = in[7:0] ;
assign n2176 =  ( n2175 ) == ( bv_8_68_n433 )  ;
assign n2177 = in[7:0] ;
assign n2178 =  ( n2177 ) == ( bv_8_67_n535 )  ;
assign n2179 = in[7:0] ;
assign n2180 =  ( n2179 ) == ( bv_8_66_n43 )  ;
assign n2181 = in[7:0] ;
assign n2182 =  ( n2181 ) == ( bv_8_65_n35 )  ;
assign n2183 = in[7:0] ;
assign n2184 =  ( n2183 ) == ( bv_8_64_n493 )  ;
assign n2185 = in[7:0] ;
assign n2186 =  ( n2185 ) == ( bv_8_63_n629 )  ;
assign n2187 = in[7:0] ;
assign n2188 =  ( n2187 ) == ( bv_8_62_n184 )  ;
assign n2189 = in[7:0] ;
assign n2190 =  ( n2189 ) == ( bv_8_61_n420 )  ;
assign n2191 = in[7:0] ;
assign n2192 =  ( n2191 ) == ( bv_8_60_n508 )  ;
assign n2193 = in[7:0] ;
assign n2194 =  ( n2193 ) == ( bv_8_59_n604 )  ;
assign n2195 = in[7:0] ;
assign n2196 =  ( n2195 ) == ( bv_8_58_n347 )  ;
assign n2197 = in[7:0] ;
assign n2198 =  ( n2197 ) == ( bv_8_57_n559 )  ;
assign n2199 = in[7:0] ;
assign n2200 =  ( n2199 ) == ( bv_8_56_n482 )  ;
assign n2201 = in[7:0] ;
assign n2202 =  ( n2201 ) == ( bv_8_55_n293 )  ;
assign n2203 = in[7:0] ;
assign n2204 =  ( n2203 ) == ( bv_8_54_n651 )  ;
assign n2205 = in[7:0] ;
assign n2206 =  ( n2205 ) == ( bv_8_53_n153 )  ;
assign n2207 = in[7:0] ;
assign n2208 =  ( n2207 ) == ( bv_8_52_n657 )  ;
assign n2209 = in[7:0] ;
assign n2210 =  ( n2209 ) == ( bv_8_51_n529 )  ;
assign n2211 = in[7:0] ;
assign n2212 =  ( n2211 ) == ( bv_8_50_n350 )  ;
assign n2213 = in[7:0] ;
assign n2214 =  ( n2213 ) == ( bv_8_49_n666 )  ;
assign n2215 = in[7:0] ;
assign n2216 =  ( n2215 ) == ( bv_8_48_n669 )  ;
assign n2217 = in[7:0] ;
assign n2218 =  ( n2217 ) == ( bv_8_47_n592 )  ;
assign n2219 = in[7:0] ;
assign n2220 =  ( n2219 ) == ( bv_8_46_n236 )  ;
assign n2221 = in[7:0] ;
assign n2222 =  ( n2221 ) == ( bv_8_45_n27 )  ;
assign n2223 = in[7:0] ;
assign n2224 =  ( n2223 ) == ( bv_8_44_n622 )  ;
assign n2225 = in[7:0] ;
assign n2226 =  ( n2225 ) == ( bv_8_43_n682 )  ;
assign n2227 = in[7:0] ;
assign n2228 =  ( n2227 ) == ( bv_8_42_n388 )  ;
assign n2229 = in[7:0] ;
assign n2230 =  ( n2229 ) == ( bv_8_41_n597 )  ;
assign n2231 = in[7:0] ;
assign n2232 =  ( n2231 ) == ( bv_8_40_n75 )  ;
assign n2233 = in[7:0] ;
assign n2234 =  ( n2233 ) == ( bv_8_39_n635 )  ;
assign n2235 = in[7:0] ;
assign n2236 =  ( n2235 ) == ( bv_8_38_n693 )  ;
assign n2237 = in[7:0] ;
assign n2238 =  ( n2237 ) == ( bv_8_37_n240 )  ;
assign n2239 = in[7:0] ;
assign n2240 =  ( n2239 ) == ( bv_8_36_n331 )  ;
assign n2241 = in[7:0] ;
assign n2242 =  ( n2241 ) == ( bv_8_35_n664 )  ;
assign n2243 = in[7:0] ;
assign n2244 =  ( n2243 ) == ( bv_8_34_n391 )  ;
assign n2245 = in[7:0] ;
assign n2246 =  ( n2245 ) == ( bv_8_33_n469 )  ;
assign n2247 = in[7:0] ;
assign n2248 =  ( n2247 ) == ( bv_8_32_n576 )  ;
assign n2249 = in[7:0] ;
assign n2250 =  ( n2249 ) == ( bv_8_31_n207 )  ;
assign n2251 = in[7:0] ;
assign n2252 =  ( n2251 ) == ( bv_8_30_n94 )  ;
assign n2253 = in[7:0] ;
assign n2254 =  ( n2253 ) == ( bv_8_29_n134 )  ;
assign n2255 = in[7:0] ;
assign n2256 =  ( n2255 ) == ( bv_8_28_n232 )  ;
assign n2257 = in[7:0] ;
assign n2258 =  ( n2257 ) == ( bv_8_27_n616 )  ;
assign n2259 = in[7:0] ;
assign n2260 =  ( n2259 ) == ( bv_8_26_n619 )  ;
assign n2261 = in[7:0] ;
assign n2262 =  ( n2261 ) == ( bv_8_25_n411 )  ;
assign n2263 = in[7:0] ;
assign n2264 =  ( n2263 ) == ( bv_8_24_n659 )  ;
assign n2265 = in[7:0] ;
assign n2266 =  ( n2265 ) == ( bv_8_23_n430 )  ;
assign n2267 = in[7:0] ;
assign n2268 =  ( n2267 ) == ( bv_8_22_n7 )  ;
assign n2269 = in[7:0] ;
assign n2270 =  ( n2269 ) == ( bv_8_21_n674 )  ;
assign n2271 = in[7:0] ;
assign n2272 =  ( n2271 ) == ( bv_8_20_n369 )  ;
assign n2273 = in[7:0] ;
assign n2274 =  ( n2273 ) == ( bv_8_19_n447 )  ;
assign n2275 = in[7:0] ;
assign n2276 =  ( n2275 ) == ( bv_8_18_n644 )  ;
assign n2277 = in[7:0] ;
assign n2278 =  ( n2277 ) == ( bv_8_17_n117 )  ;
assign n2279 = in[7:0] ;
assign n2280 =  ( n2279 ) == ( bv_8_16_n465 )  ;
assign n2281 = in[7:0] ;
assign n2282 =  ( n2281 ) == ( bv_8_15_n23 )  ;
assign n2283 = in[7:0] ;
assign n2284 =  ( n2283 ) == ( bv_8_14_n161 )  ;
assign n2285 = in[7:0] ;
assign n2286 =  ( n2285 ) == ( bv_8_13_n55 )  ;
assign n2287 = in[7:0] ;
assign n2288 =  ( n2287 ) == ( bv_8_12_n450 )  ;
assign n2289 = in[7:0] ;
assign n2290 =  ( n2289 ) == ( bv_8_11_n359 )  ;
assign n2291 = in[7:0] ;
assign n2292 =  ( n2291 ) == ( bv_8_10_n343 )  ;
assign n2293 = in[7:0] ;
assign n2294 =  ( n2293 ) == ( bv_8_9_n627 )  ;
assign n2295 = in[7:0] ;
assign n2296 =  ( n2295 ) == ( bv_8_8_n250 )  ;
assign n2297 = in[7:0] ;
assign n2298 =  ( n2297 ) == ( bv_8_7_n647 )  ;
assign n2299 = in[7:0] ;
assign n2300 =  ( n2299 ) == ( bv_8_6_n335 )  ;
assign n2301 = in[7:0] ;
assign n2302 =  ( n2301 ) == ( bv_8_5_n653 )  ;
assign n2303 = in[7:0] ;
assign n2304 =  ( n2303 ) == ( bv_8_4_n671 )  ;
assign n2305 = in[7:0] ;
assign n2306 =  ( n2305 ) == ( bv_8_3_n168 )  ;
assign n2307 = in[7:0] ;
assign n2308 =  ( n2307 ) == ( bv_8_2_n518 )  ;
assign n2309 = in[7:0] ;
assign n2310 =  ( n2309 ) == ( bv_8_1_n753 )  ;
assign n2311 = in[7:0] ;
assign n2312 =  ( n2311 ) == ( bv_8_0_n583 )  ;
assign n2313 =  ( n2312 ) ? ( bv_8_99_n537 ) : ( bv_8_0_n583 ) ;
assign n2314 =  ( n2310 ) ? ( bv_8_124_n463 ) : ( n2313 ) ;
assign n2315 =  ( n2308 ) ? ( bv_8_119_n477 ) : ( n2314 ) ;
assign n2316 =  ( n2306 ) ? ( bv_8_123_n467 ) : ( n2315 ) ;
assign n2317 =  ( n2304 ) ? ( bv_8_242_n57 ) : ( n2316 ) ;
assign n2318 =  ( n2302 ) ? ( bv_8_107_n513 ) : ( n2317 ) ;
assign n2319 =  ( n2300 ) ? ( bv_8_111_n501 ) : ( n2318 ) ;
assign n2320 =  ( n2298 ) ? ( bv_8_197_n226 ) : ( n2319 ) ;
assign n2321 =  ( n2296 ) ? ( bv_8_48_n669 ) : ( n2320 ) ;
assign n2322 =  ( n2294 ) ? ( bv_8_1_n753 ) : ( n2321 ) ;
assign n2323 =  ( n2292 ) ? ( bv_8_103_n525 ) : ( n2322 ) ;
assign n2324 =  ( n2290 ) ? ( bv_8_43_n682 ) : ( n2323 ) ;
assign n2325 =  ( n2288 ) ? ( bv_8_254_n9 ) : ( n2324 ) ;
assign n2326 =  ( n2286 ) ? ( bv_8_215_n159 ) : ( n2325 ) ;
assign n2327 =  ( n2284 ) ? ( bv_8_171_n314 ) : ( n2326 ) ;
assign n2328 =  ( n2282 ) ? ( bv_8_118_n480 ) : ( n2327 ) ;
assign n2329 =  ( n2280 ) ? ( bv_8_202_n209 ) : ( n2328 ) ;
assign n2330 =  ( n2278 ) ? ( bv_8_130_n445 ) : ( n2329 ) ;
assign n2331 =  ( n2276 ) ? ( bv_8_201_n213 ) : ( n2330 ) ;
assign n2332 =  ( n2274 ) ? ( bv_8_125_n460 ) : ( n2331 ) ;
assign n2333 =  ( n2272 ) ? ( bv_8_250_n25 ) : ( n2332 ) ;
assign n2334 =  ( n2270 ) ? ( bv_8_89_n564 ) : ( n2333 ) ;
assign n2335 =  ( n2268 ) ? ( bv_8_71_n608 ) : ( n2334 ) ;
assign n2336 =  ( n2266 ) ? ( bv_8_240_n65 ) : ( n2335 ) ;
assign n2337 =  ( n2264 ) ? ( bv_8_173_n306 ) : ( n2336 ) ;
assign n2338 =  ( n2262 ) ? ( bv_8_212_n170 ) : ( n2337 ) ;
assign n2339 =  ( n2260 ) ? ( bv_8_162_n345 ) : ( n2338 ) ;
assign n2340 =  ( n2258 ) ? ( bv_8_175_n300 ) : ( n2339 ) ;
assign n2341 =  ( n2256 ) ? ( bv_8_156_n365 ) : ( n2340 ) ;
assign n2342 =  ( n2254 ) ? ( bv_8_164_n337 ) : ( n2341 ) ;
assign n2343 =  ( n2252 ) ? ( bv_8_114_n491 ) : ( n2342 ) ;
assign n2344 =  ( n2250 ) ? ( bv_8_192_n245 ) : ( n2343 ) ;
assign n2345 =  ( n2248 ) ? ( bv_8_183_n274 ) : ( n2344 ) ;
assign n2346 =  ( n2246 ) ? ( bv_8_253_n13 ) : ( n2345 ) ;
assign n2347 =  ( n2244 ) ? ( bv_8_147_n393 ) : ( n2346 ) ;
assign n2348 =  ( n2242 ) ? ( bv_8_38_n693 ) : ( n2347 ) ;
assign n2349 =  ( n2240 ) ? ( bv_8_54_n651 ) : ( n2348 ) ;
assign n2350 =  ( n2238 ) ? ( bv_8_63_n629 ) : ( n2349 ) ;
assign n2351 =  ( n2236 ) ? ( bv_8_247_n37 ) : ( n2350 ) ;
assign n2352 =  ( n2234 ) ? ( bv_8_204_n201 ) : ( n2351 ) ;
assign n2353 =  ( n2232 ) ? ( bv_8_52_n657 ) : ( n2352 ) ;
assign n2354 =  ( n2230 ) ? ( bv_8_165_n333 ) : ( n2353 ) ;
assign n2355 =  ( n2228 ) ? ( bv_8_229_n107 ) : ( n2354 ) ;
assign n2356 =  ( n2226 ) ? ( bv_8_241_n61 ) : ( n2355 ) ;
assign n2357 =  ( n2224 ) ? ( bv_8_113_n495 ) : ( n2356 ) ;
assign n2358 =  ( n2222 ) ? ( bv_8_216_n155 ) : ( n2357 ) ;
assign n2359 =  ( n2220 ) ? ( bv_8_49_n666 ) : ( n2358 ) ;
assign n2360 =  ( n2218 ) ? ( bv_8_21_n674 ) : ( n2359 ) ;
assign n2361 =  ( n2216 ) ? ( bv_8_4_n671 ) : ( n2360 ) ;
assign n2362 =  ( n2214 ) ? ( bv_8_199_n219 ) : ( n2361 ) ;
assign n2363 =  ( n2212 ) ? ( bv_8_35_n664 ) : ( n2362 ) ;
assign n2364 =  ( n2210 ) ? ( bv_8_195_n234 ) : ( n2363 ) ;
assign n2365 =  ( n2208 ) ? ( bv_8_24_n659 ) : ( n2364 ) ;
assign n2366 =  ( n2206 ) ? ( bv_8_150_n383 ) : ( n2365 ) ;
assign n2367 =  ( n2204 ) ? ( bv_8_5_n653 ) : ( n2366 ) ;
assign n2368 =  ( n2202 ) ? ( bv_8_154_n371 ) : ( n2367 ) ;
assign n2369 =  ( n2200 ) ? ( bv_8_7_n647 ) : ( n2368 ) ;
assign n2370 =  ( n2198 ) ? ( bv_8_18_n644 ) : ( n2369 ) ;
assign n2371 =  ( n2196 ) ? ( bv_8_128_n452 ) : ( n2370 ) ;
assign n2372 =  ( n2194 ) ? ( bv_8_226_n119 ) : ( n2371 ) ;
assign n2373 =  ( n2192 ) ? ( bv_8_235_n85 ) : ( n2372 ) ;
assign n2374 =  ( n2190 ) ? ( bv_8_39_n635 ) : ( n2373 ) ;
assign n2375 =  ( n2188 ) ? ( bv_8_178_n291 ) : ( n2374 ) ;
assign n2376 =  ( n2186 ) ? ( bv_8_117_n484 ) : ( n2375 ) ;
assign n2377 =  ( n2184 ) ? ( bv_8_9_n627 ) : ( n2376 ) ;
assign n2378 =  ( n2182 ) ? ( bv_8_131_n442 ) : ( n2377 ) ;
assign n2379 =  ( n2180 ) ? ( bv_8_44_n622 ) : ( n2378 ) ;
assign n2380 =  ( n2178 ) ? ( bv_8_26_n619 ) : ( n2379 ) ;
assign n2381 =  ( n2176 ) ? ( bv_8_27_n616 ) : ( n2380 ) ;
assign n2382 =  ( n2174 ) ? ( bv_8_110_n504 ) : ( n2381 ) ;
assign n2383 =  ( n2172 ) ? ( bv_8_90_n561 ) : ( n2382 ) ;
assign n2384 =  ( n2170 ) ? ( bv_8_160_n352 ) : ( n2383 ) ;
assign n2385 =  ( n2168 ) ? ( bv_8_82_n581 ) : ( n2384 ) ;
assign n2386 =  ( n2166 ) ? ( bv_8_59_n604 ) : ( n2385 ) ;
assign n2387 =  ( n2164 ) ? ( bv_8_214_n163 ) : ( n2386 ) ;
assign n2388 =  ( n2162 ) ? ( bv_8_179_n287 ) : ( n2387 ) ;
assign n2389 =  ( n2160 ) ? ( bv_8_41_n597 ) : ( n2388 ) ;
assign n2390 =  ( n2158 ) ? ( bv_8_227_n115 ) : ( n2389 ) ;
assign n2391 =  ( n2156 ) ? ( bv_8_47_n592 ) : ( n2390 ) ;
assign n2392 =  ( n2154 ) ? ( bv_8_132_n438 ) : ( n2391 ) ;
assign n2393 =  ( n2152 ) ? ( bv_8_83_n578 ) : ( n2392 ) ;
assign n2394 =  ( n2150 ) ? ( bv_8_209_n182 ) : ( n2393 ) ;
assign n2395 =  ( n2148 ) ? ( bv_8_0_n583 ) : ( n2394 ) ;
assign n2396 =  ( n2146 ) ? ( bv_8_237_n77 ) : ( n2395 ) ;
assign n2397 =  ( n2144 ) ? ( bv_8_32_n576 ) : ( n2396 ) ;
assign n2398 =  ( n2142 ) ? ( bv_8_252_n17 ) : ( n2397 ) ;
assign n2399 =  ( n2140 ) ? ( bv_8_177_n295 ) : ( n2398 ) ;
assign n2400 =  ( n2138 ) ? ( bv_8_91_n557 ) : ( n2399 ) ;
assign n2401 =  ( n2136 ) ? ( bv_8_106_n516 ) : ( n2400 ) ;
assign n2402 =  ( n2134 ) ? ( bv_8_203_n205 ) : ( n2401 ) ;
assign n2403 =  ( n2132 ) ? ( bv_8_190_n252 ) : ( n2402 ) ;
assign n2404 =  ( n2130 ) ? ( bv_8_57_n559 ) : ( n2403 ) ;
assign n2405 =  ( n2128 ) ? ( bv_8_74_n555 ) : ( n2404 ) ;
assign n2406 =  ( n2126 ) ? ( bv_8_76_n552 ) : ( n2405 ) ;
assign n2407 =  ( n2124 ) ? ( bv_8_88_n549 ) : ( n2406 ) ;
assign n2408 =  ( n2122 ) ? ( bv_8_207_n190 ) : ( n2407 ) ;
assign n2409 =  ( n2120 ) ? ( bv_8_208_n186 ) : ( n2408 ) ;
assign n2410 =  ( n2118 ) ? ( bv_8_239_n69 ) : ( n2409 ) ;
assign n2411 =  ( n2116 ) ? ( bv_8_170_n318 ) : ( n2410 ) ;
assign n2412 =  ( n2114 ) ? ( bv_8_251_n21 ) : ( n2411 ) ;
assign n2413 =  ( n2112 ) ? ( bv_8_67_n535 ) : ( n2412 ) ;
assign n2414 =  ( n2110 ) ? ( bv_8_77_n532 ) : ( n2413 ) ;
assign n2415 =  ( n2108 ) ? ( bv_8_51_n529 ) : ( n2414 ) ;
assign n2416 =  ( n2106 ) ? ( bv_8_133_n435 ) : ( n2415 ) ;
assign n2417 =  ( n2104 ) ? ( bv_8_69_n523 ) : ( n2416 ) ;
assign n2418 =  ( n2102 ) ? ( bv_8_249_n29 ) : ( n2417 ) ;
assign n2419 =  ( n2100 ) ? ( bv_8_2_n518 ) : ( n2418 ) ;
assign n2420 =  ( n2098 ) ? ( bv_8_127_n455 ) : ( n2419 ) ;
assign n2421 =  ( n2096 ) ? ( bv_8_80_n511 ) : ( n2420 ) ;
assign n2422 =  ( n2094 ) ? ( bv_8_60_n508 ) : ( n2421 ) ;
assign n2423 =  ( n2092 ) ? ( bv_8_159_n355 ) : ( n2422 ) ;
assign n2424 =  ( n2090 ) ? ( bv_8_168_n323 ) : ( n2423 ) ;
assign n2425 =  ( n2088 ) ? ( bv_8_81_n499 ) : ( n2424 ) ;
assign n2426 =  ( n2086 ) ? ( bv_8_163_n341 ) : ( n2425 ) ;
assign n2427 =  ( n2084 ) ? ( bv_8_64_n493 ) : ( n2426 ) ;
assign n2428 =  ( n2082 ) ? ( bv_8_143_n406 ) : ( n2427 ) ;
assign n2429 =  ( n2080 ) ? ( bv_8_146_n396 ) : ( n2428 ) ;
assign n2430 =  ( n2078 ) ? ( bv_8_157_n361 ) : ( n2429 ) ;
assign n2431 =  ( n2076 ) ? ( bv_8_56_n482 ) : ( n2430 ) ;
assign n2432 =  ( n2074 ) ? ( bv_8_245_n45 ) : ( n2431 ) ;
assign n2433 =  ( n2072 ) ? ( bv_8_188_n259 ) : ( n2432 ) ;
assign n2434 =  ( n2070 ) ? ( bv_8_182_n278 ) : ( n2433 ) ;
assign n2435 =  ( n2068 ) ? ( bv_8_218_n148 ) : ( n2434 ) ;
assign n2436 =  ( n2066 ) ? ( bv_8_33_n469 ) : ( n2435 ) ;
assign n2437 =  ( n2064 ) ? ( bv_8_16_n465 ) : ( n2436 ) ;
assign n2438 =  ( n2062 ) ? ( bv_8_255_n5 ) : ( n2437 ) ;
assign n2439 =  ( n2060 ) ? ( bv_8_243_n53 ) : ( n2438 ) ;
assign n2440 =  ( n2058 ) ? ( bv_8_210_n178 ) : ( n2439 ) ;
assign n2441 =  ( n2056 ) ? ( bv_8_205_n197 ) : ( n2440 ) ;
assign n2442 =  ( n2054 ) ? ( bv_8_12_n450 ) : ( n2441 ) ;
assign n2443 =  ( n2052 ) ? ( bv_8_19_n447 ) : ( n2442 ) ;
assign n2444 =  ( n2050 ) ? ( bv_8_236_n81 ) : ( n2443 ) ;
assign n2445 =  ( n2048 ) ? ( bv_8_95_n440 ) : ( n2444 ) ;
assign n2446 =  ( n2046 ) ? ( bv_8_151_n379 ) : ( n2445 ) ;
assign n2447 =  ( n2044 ) ? ( bv_8_68_n433 ) : ( n2446 ) ;
assign n2448 =  ( n2042 ) ? ( bv_8_23_n430 ) : ( n2447 ) ;
assign n2449 =  ( n2040 ) ? ( bv_8_196_n230 ) : ( n2448 ) ;
assign n2450 =  ( n2038 ) ? ( bv_8_167_n326 ) : ( n2449 ) ;
assign n2451 =  ( n2036 ) ? ( bv_8_126_n423 ) : ( n2450 ) ;
assign n2452 =  ( n2034 ) ? ( bv_8_61_n420 ) : ( n2451 ) ;
assign n2453 =  ( n2032 ) ? ( bv_8_100_n417 ) : ( n2452 ) ;
assign n2454 =  ( n2030 ) ? ( bv_8_93_n414 ) : ( n2453 ) ;
assign n2455 =  ( n2028 ) ? ( bv_8_25_n411 ) : ( n2454 ) ;
assign n2456 =  ( n2026 ) ? ( bv_8_115_n408 ) : ( n2455 ) ;
assign n2457 =  ( n2024 ) ? ( bv_8_96_n404 ) : ( n2456 ) ;
assign n2458 =  ( n2022 ) ? ( bv_8_129_n401 ) : ( n2457 ) ;
assign n2459 =  ( n2020 ) ? ( bv_8_79_n398 ) : ( n2458 ) ;
assign n2460 =  ( n2018 ) ? ( bv_8_220_n140 ) : ( n2459 ) ;
assign n2461 =  ( n2016 ) ? ( bv_8_34_n391 ) : ( n2460 ) ;
assign n2462 =  ( n2014 ) ? ( bv_8_42_n388 ) : ( n2461 ) ;
assign n2463 =  ( n2012 ) ? ( bv_8_144_n385 ) : ( n2462 ) ;
assign n2464 =  ( n2010 ) ? ( bv_8_136_n381 ) : ( n2463 ) ;
assign n2465 =  ( n2008 ) ? ( bv_8_70_n377 ) : ( n2464 ) ;
assign n2466 =  ( n2006 ) ? ( bv_8_238_n73 ) : ( n2465 ) ;
assign n2467 =  ( n2004 ) ? ( bv_8_184_n270 ) : ( n2466 ) ;
assign n2468 =  ( n2002 ) ? ( bv_8_20_n369 ) : ( n2467 ) ;
assign n2469 =  ( n2000 ) ? ( bv_8_222_n132 ) : ( n2468 ) ;
assign n2470 =  ( n1998 ) ? ( bv_8_94_n363 ) : ( n2469 ) ;
assign n2471 =  ( n1996 ) ? ( bv_8_11_n359 ) : ( n2470 ) ;
assign n2472 =  ( n1994 ) ? ( bv_8_219_n144 ) : ( n2471 ) ;
assign n2473 =  ( n1992 ) ? ( bv_8_224_n126 ) : ( n2472 ) ;
assign n2474 =  ( n1990 ) ? ( bv_8_50_n350 ) : ( n2473 ) ;
assign n2475 =  ( n1988 ) ? ( bv_8_58_n347 ) : ( n2474 ) ;
assign n2476 =  ( n1986 ) ? ( bv_8_10_n343 ) : ( n2475 ) ;
assign n2477 =  ( n1984 ) ? ( bv_8_73_n339 ) : ( n2476 ) ;
assign n2478 =  ( n1982 ) ? ( bv_8_6_n335 ) : ( n2477 ) ;
assign n2479 =  ( n1980 ) ? ( bv_8_36_n331 ) : ( n2478 ) ;
assign n2480 =  ( n1978 ) ? ( bv_8_92_n328 ) : ( n2479 ) ;
assign n2481 =  ( n1976 ) ? ( bv_8_194_n238 ) : ( n2480 ) ;
assign n2482 =  ( n1974 ) ? ( bv_8_211_n174 ) : ( n2481 ) ;
assign n2483 =  ( n1972 ) ? ( bv_8_172_n310 ) : ( n2482 ) ;
assign n2484 =  ( n1970 ) ? ( bv_8_98_n316 ) : ( n2483 ) ;
assign n2485 =  ( n1968 ) ? ( bv_8_145_n312 ) : ( n2484 ) ;
assign n2486 =  ( n1966 ) ? ( bv_8_149_n308 ) : ( n2485 ) ;
assign n2487 =  ( n1964 ) ? ( bv_8_228_n111 ) : ( n2486 ) ;
assign n2488 =  ( n1962 ) ? ( bv_8_121_n302 ) : ( n2487 ) ;
assign n2489 =  ( n1960 ) ? ( bv_8_231_n100 ) : ( n2488 ) ;
assign n2490 =  ( n1958 ) ? ( bv_8_200_n216 ) : ( n2489 ) ;
assign n2491 =  ( n1956 ) ? ( bv_8_55_n293 ) : ( n2490 ) ;
assign n2492 =  ( n1954 ) ? ( bv_8_109_n289 ) : ( n2491 ) ;
assign n2493 =  ( n1952 ) ? ( bv_8_141_n285 ) : ( n2492 ) ;
assign n2494 =  ( n1950 ) ? ( bv_8_213_n166 ) : ( n2493 ) ;
assign n2495 =  ( n1948 ) ? ( bv_8_78_n280 ) : ( n2494 ) ;
assign n2496 =  ( n1946 ) ? ( bv_8_169_n276 ) : ( n2495 ) ;
assign n2497 =  ( n1944 ) ? ( bv_8_108_n272 ) : ( n2496 ) ;
assign n2498 =  ( n1942 ) ? ( bv_8_86_n268 ) : ( n2497 ) ;
assign n2499 =  ( n1940 ) ? ( bv_8_244_n49 ) : ( n2498 ) ;
assign n2500 =  ( n1938 ) ? ( bv_8_234_n89 ) : ( n2499 ) ;
assign n2501 =  ( n1936 ) ? ( bv_8_101_n261 ) : ( n2500 ) ;
assign n2502 =  ( n1934 ) ? ( bv_8_122_n257 ) : ( n2501 ) ;
assign n2503 =  ( n1932 ) ? ( bv_8_174_n254 ) : ( n2502 ) ;
assign n2504 =  ( n1930 ) ? ( bv_8_8_n250 ) : ( n2503 ) ;
assign n2505 =  ( n1928 ) ? ( bv_8_186_n247 ) : ( n2504 ) ;
assign n2506 =  ( n1926 ) ? ( bv_8_120_n243 ) : ( n2505 ) ;
assign n2507 =  ( n1924 ) ? ( bv_8_37_n240 ) : ( n2506 ) ;
assign n2508 =  ( n1922 ) ? ( bv_8_46_n236 ) : ( n2507 ) ;
assign n2509 =  ( n1920 ) ? ( bv_8_28_n232 ) : ( n2508 ) ;
assign n2510 =  ( n1918 ) ? ( bv_8_166_n228 ) : ( n2509 ) ;
assign n2511 =  ( n1916 ) ? ( bv_8_180_n224 ) : ( n2510 ) ;
assign n2512 =  ( n1914 ) ? ( bv_8_198_n221 ) : ( n2511 ) ;
assign n2513 =  ( n1912 ) ? ( bv_8_232_n96 ) : ( n2512 ) ;
assign n2514 =  ( n1910 ) ? ( bv_8_221_n136 ) : ( n2513 ) ;
assign n2515 =  ( n1908 ) ? ( bv_8_116_n211 ) : ( n2514 ) ;
assign n2516 =  ( n1906 ) ? ( bv_8_31_n207 ) : ( n2515 ) ;
assign n2517 =  ( n1904 ) ? ( bv_8_75_n203 ) : ( n2516 ) ;
assign n2518 =  ( n1902 ) ? ( bv_8_189_n199 ) : ( n2517 ) ;
assign n2519 =  ( n1900 ) ? ( bv_8_139_n195 ) : ( n2518 ) ;
assign n2520 =  ( n1898 ) ? ( bv_8_138_n192 ) : ( n2519 ) ;
assign n2521 =  ( n1896 ) ? ( bv_8_112_n188 ) : ( n2520 ) ;
assign n2522 =  ( n1894 ) ? ( bv_8_62_n184 ) : ( n2521 ) ;
assign n2523 =  ( n1892 ) ? ( bv_8_181_n180 ) : ( n2522 ) ;
assign n2524 =  ( n1890 ) ? ( bv_8_102_n176 ) : ( n2523 ) ;
assign n2525 =  ( n1888 ) ? ( bv_8_72_n172 ) : ( n2524 ) ;
assign n2526 =  ( n1886 ) ? ( bv_8_3_n168 ) : ( n2525 ) ;
assign n2527 =  ( n1884 ) ? ( bv_8_246_n41 ) : ( n2526 ) ;
assign n2528 =  ( n1882 ) ? ( bv_8_14_n161 ) : ( n2527 ) ;
assign n2529 =  ( n1880 ) ? ( bv_8_97_n157 ) : ( n2528 ) ;
assign n2530 =  ( n1878 ) ? ( bv_8_53_n153 ) : ( n2529 ) ;
assign n2531 =  ( n1876 ) ? ( bv_8_87_n150 ) : ( n2530 ) ;
assign n2532 =  ( n1874 ) ? ( bv_8_185_n146 ) : ( n2531 ) ;
assign n2533 =  ( n1872 ) ? ( bv_8_134_n142 ) : ( n2532 ) ;
assign n2534 =  ( n1870 ) ? ( bv_8_193_n138 ) : ( n2533 ) ;
assign n2535 =  ( n1868 ) ? ( bv_8_29_n134 ) : ( n2534 ) ;
assign n2536 =  ( n1866 ) ? ( bv_8_158_n130 ) : ( n2535 ) ;
assign n2537 =  ( n1864 ) ? ( bv_8_225_n123 ) : ( n2536 ) ;
assign n2538 =  ( n1862 ) ? ( bv_8_248_n33 ) : ( n2537 ) ;
assign n2539 =  ( n1860 ) ? ( bv_8_152_n121 ) : ( n2538 ) ;
assign n2540 =  ( n1858 ) ? ( bv_8_17_n117 ) : ( n2539 ) ;
assign n2541 =  ( n1856 ) ? ( bv_8_105_n113 ) : ( n2540 ) ;
assign n2542 =  ( n1854 ) ? ( bv_8_217_n109 ) : ( n2541 ) ;
assign n2543 =  ( n1852 ) ? ( bv_8_142_n105 ) : ( n2542 ) ;
assign n2544 =  ( n1850 ) ? ( bv_8_148_n102 ) : ( n2543 ) ;
assign n2545 =  ( n1848 ) ? ( bv_8_155_n98 ) : ( n2544 ) ;
assign n2546 =  ( n1846 ) ? ( bv_8_30_n94 ) : ( n2545 ) ;
assign n2547 =  ( n1844 ) ? ( bv_8_135_n91 ) : ( n2546 ) ;
assign n2548 =  ( n1842 ) ? ( bv_8_233_n87 ) : ( n2547 ) ;
assign n2549 =  ( n1840 ) ? ( bv_8_206_n83 ) : ( n2548 ) ;
assign n2550 =  ( n1838 ) ? ( bv_8_85_n79 ) : ( n2549 ) ;
assign n2551 =  ( n1836 ) ? ( bv_8_40_n75 ) : ( n2550 ) ;
assign n2552 =  ( n1834 ) ? ( bv_8_223_n71 ) : ( n2551 ) ;
assign n2553 =  ( n1832 ) ? ( bv_8_140_n67 ) : ( n2552 ) ;
assign n2554 =  ( n1830 ) ? ( bv_8_161_n63 ) : ( n2553 ) ;
assign n2555 =  ( n1828 ) ? ( bv_8_137_n59 ) : ( n2554 ) ;
assign n2556 =  ( n1826 ) ? ( bv_8_13_n55 ) : ( n2555 ) ;
assign n2557 =  ( n1824 ) ? ( bv_8_191_n51 ) : ( n2556 ) ;
assign n2558 =  ( n1822 ) ? ( bv_8_230_n47 ) : ( n2557 ) ;
assign n2559 =  ( n1820 ) ? ( bv_8_66_n43 ) : ( n2558 ) ;
assign n2560 =  ( n1818 ) ? ( bv_8_104_n39 ) : ( n2559 ) ;
assign n2561 =  ( n1816 ) ? ( bv_8_65_n35 ) : ( n2560 ) ;
assign n2562 =  ( n1814 ) ? ( bv_8_153_n31 ) : ( n2561 ) ;
assign n2563 =  ( n1812 ) ? ( bv_8_45_n27 ) : ( n2562 ) ;
assign n2564 =  ( n1810 ) ? ( bv_8_15_n23 ) : ( n2563 ) ;
assign n2565 =  ( n1808 ) ? ( bv_8_176_n19 ) : ( n2564 ) ;
assign n2566 =  ( n1806 ) ? ( bv_8_84_n15 ) : ( n2565 ) ;
assign n2567 =  ( n1804 ) ? ( bv_8_187_n11 ) : ( n2566 ) ;
assign n2568 =  ( n1802 ) ? ( bv_8_22_n7 ) : ( n2567 ) ;
assign n2569 =  ( n1800 ) ^ ( n2568 )  ;
assign n2570 =  { ( n1799 ) , ( n2569 ) }  ;
assign n2571 = in[103:96] ;
assign n2572 = in[31:24] ;
assign n2573 =  ( n2572 ) == ( bv_8_255_n5 )  ;
assign n2574 = in[31:24] ;
assign n2575 =  ( n2574 ) == ( bv_8_254_n9 )  ;
assign n2576 = in[31:24] ;
assign n2577 =  ( n2576 ) == ( bv_8_253_n13 )  ;
assign n2578 = in[31:24] ;
assign n2579 =  ( n2578 ) == ( bv_8_252_n17 )  ;
assign n2580 = in[31:24] ;
assign n2581 =  ( n2580 ) == ( bv_8_251_n21 )  ;
assign n2582 = in[31:24] ;
assign n2583 =  ( n2582 ) == ( bv_8_250_n25 )  ;
assign n2584 = in[31:24] ;
assign n2585 =  ( n2584 ) == ( bv_8_249_n29 )  ;
assign n2586 = in[31:24] ;
assign n2587 =  ( n2586 ) == ( bv_8_248_n33 )  ;
assign n2588 = in[31:24] ;
assign n2589 =  ( n2588 ) == ( bv_8_247_n37 )  ;
assign n2590 = in[31:24] ;
assign n2591 =  ( n2590 ) == ( bv_8_246_n41 )  ;
assign n2592 = in[31:24] ;
assign n2593 =  ( n2592 ) == ( bv_8_245_n45 )  ;
assign n2594 = in[31:24] ;
assign n2595 =  ( n2594 ) == ( bv_8_244_n49 )  ;
assign n2596 = in[31:24] ;
assign n2597 =  ( n2596 ) == ( bv_8_243_n53 )  ;
assign n2598 = in[31:24] ;
assign n2599 =  ( n2598 ) == ( bv_8_242_n57 )  ;
assign n2600 = in[31:24] ;
assign n2601 =  ( n2600 ) == ( bv_8_241_n61 )  ;
assign n2602 = in[31:24] ;
assign n2603 =  ( n2602 ) == ( bv_8_240_n65 )  ;
assign n2604 = in[31:24] ;
assign n2605 =  ( n2604 ) == ( bv_8_239_n69 )  ;
assign n2606 = in[31:24] ;
assign n2607 =  ( n2606 ) == ( bv_8_238_n73 )  ;
assign n2608 = in[31:24] ;
assign n2609 =  ( n2608 ) == ( bv_8_237_n77 )  ;
assign n2610 = in[31:24] ;
assign n2611 =  ( n2610 ) == ( bv_8_236_n81 )  ;
assign n2612 = in[31:24] ;
assign n2613 =  ( n2612 ) == ( bv_8_235_n85 )  ;
assign n2614 = in[31:24] ;
assign n2615 =  ( n2614 ) == ( bv_8_234_n89 )  ;
assign n2616 = in[31:24] ;
assign n2617 =  ( n2616 ) == ( bv_8_233_n87 )  ;
assign n2618 = in[31:24] ;
assign n2619 =  ( n2618 ) == ( bv_8_232_n96 )  ;
assign n2620 = in[31:24] ;
assign n2621 =  ( n2620 ) == ( bv_8_231_n100 )  ;
assign n2622 = in[31:24] ;
assign n2623 =  ( n2622 ) == ( bv_8_230_n47 )  ;
assign n2624 = in[31:24] ;
assign n2625 =  ( n2624 ) == ( bv_8_229_n107 )  ;
assign n2626 = in[31:24] ;
assign n2627 =  ( n2626 ) == ( bv_8_228_n111 )  ;
assign n2628 = in[31:24] ;
assign n2629 =  ( n2628 ) == ( bv_8_227_n115 )  ;
assign n2630 = in[31:24] ;
assign n2631 =  ( n2630 ) == ( bv_8_226_n119 )  ;
assign n2632 = in[31:24] ;
assign n2633 =  ( n2632 ) == ( bv_8_225_n123 )  ;
assign n2634 = in[31:24] ;
assign n2635 =  ( n2634 ) == ( bv_8_224_n126 )  ;
assign n2636 = in[31:24] ;
assign n2637 =  ( n2636 ) == ( bv_8_223_n71 )  ;
assign n2638 = in[31:24] ;
assign n2639 =  ( n2638 ) == ( bv_8_222_n132 )  ;
assign n2640 = in[31:24] ;
assign n2641 =  ( n2640 ) == ( bv_8_221_n136 )  ;
assign n2642 = in[31:24] ;
assign n2643 =  ( n2642 ) == ( bv_8_220_n140 )  ;
assign n2644 = in[31:24] ;
assign n2645 =  ( n2644 ) == ( bv_8_219_n144 )  ;
assign n2646 = in[31:24] ;
assign n2647 =  ( n2646 ) == ( bv_8_218_n148 )  ;
assign n2648 = in[31:24] ;
assign n2649 =  ( n2648 ) == ( bv_8_217_n109 )  ;
assign n2650 = in[31:24] ;
assign n2651 =  ( n2650 ) == ( bv_8_216_n155 )  ;
assign n2652 = in[31:24] ;
assign n2653 =  ( n2652 ) == ( bv_8_215_n159 )  ;
assign n2654 = in[31:24] ;
assign n2655 =  ( n2654 ) == ( bv_8_214_n163 )  ;
assign n2656 = in[31:24] ;
assign n2657 =  ( n2656 ) == ( bv_8_213_n166 )  ;
assign n2658 = in[31:24] ;
assign n2659 =  ( n2658 ) == ( bv_8_212_n170 )  ;
assign n2660 = in[31:24] ;
assign n2661 =  ( n2660 ) == ( bv_8_211_n174 )  ;
assign n2662 = in[31:24] ;
assign n2663 =  ( n2662 ) == ( bv_8_210_n178 )  ;
assign n2664 = in[31:24] ;
assign n2665 =  ( n2664 ) == ( bv_8_209_n182 )  ;
assign n2666 = in[31:24] ;
assign n2667 =  ( n2666 ) == ( bv_8_208_n186 )  ;
assign n2668 = in[31:24] ;
assign n2669 =  ( n2668 ) == ( bv_8_207_n190 )  ;
assign n2670 = in[31:24] ;
assign n2671 =  ( n2670 ) == ( bv_8_206_n83 )  ;
assign n2672 = in[31:24] ;
assign n2673 =  ( n2672 ) == ( bv_8_205_n197 )  ;
assign n2674 = in[31:24] ;
assign n2675 =  ( n2674 ) == ( bv_8_204_n201 )  ;
assign n2676 = in[31:24] ;
assign n2677 =  ( n2676 ) == ( bv_8_203_n205 )  ;
assign n2678 = in[31:24] ;
assign n2679 =  ( n2678 ) == ( bv_8_202_n209 )  ;
assign n2680 = in[31:24] ;
assign n2681 =  ( n2680 ) == ( bv_8_201_n213 )  ;
assign n2682 = in[31:24] ;
assign n2683 =  ( n2682 ) == ( bv_8_200_n216 )  ;
assign n2684 = in[31:24] ;
assign n2685 =  ( n2684 ) == ( bv_8_199_n219 )  ;
assign n2686 = in[31:24] ;
assign n2687 =  ( n2686 ) == ( bv_8_198_n221 )  ;
assign n2688 = in[31:24] ;
assign n2689 =  ( n2688 ) == ( bv_8_197_n226 )  ;
assign n2690 = in[31:24] ;
assign n2691 =  ( n2690 ) == ( bv_8_196_n230 )  ;
assign n2692 = in[31:24] ;
assign n2693 =  ( n2692 ) == ( bv_8_195_n234 )  ;
assign n2694 = in[31:24] ;
assign n2695 =  ( n2694 ) == ( bv_8_194_n238 )  ;
assign n2696 = in[31:24] ;
assign n2697 =  ( n2696 ) == ( bv_8_193_n138 )  ;
assign n2698 = in[31:24] ;
assign n2699 =  ( n2698 ) == ( bv_8_192_n245 )  ;
assign n2700 = in[31:24] ;
assign n2701 =  ( n2700 ) == ( bv_8_191_n51 )  ;
assign n2702 = in[31:24] ;
assign n2703 =  ( n2702 ) == ( bv_8_190_n252 )  ;
assign n2704 = in[31:24] ;
assign n2705 =  ( n2704 ) == ( bv_8_189_n199 )  ;
assign n2706 = in[31:24] ;
assign n2707 =  ( n2706 ) == ( bv_8_188_n259 )  ;
assign n2708 = in[31:24] ;
assign n2709 =  ( n2708 ) == ( bv_8_187_n11 )  ;
assign n2710 = in[31:24] ;
assign n2711 =  ( n2710 ) == ( bv_8_186_n247 )  ;
assign n2712 = in[31:24] ;
assign n2713 =  ( n2712 ) == ( bv_8_185_n146 )  ;
assign n2714 = in[31:24] ;
assign n2715 =  ( n2714 ) == ( bv_8_184_n270 )  ;
assign n2716 = in[31:24] ;
assign n2717 =  ( n2716 ) == ( bv_8_183_n274 )  ;
assign n2718 = in[31:24] ;
assign n2719 =  ( n2718 ) == ( bv_8_182_n278 )  ;
assign n2720 = in[31:24] ;
assign n2721 =  ( n2720 ) == ( bv_8_181_n180 )  ;
assign n2722 = in[31:24] ;
assign n2723 =  ( n2722 ) == ( bv_8_180_n224 )  ;
assign n2724 = in[31:24] ;
assign n2725 =  ( n2724 ) == ( bv_8_179_n287 )  ;
assign n2726 = in[31:24] ;
assign n2727 =  ( n2726 ) == ( bv_8_178_n291 )  ;
assign n2728 = in[31:24] ;
assign n2729 =  ( n2728 ) == ( bv_8_177_n295 )  ;
assign n2730 = in[31:24] ;
assign n2731 =  ( n2730 ) == ( bv_8_176_n19 )  ;
assign n2732 = in[31:24] ;
assign n2733 =  ( n2732 ) == ( bv_8_175_n300 )  ;
assign n2734 = in[31:24] ;
assign n2735 =  ( n2734 ) == ( bv_8_174_n254 )  ;
assign n2736 = in[31:24] ;
assign n2737 =  ( n2736 ) == ( bv_8_173_n306 )  ;
assign n2738 = in[31:24] ;
assign n2739 =  ( n2738 ) == ( bv_8_172_n310 )  ;
assign n2740 = in[31:24] ;
assign n2741 =  ( n2740 ) == ( bv_8_171_n314 )  ;
assign n2742 = in[31:24] ;
assign n2743 =  ( n2742 ) == ( bv_8_170_n318 )  ;
assign n2744 = in[31:24] ;
assign n2745 =  ( n2744 ) == ( bv_8_169_n276 )  ;
assign n2746 = in[31:24] ;
assign n2747 =  ( n2746 ) == ( bv_8_168_n323 )  ;
assign n2748 = in[31:24] ;
assign n2749 =  ( n2748 ) == ( bv_8_167_n326 )  ;
assign n2750 = in[31:24] ;
assign n2751 =  ( n2750 ) == ( bv_8_166_n228 )  ;
assign n2752 = in[31:24] ;
assign n2753 =  ( n2752 ) == ( bv_8_165_n333 )  ;
assign n2754 = in[31:24] ;
assign n2755 =  ( n2754 ) == ( bv_8_164_n337 )  ;
assign n2756 = in[31:24] ;
assign n2757 =  ( n2756 ) == ( bv_8_163_n341 )  ;
assign n2758 = in[31:24] ;
assign n2759 =  ( n2758 ) == ( bv_8_162_n345 )  ;
assign n2760 = in[31:24] ;
assign n2761 =  ( n2760 ) == ( bv_8_161_n63 )  ;
assign n2762 = in[31:24] ;
assign n2763 =  ( n2762 ) == ( bv_8_160_n352 )  ;
assign n2764 = in[31:24] ;
assign n2765 =  ( n2764 ) == ( bv_8_159_n355 )  ;
assign n2766 = in[31:24] ;
assign n2767 =  ( n2766 ) == ( bv_8_158_n130 )  ;
assign n2768 = in[31:24] ;
assign n2769 =  ( n2768 ) == ( bv_8_157_n361 )  ;
assign n2770 = in[31:24] ;
assign n2771 =  ( n2770 ) == ( bv_8_156_n365 )  ;
assign n2772 = in[31:24] ;
assign n2773 =  ( n2772 ) == ( bv_8_155_n98 )  ;
assign n2774 = in[31:24] ;
assign n2775 =  ( n2774 ) == ( bv_8_154_n371 )  ;
assign n2776 = in[31:24] ;
assign n2777 =  ( n2776 ) == ( bv_8_153_n31 )  ;
assign n2778 = in[31:24] ;
assign n2779 =  ( n2778 ) == ( bv_8_152_n121 )  ;
assign n2780 = in[31:24] ;
assign n2781 =  ( n2780 ) == ( bv_8_151_n379 )  ;
assign n2782 = in[31:24] ;
assign n2783 =  ( n2782 ) == ( bv_8_150_n383 )  ;
assign n2784 = in[31:24] ;
assign n2785 =  ( n2784 ) == ( bv_8_149_n308 )  ;
assign n2786 = in[31:24] ;
assign n2787 =  ( n2786 ) == ( bv_8_148_n102 )  ;
assign n2788 = in[31:24] ;
assign n2789 =  ( n2788 ) == ( bv_8_147_n393 )  ;
assign n2790 = in[31:24] ;
assign n2791 =  ( n2790 ) == ( bv_8_146_n396 )  ;
assign n2792 = in[31:24] ;
assign n2793 =  ( n2792 ) == ( bv_8_145_n312 )  ;
assign n2794 = in[31:24] ;
assign n2795 =  ( n2794 ) == ( bv_8_144_n385 )  ;
assign n2796 = in[31:24] ;
assign n2797 =  ( n2796 ) == ( bv_8_143_n406 )  ;
assign n2798 = in[31:24] ;
assign n2799 =  ( n2798 ) == ( bv_8_142_n105 )  ;
assign n2800 = in[31:24] ;
assign n2801 =  ( n2800 ) == ( bv_8_141_n285 )  ;
assign n2802 = in[31:24] ;
assign n2803 =  ( n2802 ) == ( bv_8_140_n67 )  ;
assign n2804 = in[31:24] ;
assign n2805 =  ( n2804 ) == ( bv_8_139_n195 )  ;
assign n2806 = in[31:24] ;
assign n2807 =  ( n2806 ) == ( bv_8_138_n192 )  ;
assign n2808 = in[31:24] ;
assign n2809 =  ( n2808 ) == ( bv_8_137_n59 )  ;
assign n2810 = in[31:24] ;
assign n2811 =  ( n2810 ) == ( bv_8_136_n381 )  ;
assign n2812 = in[31:24] ;
assign n2813 =  ( n2812 ) == ( bv_8_135_n91 )  ;
assign n2814 = in[31:24] ;
assign n2815 =  ( n2814 ) == ( bv_8_134_n142 )  ;
assign n2816 = in[31:24] ;
assign n2817 =  ( n2816 ) == ( bv_8_133_n435 )  ;
assign n2818 = in[31:24] ;
assign n2819 =  ( n2818 ) == ( bv_8_132_n438 )  ;
assign n2820 = in[31:24] ;
assign n2821 =  ( n2820 ) == ( bv_8_131_n442 )  ;
assign n2822 = in[31:24] ;
assign n2823 =  ( n2822 ) == ( bv_8_130_n445 )  ;
assign n2824 = in[31:24] ;
assign n2825 =  ( n2824 ) == ( bv_8_129_n401 )  ;
assign n2826 = in[31:24] ;
assign n2827 =  ( n2826 ) == ( bv_8_128_n452 )  ;
assign n2828 = in[31:24] ;
assign n2829 =  ( n2828 ) == ( bv_8_127_n455 )  ;
assign n2830 = in[31:24] ;
assign n2831 =  ( n2830 ) == ( bv_8_126_n423 )  ;
assign n2832 = in[31:24] ;
assign n2833 =  ( n2832 ) == ( bv_8_125_n460 )  ;
assign n2834 = in[31:24] ;
assign n2835 =  ( n2834 ) == ( bv_8_124_n463 )  ;
assign n2836 = in[31:24] ;
assign n2837 =  ( n2836 ) == ( bv_8_123_n467 )  ;
assign n2838 = in[31:24] ;
assign n2839 =  ( n2838 ) == ( bv_8_122_n257 )  ;
assign n2840 = in[31:24] ;
assign n2841 =  ( n2840 ) == ( bv_8_121_n302 )  ;
assign n2842 = in[31:24] ;
assign n2843 =  ( n2842 ) == ( bv_8_120_n243 )  ;
assign n2844 = in[31:24] ;
assign n2845 =  ( n2844 ) == ( bv_8_119_n477 )  ;
assign n2846 = in[31:24] ;
assign n2847 =  ( n2846 ) == ( bv_8_118_n480 )  ;
assign n2848 = in[31:24] ;
assign n2849 =  ( n2848 ) == ( bv_8_117_n484 )  ;
assign n2850 = in[31:24] ;
assign n2851 =  ( n2850 ) == ( bv_8_116_n211 )  ;
assign n2852 = in[31:24] ;
assign n2853 =  ( n2852 ) == ( bv_8_115_n408 )  ;
assign n2854 = in[31:24] ;
assign n2855 =  ( n2854 ) == ( bv_8_114_n491 )  ;
assign n2856 = in[31:24] ;
assign n2857 =  ( n2856 ) == ( bv_8_113_n495 )  ;
assign n2858 = in[31:24] ;
assign n2859 =  ( n2858 ) == ( bv_8_112_n188 )  ;
assign n2860 = in[31:24] ;
assign n2861 =  ( n2860 ) == ( bv_8_111_n501 )  ;
assign n2862 = in[31:24] ;
assign n2863 =  ( n2862 ) == ( bv_8_110_n504 )  ;
assign n2864 = in[31:24] ;
assign n2865 =  ( n2864 ) == ( bv_8_109_n289 )  ;
assign n2866 = in[31:24] ;
assign n2867 =  ( n2866 ) == ( bv_8_108_n272 )  ;
assign n2868 = in[31:24] ;
assign n2869 =  ( n2868 ) == ( bv_8_107_n513 )  ;
assign n2870 = in[31:24] ;
assign n2871 =  ( n2870 ) == ( bv_8_106_n516 )  ;
assign n2872 = in[31:24] ;
assign n2873 =  ( n2872 ) == ( bv_8_105_n113 )  ;
assign n2874 = in[31:24] ;
assign n2875 =  ( n2874 ) == ( bv_8_104_n39 )  ;
assign n2876 = in[31:24] ;
assign n2877 =  ( n2876 ) == ( bv_8_103_n525 )  ;
assign n2878 = in[31:24] ;
assign n2879 =  ( n2878 ) == ( bv_8_102_n176 )  ;
assign n2880 = in[31:24] ;
assign n2881 =  ( n2880 ) == ( bv_8_101_n261 )  ;
assign n2882 = in[31:24] ;
assign n2883 =  ( n2882 ) == ( bv_8_100_n417 )  ;
assign n2884 = in[31:24] ;
assign n2885 =  ( n2884 ) == ( bv_8_99_n537 )  ;
assign n2886 = in[31:24] ;
assign n2887 =  ( n2886 ) == ( bv_8_98_n316 )  ;
assign n2888 = in[31:24] ;
assign n2889 =  ( n2888 ) == ( bv_8_97_n157 )  ;
assign n2890 = in[31:24] ;
assign n2891 =  ( n2890 ) == ( bv_8_96_n404 )  ;
assign n2892 = in[31:24] ;
assign n2893 =  ( n2892 ) == ( bv_8_95_n440 )  ;
assign n2894 = in[31:24] ;
assign n2895 =  ( n2894 ) == ( bv_8_94_n363 )  ;
assign n2896 = in[31:24] ;
assign n2897 =  ( n2896 ) == ( bv_8_93_n414 )  ;
assign n2898 = in[31:24] ;
assign n2899 =  ( n2898 ) == ( bv_8_92_n328 )  ;
assign n2900 = in[31:24] ;
assign n2901 =  ( n2900 ) == ( bv_8_91_n557 )  ;
assign n2902 = in[31:24] ;
assign n2903 =  ( n2902 ) == ( bv_8_90_n561 )  ;
assign n2904 = in[31:24] ;
assign n2905 =  ( n2904 ) == ( bv_8_89_n564 )  ;
assign n2906 = in[31:24] ;
assign n2907 =  ( n2906 ) == ( bv_8_88_n549 )  ;
assign n2908 = in[31:24] ;
assign n2909 =  ( n2908 ) == ( bv_8_87_n150 )  ;
assign n2910 = in[31:24] ;
assign n2911 =  ( n2910 ) == ( bv_8_86_n268 )  ;
assign n2912 = in[31:24] ;
assign n2913 =  ( n2912 ) == ( bv_8_85_n79 )  ;
assign n2914 = in[31:24] ;
assign n2915 =  ( n2914 ) == ( bv_8_84_n15 )  ;
assign n2916 = in[31:24] ;
assign n2917 =  ( n2916 ) == ( bv_8_83_n578 )  ;
assign n2918 = in[31:24] ;
assign n2919 =  ( n2918 ) == ( bv_8_82_n581 )  ;
assign n2920 = in[31:24] ;
assign n2921 =  ( n2920 ) == ( bv_8_81_n499 )  ;
assign n2922 = in[31:24] ;
assign n2923 =  ( n2922 ) == ( bv_8_80_n511 )  ;
assign n2924 = in[31:24] ;
assign n2925 =  ( n2924 ) == ( bv_8_79_n398 )  ;
assign n2926 = in[31:24] ;
assign n2927 =  ( n2926 ) == ( bv_8_78_n280 )  ;
assign n2928 = in[31:24] ;
assign n2929 =  ( n2928 ) == ( bv_8_77_n532 )  ;
assign n2930 = in[31:24] ;
assign n2931 =  ( n2930 ) == ( bv_8_76_n552 )  ;
assign n2932 = in[31:24] ;
assign n2933 =  ( n2932 ) == ( bv_8_75_n203 )  ;
assign n2934 = in[31:24] ;
assign n2935 =  ( n2934 ) == ( bv_8_74_n555 )  ;
assign n2936 = in[31:24] ;
assign n2937 =  ( n2936 ) == ( bv_8_73_n339 )  ;
assign n2938 = in[31:24] ;
assign n2939 =  ( n2938 ) == ( bv_8_72_n172 )  ;
assign n2940 = in[31:24] ;
assign n2941 =  ( n2940 ) == ( bv_8_71_n608 )  ;
assign n2942 = in[31:24] ;
assign n2943 =  ( n2942 ) == ( bv_8_70_n377 )  ;
assign n2944 = in[31:24] ;
assign n2945 =  ( n2944 ) == ( bv_8_69_n523 )  ;
assign n2946 = in[31:24] ;
assign n2947 =  ( n2946 ) == ( bv_8_68_n433 )  ;
assign n2948 = in[31:24] ;
assign n2949 =  ( n2948 ) == ( bv_8_67_n535 )  ;
assign n2950 = in[31:24] ;
assign n2951 =  ( n2950 ) == ( bv_8_66_n43 )  ;
assign n2952 = in[31:24] ;
assign n2953 =  ( n2952 ) == ( bv_8_65_n35 )  ;
assign n2954 = in[31:24] ;
assign n2955 =  ( n2954 ) == ( bv_8_64_n493 )  ;
assign n2956 = in[31:24] ;
assign n2957 =  ( n2956 ) == ( bv_8_63_n629 )  ;
assign n2958 = in[31:24] ;
assign n2959 =  ( n2958 ) == ( bv_8_62_n184 )  ;
assign n2960 = in[31:24] ;
assign n2961 =  ( n2960 ) == ( bv_8_61_n420 )  ;
assign n2962 = in[31:24] ;
assign n2963 =  ( n2962 ) == ( bv_8_60_n508 )  ;
assign n2964 = in[31:24] ;
assign n2965 =  ( n2964 ) == ( bv_8_59_n604 )  ;
assign n2966 = in[31:24] ;
assign n2967 =  ( n2966 ) == ( bv_8_58_n347 )  ;
assign n2968 = in[31:24] ;
assign n2969 =  ( n2968 ) == ( bv_8_57_n559 )  ;
assign n2970 = in[31:24] ;
assign n2971 =  ( n2970 ) == ( bv_8_56_n482 )  ;
assign n2972 = in[31:24] ;
assign n2973 =  ( n2972 ) == ( bv_8_55_n293 )  ;
assign n2974 = in[31:24] ;
assign n2975 =  ( n2974 ) == ( bv_8_54_n651 )  ;
assign n2976 = in[31:24] ;
assign n2977 =  ( n2976 ) == ( bv_8_53_n153 )  ;
assign n2978 = in[31:24] ;
assign n2979 =  ( n2978 ) == ( bv_8_52_n657 )  ;
assign n2980 = in[31:24] ;
assign n2981 =  ( n2980 ) == ( bv_8_51_n529 )  ;
assign n2982 = in[31:24] ;
assign n2983 =  ( n2982 ) == ( bv_8_50_n350 )  ;
assign n2984 = in[31:24] ;
assign n2985 =  ( n2984 ) == ( bv_8_49_n666 )  ;
assign n2986 = in[31:24] ;
assign n2987 =  ( n2986 ) == ( bv_8_48_n669 )  ;
assign n2988 = in[31:24] ;
assign n2989 =  ( n2988 ) == ( bv_8_47_n592 )  ;
assign n2990 = in[31:24] ;
assign n2991 =  ( n2990 ) == ( bv_8_46_n236 )  ;
assign n2992 = in[31:24] ;
assign n2993 =  ( n2992 ) == ( bv_8_45_n27 )  ;
assign n2994 = in[31:24] ;
assign n2995 =  ( n2994 ) == ( bv_8_44_n622 )  ;
assign n2996 = in[31:24] ;
assign n2997 =  ( n2996 ) == ( bv_8_43_n682 )  ;
assign n2998 = in[31:24] ;
assign n2999 =  ( n2998 ) == ( bv_8_42_n388 )  ;
assign n3000 = in[31:24] ;
assign n3001 =  ( n3000 ) == ( bv_8_41_n597 )  ;
assign n3002 = in[31:24] ;
assign n3003 =  ( n3002 ) == ( bv_8_40_n75 )  ;
assign n3004 = in[31:24] ;
assign n3005 =  ( n3004 ) == ( bv_8_39_n635 )  ;
assign n3006 = in[31:24] ;
assign n3007 =  ( n3006 ) == ( bv_8_38_n693 )  ;
assign n3008 = in[31:24] ;
assign n3009 =  ( n3008 ) == ( bv_8_37_n240 )  ;
assign n3010 = in[31:24] ;
assign n3011 =  ( n3010 ) == ( bv_8_36_n331 )  ;
assign n3012 = in[31:24] ;
assign n3013 =  ( n3012 ) == ( bv_8_35_n664 )  ;
assign n3014 = in[31:24] ;
assign n3015 =  ( n3014 ) == ( bv_8_34_n391 )  ;
assign n3016 = in[31:24] ;
assign n3017 =  ( n3016 ) == ( bv_8_33_n469 )  ;
assign n3018 = in[31:24] ;
assign n3019 =  ( n3018 ) == ( bv_8_32_n576 )  ;
assign n3020 = in[31:24] ;
assign n3021 =  ( n3020 ) == ( bv_8_31_n207 )  ;
assign n3022 = in[31:24] ;
assign n3023 =  ( n3022 ) == ( bv_8_30_n94 )  ;
assign n3024 = in[31:24] ;
assign n3025 =  ( n3024 ) == ( bv_8_29_n134 )  ;
assign n3026 = in[31:24] ;
assign n3027 =  ( n3026 ) == ( bv_8_28_n232 )  ;
assign n3028 = in[31:24] ;
assign n3029 =  ( n3028 ) == ( bv_8_27_n616 )  ;
assign n3030 = in[31:24] ;
assign n3031 =  ( n3030 ) == ( bv_8_26_n619 )  ;
assign n3032 = in[31:24] ;
assign n3033 =  ( n3032 ) == ( bv_8_25_n411 )  ;
assign n3034 = in[31:24] ;
assign n3035 =  ( n3034 ) == ( bv_8_24_n659 )  ;
assign n3036 = in[31:24] ;
assign n3037 =  ( n3036 ) == ( bv_8_23_n430 )  ;
assign n3038 = in[31:24] ;
assign n3039 =  ( n3038 ) == ( bv_8_22_n7 )  ;
assign n3040 = in[31:24] ;
assign n3041 =  ( n3040 ) == ( bv_8_21_n674 )  ;
assign n3042 = in[31:24] ;
assign n3043 =  ( n3042 ) == ( bv_8_20_n369 )  ;
assign n3044 = in[31:24] ;
assign n3045 =  ( n3044 ) == ( bv_8_19_n447 )  ;
assign n3046 = in[31:24] ;
assign n3047 =  ( n3046 ) == ( bv_8_18_n644 )  ;
assign n3048 = in[31:24] ;
assign n3049 =  ( n3048 ) == ( bv_8_17_n117 )  ;
assign n3050 = in[31:24] ;
assign n3051 =  ( n3050 ) == ( bv_8_16_n465 )  ;
assign n3052 = in[31:24] ;
assign n3053 =  ( n3052 ) == ( bv_8_15_n23 )  ;
assign n3054 = in[31:24] ;
assign n3055 =  ( n3054 ) == ( bv_8_14_n161 )  ;
assign n3056 = in[31:24] ;
assign n3057 =  ( n3056 ) == ( bv_8_13_n55 )  ;
assign n3058 = in[31:24] ;
assign n3059 =  ( n3058 ) == ( bv_8_12_n450 )  ;
assign n3060 = in[31:24] ;
assign n3061 =  ( n3060 ) == ( bv_8_11_n359 )  ;
assign n3062 = in[31:24] ;
assign n3063 =  ( n3062 ) == ( bv_8_10_n343 )  ;
assign n3064 = in[31:24] ;
assign n3065 =  ( n3064 ) == ( bv_8_9_n627 )  ;
assign n3066 = in[31:24] ;
assign n3067 =  ( n3066 ) == ( bv_8_8_n250 )  ;
assign n3068 = in[31:24] ;
assign n3069 =  ( n3068 ) == ( bv_8_7_n647 )  ;
assign n3070 = in[31:24] ;
assign n3071 =  ( n3070 ) == ( bv_8_6_n335 )  ;
assign n3072 = in[31:24] ;
assign n3073 =  ( n3072 ) == ( bv_8_5_n653 )  ;
assign n3074 = in[31:24] ;
assign n3075 =  ( n3074 ) == ( bv_8_4_n671 )  ;
assign n3076 = in[31:24] ;
assign n3077 =  ( n3076 ) == ( bv_8_3_n168 )  ;
assign n3078 = in[31:24] ;
assign n3079 =  ( n3078 ) == ( bv_8_2_n518 )  ;
assign n3080 = in[31:24] ;
assign n3081 =  ( n3080 ) == ( bv_8_1_n753 )  ;
assign n3082 = in[31:24] ;
assign n3083 =  ( n3082 ) == ( bv_8_0_n583 )  ;
assign n3084 =  ( n3083 ) ? ( bv_8_99_n537 ) : ( bv_8_0_n583 ) ;
assign n3085 =  ( n3081 ) ? ( bv_8_124_n463 ) : ( n3084 ) ;
assign n3086 =  ( n3079 ) ? ( bv_8_119_n477 ) : ( n3085 ) ;
assign n3087 =  ( n3077 ) ? ( bv_8_123_n467 ) : ( n3086 ) ;
assign n3088 =  ( n3075 ) ? ( bv_8_242_n57 ) : ( n3087 ) ;
assign n3089 =  ( n3073 ) ? ( bv_8_107_n513 ) : ( n3088 ) ;
assign n3090 =  ( n3071 ) ? ( bv_8_111_n501 ) : ( n3089 ) ;
assign n3091 =  ( n3069 ) ? ( bv_8_197_n226 ) : ( n3090 ) ;
assign n3092 =  ( n3067 ) ? ( bv_8_48_n669 ) : ( n3091 ) ;
assign n3093 =  ( n3065 ) ? ( bv_8_1_n753 ) : ( n3092 ) ;
assign n3094 =  ( n3063 ) ? ( bv_8_103_n525 ) : ( n3093 ) ;
assign n3095 =  ( n3061 ) ? ( bv_8_43_n682 ) : ( n3094 ) ;
assign n3096 =  ( n3059 ) ? ( bv_8_254_n9 ) : ( n3095 ) ;
assign n3097 =  ( n3057 ) ? ( bv_8_215_n159 ) : ( n3096 ) ;
assign n3098 =  ( n3055 ) ? ( bv_8_171_n314 ) : ( n3097 ) ;
assign n3099 =  ( n3053 ) ? ( bv_8_118_n480 ) : ( n3098 ) ;
assign n3100 =  ( n3051 ) ? ( bv_8_202_n209 ) : ( n3099 ) ;
assign n3101 =  ( n3049 ) ? ( bv_8_130_n445 ) : ( n3100 ) ;
assign n3102 =  ( n3047 ) ? ( bv_8_201_n213 ) : ( n3101 ) ;
assign n3103 =  ( n3045 ) ? ( bv_8_125_n460 ) : ( n3102 ) ;
assign n3104 =  ( n3043 ) ? ( bv_8_250_n25 ) : ( n3103 ) ;
assign n3105 =  ( n3041 ) ? ( bv_8_89_n564 ) : ( n3104 ) ;
assign n3106 =  ( n3039 ) ? ( bv_8_71_n608 ) : ( n3105 ) ;
assign n3107 =  ( n3037 ) ? ( bv_8_240_n65 ) : ( n3106 ) ;
assign n3108 =  ( n3035 ) ? ( bv_8_173_n306 ) : ( n3107 ) ;
assign n3109 =  ( n3033 ) ? ( bv_8_212_n170 ) : ( n3108 ) ;
assign n3110 =  ( n3031 ) ? ( bv_8_162_n345 ) : ( n3109 ) ;
assign n3111 =  ( n3029 ) ? ( bv_8_175_n300 ) : ( n3110 ) ;
assign n3112 =  ( n3027 ) ? ( bv_8_156_n365 ) : ( n3111 ) ;
assign n3113 =  ( n3025 ) ? ( bv_8_164_n337 ) : ( n3112 ) ;
assign n3114 =  ( n3023 ) ? ( bv_8_114_n491 ) : ( n3113 ) ;
assign n3115 =  ( n3021 ) ? ( bv_8_192_n245 ) : ( n3114 ) ;
assign n3116 =  ( n3019 ) ? ( bv_8_183_n274 ) : ( n3115 ) ;
assign n3117 =  ( n3017 ) ? ( bv_8_253_n13 ) : ( n3116 ) ;
assign n3118 =  ( n3015 ) ? ( bv_8_147_n393 ) : ( n3117 ) ;
assign n3119 =  ( n3013 ) ? ( bv_8_38_n693 ) : ( n3118 ) ;
assign n3120 =  ( n3011 ) ? ( bv_8_54_n651 ) : ( n3119 ) ;
assign n3121 =  ( n3009 ) ? ( bv_8_63_n629 ) : ( n3120 ) ;
assign n3122 =  ( n3007 ) ? ( bv_8_247_n37 ) : ( n3121 ) ;
assign n3123 =  ( n3005 ) ? ( bv_8_204_n201 ) : ( n3122 ) ;
assign n3124 =  ( n3003 ) ? ( bv_8_52_n657 ) : ( n3123 ) ;
assign n3125 =  ( n3001 ) ? ( bv_8_165_n333 ) : ( n3124 ) ;
assign n3126 =  ( n2999 ) ? ( bv_8_229_n107 ) : ( n3125 ) ;
assign n3127 =  ( n2997 ) ? ( bv_8_241_n61 ) : ( n3126 ) ;
assign n3128 =  ( n2995 ) ? ( bv_8_113_n495 ) : ( n3127 ) ;
assign n3129 =  ( n2993 ) ? ( bv_8_216_n155 ) : ( n3128 ) ;
assign n3130 =  ( n2991 ) ? ( bv_8_49_n666 ) : ( n3129 ) ;
assign n3131 =  ( n2989 ) ? ( bv_8_21_n674 ) : ( n3130 ) ;
assign n3132 =  ( n2987 ) ? ( bv_8_4_n671 ) : ( n3131 ) ;
assign n3133 =  ( n2985 ) ? ( bv_8_199_n219 ) : ( n3132 ) ;
assign n3134 =  ( n2983 ) ? ( bv_8_35_n664 ) : ( n3133 ) ;
assign n3135 =  ( n2981 ) ? ( bv_8_195_n234 ) : ( n3134 ) ;
assign n3136 =  ( n2979 ) ? ( bv_8_24_n659 ) : ( n3135 ) ;
assign n3137 =  ( n2977 ) ? ( bv_8_150_n383 ) : ( n3136 ) ;
assign n3138 =  ( n2975 ) ? ( bv_8_5_n653 ) : ( n3137 ) ;
assign n3139 =  ( n2973 ) ? ( bv_8_154_n371 ) : ( n3138 ) ;
assign n3140 =  ( n2971 ) ? ( bv_8_7_n647 ) : ( n3139 ) ;
assign n3141 =  ( n2969 ) ? ( bv_8_18_n644 ) : ( n3140 ) ;
assign n3142 =  ( n2967 ) ? ( bv_8_128_n452 ) : ( n3141 ) ;
assign n3143 =  ( n2965 ) ? ( bv_8_226_n119 ) : ( n3142 ) ;
assign n3144 =  ( n2963 ) ? ( bv_8_235_n85 ) : ( n3143 ) ;
assign n3145 =  ( n2961 ) ? ( bv_8_39_n635 ) : ( n3144 ) ;
assign n3146 =  ( n2959 ) ? ( bv_8_178_n291 ) : ( n3145 ) ;
assign n3147 =  ( n2957 ) ? ( bv_8_117_n484 ) : ( n3146 ) ;
assign n3148 =  ( n2955 ) ? ( bv_8_9_n627 ) : ( n3147 ) ;
assign n3149 =  ( n2953 ) ? ( bv_8_131_n442 ) : ( n3148 ) ;
assign n3150 =  ( n2951 ) ? ( bv_8_44_n622 ) : ( n3149 ) ;
assign n3151 =  ( n2949 ) ? ( bv_8_26_n619 ) : ( n3150 ) ;
assign n3152 =  ( n2947 ) ? ( bv_8_27_n616 ) : ( n3151 ) ;
assign n3153 =  ( n2945 ) ? ( bv_8_110_n504 ) : ( n3152 ) ;
assign n3154 =  ( n2943 ) ? ( bv_8_90_n561 ) : ( n3153 ) ;
assign n3155 =  ( n2941 ) ? ( bv_8_160_n352 ) : ( n3154 ) ;
assign n3156 =  ( n2939 ) ? ( bv_8_82_n581 ) : ( n3155 ) ;
assign n3157 =  ( n2937 ) ? ( bv_8_59_n604 ) : ( n3156 ) ;
assign n3158 =  ( n2935 ) ? ( bv_8_214_n163 ) : ( n3157 ) ;
assign n3159 =  ( n2933 ) ? ( bv_8_179_n287 ) : ( n3158 ) ;
assign n3160 =  ( n2931 ) ? ( bv_8_41_n597 ) : ( n3159 ) ;
assign n3161 =  ( n2929 ) ? ( bv_8_227_n115 ) : ( n3160 ) ;
assign n3162 =  ( n2927 ) ? ( bv_8_47_n592 ) : ( n3161 ) ;
assign n3163 =  ( n2925 ) ? ( bv_8_132_n438 ) : ( n3162 ) ;
assign n3164 =  ( n2923 ) ? ( bv_8_83_n578 ) : ( n3163 ) ;
assign n3165 =  ( n2921 ) ? ( bv_8_209_n182 ) : ( n3164 ) ;
assign n3166 =  ( n2919 ) ? ( bv_8_0_n583 ) : ( n3165 ) ;
assign n3167 =  ( n2917 ) ? ( bv_8_237_n77 ) : ( n3166 ) ;
assign n3168 =  ( n2915 ) ? ( bv_8_32_n576 ) : ( n3167 ) ;
assign n3169 =  ( n2913 ) ? ( bv_8_252_n17 ) : ( n3168 ) ;
assign n3170 =  ( n2911 ) ? ( bv_8_177_n295 ) : ( n3169 ) ;
assign n3171 =  ( n2909 ) ? ( bv_8_91_n557 ) : ( n3170 ) ;
assign n3172 =  ( n2907 ) ? ( bv_8_106_n516 ) : ( n3171 ) ;
assign n3173 =  ( n2905 ) ? ( bv_8_203_n205 ) : ( n3172 ) ;
assign n3174 =  ( n2903 ) ? ( bv_8_190_n252 ) : ( n3173 ) ;
assign n3175 =  ( n2901 ) ? ( bv_8_57_n559 ) : ( n3174 ) ;
assign n3176 =  ( n2899 ) ? ( bv_8_74_n555 ) : ( n3175 ) ;
assign n3177 =  ( n2897 ) ? ( bv_8_76_n552 ) : ( n3176 ) ;
assign n3178 =  ( n2895 ) ? ( bv_8_88_n549 ) : ( n3177 ) ;
assign n3179 =  ( n2893 ) ? ( bv_8_207_n190 ) : ( n3178 ) ;
assign n3180 =  ( n2891 ) ? ( bv_8_208_n186 ) : ( n3179 ) ;
assign n3181 =  ( n2889 ) ? ( bv_8_239_n69 ) : ( n3180 ) ;
assign n3182 =  ( n2887 ) ? ( bv_8_170_n318 ) : ( n3181 ) ;
assign n3183 =  ( n2885 ) ? ( bv_8_251_n21 ) : ( n3182 ) ;
assign n3184 =  ( n2883 ) ? ( bv_8_67_n535 ) : ( n3183 ) ;
assign n3185 =  ( n2881 ) ? ( bv_8_77_n532 ) : ( n3184 ) ;
assign n3186 =  ( n2879 ) ? ( bv_8_51_n529 ) : ( n3185 ) ;
assign n3187 =  ( n2877 ) ? ( bv_8_133_n435 ) : ( n3186 ) ;
assign n3188 =  ( n2875 ) ? ( bv_8_69_n523 ) : ( n3187 ) ;
assign n3189 =  ( n2873 ) ? ( bv_8_249_n29 ) : ( n3188 ) ;
assign n3190 =  ( n2871 ) ? ( bv_8_2_n518 ) : ( n3189 ) ;
assign n3191 =  ( n2869 ) ? ( bv_8_127_n455 ) : ( n3190 ) ;
assign n3192 =  ( n2867 ) ? ( bv_8_80_n511 ) : ( n3191 ) ;
assign n3193 =  ( n2865 ) ? ( bv_8_60_n508 ) : ( n3192 ) ;
assign n3194 =  ( n2863 ) ? ( bv_8_159_n355 ) : ( n3193 ) ;
assign n3195 =  ( n2861 ) ? ( bv_8_168_n323 ) : ( n3194 ) ;
assign n3196 =  ( n2859 ) ? ( bv_8_81_n499 ) : ( n3195 ) ;
assign n3197 =  ( n2857 ) ? ( bv_8_163_n341 ) : ( n3196 ) ;
assign n3198 =  ( n2855 ) ? ( bv_8_64_n493 ) : ( n3197 ) ;
assign n3199 =  ( n2853 ) ? ( bv_8_143_n406 ) : ( n3198 ) ;
assign n3200 =  ( n2851 ) ? ( bv_8_146_n396 ) : ( n3199 ) ;
assign n3201 =  ( n2849 ) ? ( bv_8_157_n361 ) : ( n3200 ) ;
assign n3202 =  ( n2847 ) ? ( bv_8_56_n482 ) : ( n3201 ) ;
assign n3203 =  ( n2845 ) ? ( bv_8_245_n45 ) : ( n3202 ) ;
assign n3204 =  ( n2843 ) ? ( bv_8_188_n259 ) : ( n3203 ) ;
assign n3205 =  ( n2841 ) ? ( bv_8_182_n278 ) : ( n3204 ) ;
assign n3206 =  ( n2839 ) ? ( bv_8_218_n148 ) : ( n3205 ) ;
assign n3207 =  ( n2837 ) ? ( bv_8_33_n469 ) : ( n3206 ) ;
assign n3208 =  ( n2835 ) ? ( bv_8_16_n465 ) : ( n3207 ) ;
assign n3209 =  ( n2833 ) ? ( bv_8_255_n5 ) : ( n3208 ) ;
assign n3210 =  ( n2831 ) ? ( bv_8_243_n53 ) : ( n3209 ) ;
assign n3211 =  ( n2829 ) ? ( bv_8_210_n178 ) : ( n3210 ) ;
assign n3212 =  ( n2827 ) ? ( bv_8_205_n197 ) : ( n3211 ) ;
assign n3213 =  ( n2825 ) ? ( bv_8_12_n450 ) : ( n3212 ) ;
assign n3214 =  ( n2823 ) ? ( bv_8_19_n447 ) : ( n3213 ) ;
assign n3215 =  ( n2821 ) ? ( bv_8_236_n81 ) : ( n3214 ) ;
assign n3216 =  ( n2819 ) ? ( bv_8_95_n440 ) : ( n3215 ) ;
assign n3217 =  ( n2817 ) ? ( bv_8_151_n379 ) : ( n3216 ) ;
assign n3218 =  ( n2815 ) ? ( bv_8_68_n433 ) : ( n3217 ) ;
assign n3219 =  ( n2813 ) ? ( bv_8_23_n430 ) : ( n3218 ) ;
assign n3220 =  ( n2811 ) ? ( bv_8_196_n230 ) : ( n3219 ) ;
assign n3221 =  ( n2809 ) ? ( bv_8_167_n326 ) : ( n3220 ) ;
assign n3222 =  ( n2807 ) ? ( bv_8_126_n423 ) : ( n3221 ) ;
assign n3223 =  ( n2805 ) ? ( bv_8_61_n420 ) : ( n3222 ) ;
assign n3224 =  ( n2803 ) ? ( bv_8_100_n417 ) : ( n3223 ) ;
assign n3225 =  ( n2801 ) ? ( bv_8_93_n414 ) : ( n3224 ) ;
assign n3226 =  ( n2799 ) ? ( bv_8_25_n411 ) : ( n3225 ) ;
assign n3227 =  ( n2797 ) ? ( bv_8_115_n408 ) : ( n3226 ) ;
assign n3228 =  ( n2795 ) ? ( bv_8_96_n404 ) : ( n3227 ) ;
assign n3229 =  ( n2793 ) ? ( bv_8_129_n401 ) : ( n3228 ) ;
assign n3230 =  ( n2791 ) ? ( bv_8_79_n398 ) : ( n3229 ) ;
assign n3231 =  ( n2789 ) ? ( bv_8_220_n140 ) : ( n3230 ) ;
assign n3232 =  ( n2787 ) ? ( bv_8_34_n391 ) : ( n3231 ) ;
assign n3233 =  ( n2785 ) ? ( bv_8_42_n388 ) : ( n3232 ) ;
assign n3234 =  ( n2783 ) ? ( bv_8_144_n385 ) : ( n3233 ) ;
assign n3235 =  ( n2781 ) ? ( bv_8_136_n381 ) : ( n3234 ) ;
assign n3236 =  ( n2779 ) ? ( bv_8_70_n377 ) : ( n3235 ) ;
assign n3237 =  ( n2777 ) ? ( bv_8_238_n73 ) : ( n3236 ) ;
assign n3238 =  ( n2775 ) ? ( bv_8_184_n270 ) : ( n3237 ) ;
assign n3239 =  ( n2773 ) ? ( bv_8_20_n369 ) : ( n3238 ) ;
assign n3240 =  ( n2771 ) ? ( bv_8_222_n132 ) : ( n3239 ) ;
assign n3241 =  ( n2769 ) ? ( bv_8_94_n363 ) : ( n3240 ) ;
assign n3242 =  ( n2767 ) ? ( bv_8_11_n359 ) : ( n3241 ) ;
assign n3243 =  ( n2765 ) ? ( bv_8_219_n144 ) : ( n3242 ) ;
assign n3244 =  ( n2763 ) ? ( bv_8_224_n126 ) : ( n3243 ) ;
assign n3245 =  ( n2761 ) ? ( bv_8_50_n350 ) : ( n3244 ) ;
assign n3246 =  ( n2759 ) ? ( bv_8_58_n347 ) : ( n3245 ) ;
assign n3247 =  ( n2757 ) ? ( bv_8_10_n343 ) : ( n3246 ) ;
assign n3248 =  ( n2755 ) ? ( bv_8_73_n339 ) : ( n3247 ) ;
assign n3249 =  ( n2753 ) ? ( bv_8_6_n335 ) : ( n3248 ) ;
assign n3250 =  ( n2751 ) ? ( bv_8_36_n331 ) : ( n3249 ) ;
assign n3251 =  ( n2749 ) ? ( bv_8_92_n328 ) : ( n3250 ) ;
assign n3252 =  ( n2747 ) ? ( bv_8_194_n238 ) : ( n3251 ) ;
assign n3253 =  ( n2745 ) ? ( bv_8_211_n174 ) : ( n3252 ) ;
assign n3254 =  ( n2743 ) ? ( bv_8_172_n310 ) : ( n3253 ) ;
assign n3255 =  ( n2741 ) ? ( bv_8_98_n316 ) : ( n3254 ) ;
assign n3256 =  ( n2739 ) ? ( bv_8_145_n312 ) : ( n3255 ) ;
assign n3257 =  ( n2737 ) ? ( bv_8_149_n308 ) : ( n3256 ) ;
assign n3258 =  ( n2735 ) ? ( bv_8_228_n111 ) : ( n3257 ) ;
assign n3259 =  ( n2733 ) ? ( bv_8_121_n302 ) : ( n3258 ) ;
assign n3260 =  ( n2731 ) ? ( bv_8_231_n100 ) : ( n3259 ) ;
assign n3261 =  ( n2729 ) ? ( bv_8_200_n216 ) : ( n3260 ) ;
assign n3262 =  ( n2727 ) ? ( bv_8_55_n293 ) : ( n3261 ) ;
assign n3263 =  ( n2725 ) ? ( bv_8_109_n289 ) : ( n3262 ) ;
assign n3264 =  ( n2723 ) ? ( bv_8_141_n285 ) : ( n3263 ) ;
assign n3265 =  ( n2721 ) ? ( bv_8_213_n166 ) : ( n3264 ) ;
assign n3266 =  ( n2719 ) ? ( bv_8_78_n280 ) : ( n3265 ) ;
assign n3267 =  ( n2717 ) ? ( bv_8_169_n276 ) : ( n3266 ) ;
assign n3268 =  ( n2715 ) ? ( bv_8_108_n272 ) : ( n3267 ) ;
assign n3269 =  ( n2713 ) ? ( bv_8_86_n268 ) : ( n3268 ) ;
assign n3270 =  ( n2711 ) ? ( bv_8_244_n49 ) : ( n3269 ) ;
assign n3271 =  ( n2709 ) ? ( bv_8_234_n89 ) : ( n3270 ) ;
assign n3272 =  ( n2707 ) ? ( bv_8_101_n261 ) : ( n3271 ) ;
assign n3273 =  ( n2705 ) ? ( bv_8_122_n257 ) : ( n3272 ) ;
assign n3274 =  ( n2703 ) ? ( bv_8_174_n254 ) : ( n3273 ) ;
assign n3275 =  ( n2701 ) ? ( bv_8_8_n250 ) : ( n3274 ) ;
assign n3276 =  ( n2699 ) ? ( bv_8_186_n247 ) : ( n3275 ) ;
assign n3277 =  ( n2697 ) ? ( bv_8_120_n243 ) : ( n3276 ) ;
assign n3278 =  ( n2695 ) ? ( bv_8_37_n240 ) : ( n3277 ) ;
assign n3279 =  ( n2693 ) ? ( bv_8_46_n236 ) : ( n3278 ) ;
assign n3280 =  ( n2691 ) ? ( bv_8_28_n232 ) : ( n3279 ) ;
assign n3281 =  ( n2689 ) ? ( bv_8_166_n228 ) : ( n3280 ) ;
assign n3282 =  ( n2687 ) ? ( bv_8_180_n224 ) : ( n3281 ) ;
assign n3283 =  ( n2685 ) ? ( bv_8_198_n221 ) : ( n3282 ) ;
assign n3284 =  ( n2683 ) ? ( bv_8_232_n96 ) : ( n3283 ) ;
assign n3285 =  ( n2681 ) ? ( bv_8_221_n136 ) : ( n3284 ) ;
assign n3286 =  ( n2679 ) ? ( bv_8_116_n211 ) : ( n3285 ) ;
assign n3287 =  ( n2677 ) ? ( bv_8_31_n207 ) : ( n3286 ) ;
assign n3288 =  ( n2675 ) ? ( bv_8_75_n203 ) : ( n3287 ) ;
assign n3289 =  ( n2673 ) ? ( bv_8_189_n199 ) : ( n3288 ) ;
assign n3290 =  ( n2671 ) ? ( bv_8_139_n195 ) : ( n3289 ) ;
assign n3291 =  ( n2669 ) ? ( bv_8_138_n192 ) : ( n3290 ) ;
assign n3292 =  ( n2667 ) ? ( bv_8_112_n188 ) : ( n3291 ) ;
assign n3293 =  ( n2665 ) ? ( bv_8_62_n184 ) : ( n3292 ) ;
assign n3294 =  ( n2663 ) ? ( bv_8_181_n180 ) : ( n3293 ) ;
assign n3295 =  ( n2661 ) ? ( bv_8_102_n176 ) : ( n3294 ) ;
assign n3296 =  ( n2659 ) ? ( bv_8_72_n172 ) : ( n3295 ) ;
assign n3297 =  ( n2657 ) ? ( bv_8_3_n168 ) : ( n3296 ) ;
assign n3298 =  ( n2655 ) ? ( bv_8_246_n41 ) : ( n3297 ) ;
assign n3299 =  ( n2653 ) ? ( bv_8_14_n161 ) : ( n3298 ) ;
assign n3300 =  ( n2651 ) ? ( bv_8_97_n157 ) : ( n3299 ) ;
assign n3301 =  ( n2649 ) ? ( bv_8_53_n153 ) : ( n3300 ) ;
assign n3302 =  ( n2647 ) ? ( bv_8_87_n150 ) : ( n3301 ) ;
assign n3303 =  ( n2645 ) ? ( bv_8_185_n146 ) : ( n3302 ) ;
assign n3304 =  ( n2643 ) ? ( bv_8_134_n142 ) : ( n3303 ) ;
assign n3305 =  ( n2641 ) ? ( bv_8_193_n138 ) : ( n3304 ) ;
assign n3306 =  ( n2639 ) ? ( bv_8_29_n134 ) : ( n3305 ) ;
assign n3307 =  ( n2637 ) ? ( bv_8_158_n130 ) : ( n3306 ) ;
assign n3308 =  ( n2635 ) ? ( bv_8_225_n123 ) : ( n3307 ) ;
assign n3309 =  ( n2633 ) ? ( bv_8_248_n33 ) : ( n3308 ) ;
assign n3310 =  ( n2631 ) ? ( bv_8_152_n121 ) : ( n3309 ) ;
assign n3311 =  ( n2629 ) ? ( bv_8_17_n117 ) : ( n3310 ) ;
assign n3312 =  ( n2627 ) ? ( bv_8_105_n113 ) : ( n3311 ) ;
assign n3313 =  ( n2625 ) ? ( bv_8_217_n109 ) : ( n3312 ) ;
assign n3314 =  ( n2623 ) ? ( bv_8_142_n105 ) : ( n3313 ) ;
assign n3315 =  ( n2621 ) ? ( bv_8_148_n102 ) : ( n3314 ) ;
assign n3316 =  ( n2619 ) ? ( bv_8_155_n98 ) : ( n3315 ) ;
assign n3317 =  ( n2617 ) ? ( bv_8_30_n94 ) : ( n3316 ) ;
assign n3318 =  ( n2615 ) ? ( bv_8_135_n91 ) : ( n3317 ) ;
assign n3319 =  ( n2613 ) ? ( bv_8_233_n87 ) : ( n3318 ) ;
assign n3320 =  ( n2611 ) ? ( bv_8_206_n83 ) : ( n3319 ) ;
assign n3321 =  ( n2609 ) ? ( bv_8_85_n79 ) : ( n3320 ) ;
assign n3322 =  ( n2607 ) ? ( bv_8_40_n75 ) : ( n3321 ) ;
assign n3323 =  ( n2605 ) ? ( bv_8_223_n71 ) : ( n3322 ) ;
assign n3324 =  ( n2603 ) ? ( bv_8_140_n67 ) : ( n3323 ) ;
assign n3325 =  ( n2601 ) ? ( bv_8_161_n63 ) : ( n3324 ) ;
assign n3326 =  ( n2599 ) ? ( bv_8_137_n59 ) : ( n3325 ) ;
assign n3327 =  ( n2597 ) ? ( bv_8_13_n55 ) : ( n3326 ) ;
assign n3328 =  ( n2595 ) ? ( bv_8_191_n51 ) : ( n3327 ) ;
assign n3329 =  ( n2593 ) ? ( bv_8_230_n47 ) : ( n3328 ) ;
assign n3330 =  ( n2591 ) ? ( bv_8_66_n43 ) : ( n3329 ) ;
assign n3331 =  ( n2589 ) ? ( bv_8_104_n39 ) : ( n3330 ) ;
assign n3332 =  ( n2587 ) ? ( bv_8_65_n35 ) : ( n3331 ) ;
assign n3333 =  ( n2585 ) ? ( bv_8_153_n31 ) : ( n3332 ) ;
assign n3334 =  ( n2583 ) ? ( bv_8_45_n27 ) : ( n3333 ) ;
assign n3335 =  ( n2581 ) ? ( bv_8_15_n23 ) : ( n3334 ) ;
assign n3336 =  ( n2579 ) ? ( bv_8_176_n19 ) : ( n3335 ) ;
assign n3337 =  ( n2577 ) ? ( bv_8_84_n15 ) : ( n3336 ) ;
assign n3338 =  ( n2575 ) ? ( bv_8_187_n11 ) : ( n3337 ) ;
assign n3339 =  ( n2573 ) ? ( bv_8_22_n7 ) : ( n3338 ) ;
assign n3340 =  ( n2571 ) ^ ( n3339 )  ;
assign n3341 =  { ( n2570 ) , ( n3340 ) }  ;
assign n3342 = in[127:120] ;
assign n3343 =  ( n3342 ) ^ ( rcon )  ;
assign n3344 = in[95:88] ;
assign n3345 =  ( n3343 ) ^ ( n3344 )  ;
assign n3346 =  ( n3345 ) ^ ( n1027 )  ;
assign n3347 =  { ( n3341 ) , ( n3346 ) }  ;
assign n3348 = in[119:112] ;
assign n3349 = in[87:80] ;
assign n3350 =  ( n3348 ) ^ ( n3349 )  ;
assign n3351 =  ( n3350 ) ^ ( n1797 )  ;
assign n3352 =  { ( n3347 ) , ( n3351 ) }  ;
assign n3353 = in[111:104] ;
assign n3354 = in[79:72] ;
assign n3355 =  ( n3353 ) ^ ( n3354 )  ;
assign n3356 =  ( n3355 ) ^ ( n2568 )  ;
assign n3357 =  { ( n3352 ) , ( n3356 ) }  ;
assign n3358 = in[103:96] ;
assign n3359 = in[71:64] ;
assign n3360 =  ( n3358 ) ^ ( n3359 )  ;
assign n3361 =  ( n3360 ) ^ ( n3339 )  ;
assign n3362 =  { ( n3357 ) , ( n3361 ) }  ;
assign n3363 = in[127:120] ;
assign n3364 =  ( n3363 ) ^ ( rcon )  ;
assign n3365 = in[95:88] ;
assign n3366 =  ( n3364 ) ^ ( n3365 )  ;
assign n3367 = in[63:56] ;
assign n3368 =  ( n3366 ) ^ ( n3367 )  ;
assign n3369 =  ( n3368 ) ^ ( n1027 )  ;
assign n3370 =  { ( n3362 ) , ( n3369 ) }  ;
assign n3371 = in[119:112] ;
assign n3372 = in[87:80] ;
assign n3373 =  ( n3371 ) ^ ( n3372 )  ;
assign n3374 = in[55:48] ;
assign n3375 =  ( n3373 ) ^ ( n3374 )  ;
assign n3376 =  ( n3375 ) ^ ( n1797 )  ;
assign n3377 =  { ( n3370 ) , ( n3376 ) }  ;
assign n3378 = in[111:104] ;
assign n3379 = in[79:72] ;
assign n3380 =  ( n3378 ) ^ ( n3379 )  ;
assign n3381 = in[47:40] ;
assign n3382 =  ( n3380 ) ^ ( n3381 )  ;
assign n3383 =  ( n3382 ) ^ ( n2568 )  ;
assign n3384 =  { ( n3377 ) , ( n3383 ) }  ;
assign n3385 = in[103:96] ;
assign n3386 = in[71:64] ;
assign n3387 =  ( n3385 ) ^ ( n3386 )  ;
assign n3388 = in[39:32] ;
assign n3389 =  ( n3387 ) ^ ( n3388 )  ;
assign n3390 =  ( n3389 ) ^ ( n3339 )  ;
assign n3391 =  { ( n3384 ) , ( n3390 ) }  ;
assign n3392 = in[127:120] ;
assign n3393 =  ( n3392 ) ^ ( rcon )  ;
assign n3394 = in[95:88] ;
assign n3395 =  ( n3393 ) ^ ( n3394 )  ;
assign n3396 = in[63:56] ;
assign n3397 =  ( n3395 ) ^ ( n3396 )  ;
assign n3398 = in[31:24] ;
assign n3399 =  ( n3397 ) ^ ( n3398 )  ;
assign n3400 =  ( n3399 ) ^ ( n1027 )  ;
assign n3401 =  { ( n3391 ) , ( n3400 ) }  ;
assign n3402 = in[119:112] ;
assign n3403 = in[87:80] ;
assign n3404 =  ( n3402 ) ^ ( n3403 )  ;
assign n3405 = in[55:48] ;
assign n3406 =  ( n3404 ) ^ ( n3405 )  ;
assign n3407 = in[23:16] ;
assign n3408 =  ( n3406 ) ^ ( n3407 )  ;
assign n3409 =  ( n3408 ) ^ ( n1797 )  ;
assign n3410 =  { ( n3401 ) , ( n3409 ) }  ;
assign n3411 = in[111:104] ;
assign n3412 = in[79:72] ;
assign n3413 =  ( n3411 ) ^ ( n3412 )  ;
assign n3414 = in[47:40] ;
assign n3415 =  ( n3413 ) ^ ( n3414 )  ;
assign n3416 = in[15:8] ;
assign n3417 =  ( n3415 ) ^ ( n3416 )  ;
assign n3418 =  ( n3417 ) ^ ( n2568 )  ;
assign n3419 =  { ( n3410 ) , ( n3418 ) }  ;
assign n3420 = in[103:96] ;
assign n3421 = in[71:64] ;
assign n3422 =  ( n3420 ) ^ ( n3421 )  ;
assign n3423 = in[39:32] ;
assign n3424 =  ( n3422 ) ^ ( n3423 )  ;
assign n3425 = in[7:0] ;
assign n3426 =  ( n3424 ) ^ ( n3425 )  ;
assign n3427 =  ( n3426 ) ^ ( n3339 )  ;
assign n3428 =  { ( n3419 ) , ( n3427 ) }  ;
assign n3429 =  ( bv_128_0_n1 ) + ( n3428 )  ;
always @(posedge clk) begin
   if(rst) begin
       __COUNTER_start__n0 <= 0;
   end
   else if(__ILA_bar_valid__) begin
       if ( __ILA_bar_decode_of_i1__ ) begin 
           __COUNTER_start__n0 <= 1; end
       else if( (__COUNTER_start__n0 >= 1 ) && ( __COUNTER_start__n0 < 255 )) begin
           __COUNTER_start__n0 <= __COUNTER_start__n0 + 1; end
       if (__ILA_bar_decode_of_i1__) begin
           in <= in ;
       end
       if (__ILA_bar_decode_of_i1__) begin
           rcon <= rcon ;
       end
       if (__ILA_bar_decode_of_i1__) begin
           out_1 <= n3429 ;
       end
   end
end
endmodule
