module NV_NVDLA_RT_csc2cmac_a(nvdla_core_clk, nvdla_core_rstn, sc2mac_wt_src_pvld, sc2mac_wt_src_mask, sc2mac_wt_src_data0, sc2mac_wt_src_data1, sc2mac_wt_src_data2, sc2mac_wt_src_data3, sc2mac_wt_src_data4, sc2mac_wt_src_data5, sc2mac_wt_src_data6, sc2mac_wt_src_data7, sc2mac_wt_src_data8, sc2mac_wt_src_data9, sc2mac_wt_src_data10, sc2mac_wt_src_data11, sc2mac_wt_src_data12, sc2mac_wt_src_data13, sc2mac_wt_src_data14, sc2mac_wt_src_data15, sc2mac_wt_src_data16, sc2mac_wt_src_data17, sc2mac_wt_src_data18, sc2mac_wt_src_data19, sc2mac_wt_src_data20, sc2mac_wt_src_data21, sc2mac_wt_src_data22, sc2mac_wt_src_data23, sc2mac_wt_src_data24, sc2mac_wt_src_data25, sc2mac_wt_src_data26, sc2mac_wt_src_data27, sc2mac_wt_src_data28, sc2mac_wt_src_data29, sc2mac_wt_src_data30, sc2mac_wt_src_data31, sc2mac_wt_src_data32, sc2mac_wt_src_data33, sc2mac_wt_src_data34, sc2mac_wt_src_data35, sc2mac_wt_src_data36, sc2mac_wt_src_data37, sc2mac_wt_src_data38, sc2mac_wt_src_data39, sc2mac_wt_src_data40, sc2mac_wt_src_data41, sc2mac_wt_src_data42, sc2mac_wt_src_data43, sc2mac_wt_src_data44, sc2mac_wt_src_data45, sc2mac_wt_src_data46, sc2mac_wt_src_data47, sc2mac_wt_src_data48, sc2mac_wt_src_data49, sc2mac_wt_src_data50, sc2mac_wt_src_data51, sc2mac_wt_src_data52, sc2mac_wt_src_data53, sc2mac_wt_src_data54, sc2mac_wt_src_data55, sc2mac_wt_src_data56, sc2mac_wt_src_data57, sc2mac_wt_src_data58, sc2mac_wt_src_data59, sc2mac_wt_src_data60, sc2mac_wt_src_data61, sc2mac_wt_src_data62, sc2mac_wt_src_data63, sc2mac_wt_src_data64, sc2mac_wt_src_data65, sc2mac_wt_src_data66, sc2mac_wt_src_data67, sc2mac_wt_src_data68, sc2mac_wt_src_data69, sc2mac_wt_src_data70, sc2mac_wt_src_data71, sc2mac_wt_src_data72, sc2mac_wt_src_data73, sc2mac_wt_src_data74, sc2mac_wt_src_data75, sc2mac_wt_src_data76, sc2mac_wt_src_data77, sc2mac_wt_src_data78, sc2mac_wt_src_data79, sc2mac_wt_src_data80, sc2mac_wt_src_data81, sc2mac_wt_src_data82, sc2mac_wt_src_data83, sc2mac_wt_src_data84, sc2mac_wt_src_data85, sc2mac_wt_src_data86, sc2mac_wt_src_data87, sc2mac_wt_src_data88, sc2mac_wt_src_data89, sc2mac_wt_src_data90, sc2mac_wt_src_data91, sc2mac_wt_src_data92, sc2mac_wt_src_data93, sc2mac_wt_src_data94, sc2mac_wt_src_data95, sc2mac_wt_src_data96, sc2mac_wt_src_data97, sc2mac_wt_src_data98, sc2mac_wt_src_data99, sc2mac_wt_src_data100, sc2mac_wt_src_data101, sc2mac_wt_src_data102, sc2mac_wt_src_data103, sc2mac_wt_src_data104, sc2mac_wt_src_data105, sc2mac_wt_src_data106, sc2mac_wt_src_data107, sc2mac_wt_src_data108, sc2mac_wt_src_data109, sc2mac_wt_src_data110, sc2mac_wt_src_data111, sc2mac_wt_src_data112, sc2mac_wt_src_data113, sc2mac_wt_src_data114, sc2mac_wt_src_data115, sc2mac_wt_src_data116, sc2mac_wt_src_data117, sc2mac_wt_src_data118, sc2mac_wt_src_data119, sc2mac_wt_src_data120, sc2mac_wt_src_data121, sc2mac_wt_src_data122, sc2mac_wt_src_data123, sc2mac_wt_src_data124, sc2mac_wt_src_data125, sc2mac_wt_src_data126, sc2mac_wt_src_data127, sc2mac_wt_src_sel, sc2mac_dat_src_pvld, sc2mac_dat_src_mask, sc2mac_dat_src_data0, sc2mac_dat_src_data1, sc2mac_dat_src_data2, sc2mac_dat_src_data3, sc2mac_dat_src_data4, sc2mac_dat_src_data5, sc2mac_dat_src_data6, sc2mac_dat_src_data7, sc2mac_dat_src_data8, sc2mac_dat_src_data9, sc2mac_dat_src_data10, sc2mac_dat_src_data11, sc2mac_dat_src_data12, sc2mac_dat_src_data13, sc2mac_dat_src_data14, sc2mac_dat_src_data15, sc2mac_dat_src_data16, sc2mac_dat_src_data17, sc2mac_dat_src_data18, sc2mac_dat_src_data19, sc2mac_dat_src_data20, sc2mac_dat_src_data21, sc2mac_dat_src_data22, sc2mac_dat_src_data23, sc2mac_dat_src_data24, sc2mac_dat_src_data25, sc2mac_dat_src_data26, sc2mac_dat_src_data27, sc2mac_dat_src_data28, sc2mac_dat_src_data29, sc2mac_dat_src_data30, sc2mac_dat_src_data31, sc2mac_dat_src_data32, sc2mac_dat_src_data33, sc2mac_dat_src_data34, sc2mac_dat_src_data35, sc2mac_dat_src_data36, sc2mac_dat_src_data37, sc2mac_dat_src_data38, sc2mac_dat_src_data39, sc2mac_dat_src_data40, sc2mac_dat_src_data41, sc2mac_dat_src_data42, sc2mac_dat_src_data43, sc2mac_dat_src_data44, sc2mac_dat_src_data45, sc2mac_dat_src_data46, sc2mac_dat_src_data47, sc2mac_dat_src_data48, sc2mac_dat_src_data49, sc2mac_dat_src_data50, sc2mac_dat_src_data51, sc2mac_dat_src_data52, sc2mac_dat_src_data53, sc2mac_dat_src_data54, sc2mac_dat_src_data55, sc2mac_dat_src_data56, sc2mac_dat_src_data57, sc2mac_dat_src_data58, sc2mac_dat_src_data59, sc2mac_dat_src_data60, sc2mac_dat_src_data61, sc2mac_dat_src_data62, sc2mac_dat_src_data63, sc2mac_dat_src_data64, sc2mac_dat_src_data65, sc2mac_dat_src_data66, sc2mac_dat_src_data67, sc2mac_dat_src_data68, sc2mac_dat_src_data69, sc2mac_dat_src_data70, sc2mac_dat_src_data71, sc2mac_dat_src_data72, sc2mac_dat_src_data73, sc2mac_dat_src_data74, sc2mac_dat_src_data75, sc2mac_dat_src_data76, sc2mac_dat_src_data77, sc2mac_dat_src_data78, sc2mac_dat_src_data79, sc2mac_dat_src_data80, sc2mac_dat_src_data81, sc2mac_dat_src_data82, sc2mac_dat_src_data83, sc2mac_dat_src_data84, sc2mac_dat_src_data85, sc2mac_dat_src_data86, sc2mac_dat_src_data87, sc2mac_dat_src_data88, sc2mac_dat_src_data89, sc2mac_dat_src_data90, sc2mac_dat_src_data91, sc2mac_dat_src_data92, sc2mac_dat_src_data93, sc2mac_dat_src_data94, sc2mac_dat_src_data95, sc2mac_dat_src_data96, sc2mac_dat_src_data97, sc2mac_dat_src_data98, sc2mac_dat_src_data99, sc2mac_dat_src_data100, sc2mac_dat_src_data101, sc2mac_dat_src_data102, sc2mac_dat_src_data103, sc2mac_dat_src_data104, sc2mac_dat_src_data105, sc2mac_dat_src_data106, sc2mac_dat_src_data107, sc2mac_dat_src_data108, sc2mac_dat_src_data109, sc2mac_dat_src_data110, sc2mac_dat_src_data111, sc2mac_dat_src_data112, sc2mac_dat_src_data113, sc2mac_dat_src_data114, sc2mac_dat_src_data115, sc2mac_dat_src_data116, sc2mac_dat_src_data117, sc2mac_dat_src_data118, sc2mac_dat_src_data119, sc2mac_dat_src_data120, sc2mac_dat_src_data121, sc2mac_dat_src_data122, sc2mac_dat_src_data123, sc2mac_dat_src_data124, sc2mac_dat_src_data125, sc2mac_dat_src_data126, sc2mac_dat_src_data127, sc2mac_dat_src_pd, sc2mac_wt_dst_pvld, sc2mac_wt_dst_mask, sc2mac_wt_dst_data0, sc2mac_wt_dst_data1, sc2mac_wt_dst_data2, sc2mac_wt_dst_data3, sc2mac_wt_dst_data4, sc2mac_wt_dst_data5, sc2mac_wt_dst_data6, sc2mac_wt_dst_data7, sc2mac_wt_dst_data8, sc2mac_wt_dst_data9, sc2mac_wt_dst_data10, sc2mac_wt_dst_data11, sc2mac_wt_dst_data12, sc2mac_wt_dst_data13, sc2mac_wt_dst_data14, sc2mac_wt_dst_data15, sc2mac_wt_dst_data16, sc2mac_wt_dst_data17, sc2mac_wt_dst_data18, sc2mac_wt_dst_data19, sc2mac_wt_dst_data20, sc2mac_wt_dst_data21, sc2mac_wt_dst_data22, sc2mac_wt_dst_data23, sc2mac_wt_dst_data24, sc2mac_wt_dst_data25, sc2mac_wt_dst_data26, sc2mac_wt_dst_data27, sc2mac_wt_dst_data28, sc2mac_wt_dst_data29, sc2mac_wt_dst_data30, sc2mac_wt_dst_data31, sc2mac_wt_dst_data32, sc2mac_wt_dst_data33, sc2mac_wt_dst_data34, sc2mac_wt_dst_data35, sc2mac_wt_dst_data36, sc2mac_wt_dst_data37, sc2mac_wt_dst_data38, sc2mac_wt_dst_data39, sc2mac_wt_dst_data40, sc2mac_wt_dst_data41, sc2mac_wt_dst_data42, sc2mac_wt_dst_data43, sc2mac_wt_dst_data44, sc2mac_wt_dst_data45, sc2mac_wt_dst_data46, sc2mac_wt_dst_data47, sc2mac_wt_dst_data48, sc2mac_wt_dst_data49, sc2mac_wt_dst_data50, sc2mac_wt_dst_data51, sc2mac_wt_dst_data52, sc2mac_wt_dst_data53, sc2mac_wt_dst_data54, sc2mac_wt_dst_data55, sc2mac_wt_dst_data56, sc2mac_wt_dst_data57, sc2mac_wt_dst_data58, sc2mac_wt_dst_data59, sc2mac_wt_dst_data60, sc2mac_wt_dst_data61, sc2mac_wt_dst_data62, sc2mac_wt_dst_data63, sc2mac_wt_dst_data64, sc2mac_wt_dst_data65, sc2mac_wt_dst_data66, sc2mac_wt_dst_data67, sc2mac_wt_dst_data68, sc2mac_wt_dst_data69, sc2mac_wt_dst_data70, sc2mac_wt_dst_data71, sc2mac_wt_dst_data72, sc2mac_wt_dst_data73, sc2mac_wt_dst_data74, sc2mac_wt_dst_data75, sc2mac_wt_dst_data76, sc2mac_wt_dst_data77, sc2mac_wt_dst_data78, sc2mac_wt_dst_data79, sc2mac_wt_dst_data80, sc2mac_wt_dst_data81, sc2mac_wt_dst_data82, sc2mac_wt_dst_data83, sc2mac_wt_dst_data84, sc2mac_wt_dst_data85, sc2mac_wt_dst_data86, sc2mac_wt_dst_data87, sc2mac_wt_dst_data88, sc2mac_wt_dst_data89, sc2mac_wt_dst_data90, sc2mac_wt_dst_data91, sc2mac_wt_dst_data92, sc2mac_wt_dst_data93, sc2mac_wt_dst_data94, sc2mac_wt_dst_data95, sc2mac_wt_dst_data96, sc2mac_wt_dst_data97, sc2mac_wt_dst_data98, sc2mac_wt_dst_data99, sc2mac_wt_dst_data100, sc2mac_wt_dst_data101, sc2mac_wt_dst_data102, sc2mac_wt_dst_data103, sc2mac_wt_dst_data104, sc2mac_wt_dst_data105, sc2mac_wt_dst_data106, sc2mac_wt_dst_data107, sc2mac_wt_dst_data108, sc2mac_wt_dst_data109, sc2mac_wt_dst_data110, sc2mac_wt_dst_data111, sc2mac_wt_dst_data112, sc2mac_wt_dst_data113, sc2mac_wt_dst_data114, sc2mac_wt_dst_data115, sc2mac_wt_dst_data116, sc2mac_wt_dst_data117, sc2mac_wt_dst_data118, sc2mac_wt_dst_data119, sc2mac_wt_dst_data120, sc2mac_wt_dst_data121, sc2mac_wt_dst_data122, sc2mac_wt_dst_data123, sc2mac_wt_dst_data124, sc2mac_wt_dst_data125, sc2mac_wt_dst_data126, sc2mac_wt_dst_data127, sc2mac_wt_dst_sel, sc2mac_dat_dst_pvld, sc2mac_dat_dst_mask, sc2mac_dat_dst_data0, sc2mac_dat_dst_data1, sc2mac_dat_dst_data2, sc2mac_dat_dst_data3, sc2mac_dat_dst_data4, sc2mac_dat_dst_data5, sc2mac_dat_dst_data6, sc2mac_dat_dst_data7, sc2mac_dat_dst_data8, sc2mac_dat_dst_data9, sc2mac_dat_dst_data10, sc2mac_dat_dst_data11, sc2mac_dat_dst_data12, sc2mac_dat_dst_data13, sc2mac_dat_dst_data14, sc2mac_dat_dst_data15, sc2mac_dat_dst_data16, sc2mac_dat_dst_data17, sc2mac_dat_dst_data18, sc2mac_dat_dst_data19, sc2mac_dat_dst_data20, sc2mac_dat_dst_data21, sc2mac_dat_dst_data22, sc2mac_dat_dst_data23, sc2mac_dat_dst_data24, sc2mac_dat_dst_data25, sc2mac_dat_dst_data26, sc2mac_dat_dst_data27, sc2mac_dat_dst_data28, sc2mac_dat_dst_data29, sc2mac_dat_dst_data30, sc2mac_dat_dst_data31, sc2mac_dat_dst_data32, sc2mac_dat_dst_data33, sc2mac_dat_dst_data34, sc2mac_dat_dst_data35, sc2mac_dat_dst_data36, sc2mac_dat_dst_data37, sc2mac_dat_dst_data38, sc2mac_dat_dst_data39, sc2mac_dat_dst_data40, sc2mac_dat_dst_data41, sc2mac_dat_dst_data42, sc2mac_dat_dst_data43, sc2mac_dat_dst_data44, sc2mac_dat_dst_data45, sc2mac_dat_dst_data46, sc2mac_dat_dst_data47, sc2mac_dat_dst_data48, sc2mac_dat_dst_data49, sc2mac_dat_dst_data50, sc2mac_dat_dst_data51, sc2mac_dat_dst_data52, sc2mac_dat_dst_data53, sc2mac_dat_dst_data54, sc2mac_dat_dst_data55, sc2mac_dat_dst_data56, sc2mac_dat_dst_data57, sc2mac_dat_dst_data58, sc2mac_dat_dst_data59, sc2mac_dat_dst_data60, sc2mac_dat_dst_data61, sc2mac_dat_dst_data62, sc2mac_dat_dst_data63, sc2mac_dat_dst_data64, sc2mac_dat_dst_data65, sc2mac_dat_dst_data66, sc2mac_dat_dst_data67, sc2mac_dat_dst_data68, sc2mac_dat_dst_data69, sc2mac_dat_dst_data70, sc2mac_dat_dst_data71, sc2mac_dat_dst_data72, sc2mac_dat_dst_data73, sc2mac_dat_dst_data74, sc2mac_dat_dst_data75, sc2mac_dat_dst_data76, sc2mac_dat_dst_data77, sc2mac_dat_dst_data78, sc2mac_dat_dst_data79, sc2mac_dat_dst_data80, sc2mac_dat_dst_data81, sc2mac_dat_dst_data82, sc2mac_dat_dst_data83, sc2mac_dat_dst_data84, sc2mac_dat_dst_data85, sc2mac_dat_dst_data86, sc2mac_dat_dst_data87, sc2mac_dat_dst_data88, sc2mac_dat_dst_data89, sc2mac_dat_dst_data90, sc2mac_dat_dst_data91, sc2mac_dat_dst_data92, sc2mac_dat_dst_data93, sc2mac_dat_dst_data94, sc2mac_dat_dst_data95, sc2mac_dat_dst_data96, sc2mac_dat_dst_data97, sc2mac_dat_dst_data98, sc2mac_dat_dst_data99, sc2mac_dat_dst_data100, sc2mac_dat_dst_data101, sc2mac_dat_dst_data102, sc2mac_dat_dst_data103, sc2mac_dat_dst_data104, sc2mac_dat_dst_data105, sc2mac_dat_dst_data106, sc2mac_dat_dst_data107, sc2mac_dat_dst_data108, sc2mac_dat_dst_data109, sc2mac_dat_dst_data110, sc2mac_dat_dst_data111, sc2mac_dat_dst_data112, sc2mac_dat_dst_data113, sc2mac_dat_dst_data114, sc2mac_dat_dst_data115, sc2mac_dat_dst_data116, sc2mac_dat_dst_data117, sc2mac_dat_dst_data118, sc2mac_dat_dst_data119, sc2mac_dat_dst_data120, sc2mac_dat_dst_data121, sc2mac_dat_dst_data122, sc2mac_dat_dst_data123, sc2mac_dat_dst_data124, sc2mac_dat_dst_data125, sc2mac_dat_dst_data126, sc2mac_dat_dst_data127, sc2mac_dat_dst_pd);
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:3652" *)
  wire [7:0] _0000_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:6470" *)
  wire [7:0] _0001_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:4652" *)
  wire [7:0] _0002_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:7470" *)
  wire [7:0] _0003_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:4662" *)
  wire [7:0] _0004_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:7480" *)
  wire [7:0] _0005_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:4672" *)
  wire [7:0] _0006_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:7490" *)
  wire [7:0] _0007_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:4682" *)
  wire [7:0] _0008_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:7500" *)
  wire [7:0] _0009_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:4692" *)
  wire [7:0] _0010_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:7510" *)
  wire [7:0] _0011_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:4702" *)
  wire [7:0] _0012_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:7520" *)
  wire [7:0] _0013_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:4712" *)
  wire [7:0] _0014_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:7530" *)
  wire [7:0] _0015_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:4722" *)
  wire [7:0] _0016_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:7540" *)
  wire [7:0] _0017_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:4732" *)
  wire [7:0] _0018_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:7550" *)
  wire [7:0] _0019_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:4742" *)
  wire [7:0] _0020_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:7560" *)
  wire [7:0] _0021_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:3752" *)
  wire [7:0] _0022_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:6570" *)
  wire [7:0] _0023_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:4752" *)
  wire [7:0] _0024_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:7570" *)
  wire [7:0] _0025_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:4762" *)
  wire [7:0] _0026_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:7580" *)
  wire [7:0] _0027_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:4772" *)
  wire [7:0] _0028_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:7590" *)
  wire [7:0] _0029_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:4782" *)
  wire [7:0] _0030_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:7600" *)
  wire [7:0] _0031_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:4792" *)
  wire [7:0] _0032_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:7610" *)
  wire [7:0] _0033_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:4802" *)
  wire [7:0] _0034_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:7620" *)
  wire [7:0] _0035_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:4812" *)
  wire [7:0] _0036_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:7630" *)
  wire [7:0] _0037_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:4822" *)
  wire [7:0] _0038_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:7640" *)
  wire [7:0] _0039_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:4832" *)
  wire [7:0] _0040_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:7650" *)
  wire [7:0] _0041_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:4842" *)
  wire [7:0] _0042_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:7660" *)
  wire [7:0] _0043_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:3762" *)
  wire [7:0] _0044_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:6580" *)
  wire [7:0] _0045_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:4852" *)
  wire [7:0] _0046_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:7670" *)
  wire [7:0] _0047_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:4862" *)
  wire [7:0] _0048_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:7680" *)
  wire [7:0] _0049_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:4872" *)
  wire [7:0] _0050_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:7690" *)
  wire [7:0] _0051_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:4882" *)
  wire [7:0] _0052_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:7700" *)
  wire [7:0] _0053_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:4892" *)
  wire [7:0] _0054_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:7710" *)
  wire [7:0] _0055_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:4902" *)
  wire [7:0] _0056_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:7720" *)
  wire [7:0] _0057_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:4912" *)
  wire [7:0] _0058_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:7730" *)
  wire [7:0] _0059_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:4922" *)
  wire [7:0] _0060_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:7740" *)
  wire [7:0] _0061_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:3772" *)
  wire [7:0] _0062_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:6590" *)
  wire [7:0] _0063_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:3782" *)
  wire [7:0] _0064_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:6600" *)
  wire [7:0] _0065_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:3792" *)
  wire [7:0] _0066_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:6610" *)
  wire [7:0] _0067_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:3802" *)
  wire [7:0] _0068_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:6620" *)
  wire [7:0] _0069_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:3812" *)
  wire [7:0] _0070_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:6630" *)
  wire [7:0] _0071_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:3822" *)
  wire [7:0] _0072_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:6640" *)
  wire [7:0] _0073_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:3832" *)
  wire [7:0] _0074_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:6650" *)
  wire [7:0] _0075_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:3842" *)
  wire [7:0] _0076_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:6660" *)
  wire [7:0] _0077_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:3662" *)
  wire [7:0] _0078_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:6480" *)
  wire [7:0] _0079_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:3852" *)
  wire [7:0] _0080_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:6670" *)
  wire [7:0] _0081_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:3862" *)
  wire [7:0] _0082_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:6680" *)
  wire [7:0] _0083_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:3872" *)
  wire [7:0] _0084_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:6690" *)
  wire [7:0] _0085_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:3882" *)
  wire [7:0] _0086_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:6700" *)
  wire [7:0] _0087_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:3892" *)
  wire [7:0] _0088_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:6710" *)
  wire [7:0] _0089_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:3902" *)
  wire [7:0] _0090_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:6720" *)
  wire [7:0] _0091_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:3912" *)
  wire [7:0] _0092_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:6730" *)
  wire [7:0] _0093_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:3922" *)
  wire [7:0] _0094_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:6740" *)
  wire [7:0] _0095_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:3932" *)
  wire [7:0] _0096_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:6750" *)
  wire [7:0] _0097_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:3942" *)
  wire [7:0] _0098_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:6760" *)
  wire [7:0] _0099_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:3672" *)
  wire [7:0] _0100_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:6490" *)
  wire [7:0] _0101_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:3952" *)
  wire [7:0] _0102_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:6770" *)
  wire [7:0] _0103_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:3962" *)
  wire [7:0] _0104_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:6780" *)
  wire [7:0] _0105_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:3972" *)
  wire [7:0] _0106_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:6790" *)
  wire [7:0] _0107_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:3982" *)
  wire [7:0] _0108_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:6800" *)
  wire [7:0] _0109_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:3992" *)
  wire [7:0] _0110_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:6810" *)
  wire [7:0] _0111_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:4002" *)
  wire [7:0] _0112_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:6820" *)
  wire [7:0] _0113_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:4012" *)
  wire [7:0] _0114_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:6830" *)
  wire [7:0] _0115_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:4022" *)
  wire [7:0] _0116_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:6840" *)
  wire [7:0] _0117_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:4032" *)
  wire [7:0] _0118_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:6850" *)
  wire [7:0] _0119_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:4042" *)
  wire [7:0] _0120_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:6860" *)
  wire [7:0] _0121_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:3682" *)
  wire [7:0] _0122_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:6500" *)
  wire [7:0] _0123_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:4052" *)
  wire [7:0] _0124_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:6870" *)
  wire [7:0] _0125_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:4062" *)
  wire [7:0] _0126_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:6880" *)
  wire [7:0] _0127_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:4072" *)
  wire [7:0] _0128_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:6890" *)
  wire [7:0] _0129_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:4082" *)
  wire [7:0] _0130_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:6900" *)
  wire [7:0] _0131_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:4092" *)
  wire [7:0] _0132_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:6910" *)
  wire [7:0] _0133_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:4102" *)
  wire [7:0] _0134_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:6920" *)
  wire [7:0] _0135_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:4112" *)
  wire [7:0] _0136_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:6930" *)
  wire [7:0] _0137_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:4122" *)
  wire [7:0] _0138_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:6940" *)
  wire [7:0] _0139_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:4132" *)
  wire [7:0] _0140_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:6950" *)
  wire [7:0] _0141_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:4142" *)
  wire [7:0] _0142_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:6960" *)
  wire [7:0] _0143_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:3692" *)
  wire [7:0] _0144_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:6510" *)
  wire [7:0] _0145_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:4152" *)
  wire [7:0] _0146_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:6970" *)
  wire [7:0] _0147_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:4162" *)
  wire [7:0] _0148_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:6980" *)
  wire [7:0] _0149_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:4172" *)
  wire [7:0] _0150_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:6990" *)
  wire [7:0] _0151_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:4182" *)
  wire [7:0] _0152_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:7000" *)
  wire [7:0] _0153_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:4192" *)
  wire [7:0] _0154_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:7010" *)
  wire [7:0] _0155_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:4202" *)
  wire [7:0] _0156_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:7020" *)
  wire [7:0] _0157_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:4212" *)
  wire [7:0] _0158_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:7030" *)
  wire [7:0] _0159_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:4222" *)
  wire [7:0] _0160_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:7040" *)
  wire [7:0] _0161_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:4232" *)
  wire [7:0] _0162_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:7050" *)
  wire [7:0] _0163_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:4242" *)
  wire [7:0] _0164_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:7060" *)
  wire [7:0] _0165_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:3702" *)
  wire [7:0] _0166_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:6520" *)
  wire [7:0] _0167_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:4252" *)
  wire [7:0] _0168_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:7070" *)
  wire [7:0] _0169_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:4262" *)
  wire [7:0] _0170_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:7080" *)
  wire [7:0] _0171_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:4272" *)
  wire [7:0] _0172_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:7090" *)
  wire [7:0] _0173_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:4282" *)
  wire [7:0] _0174_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:7100" *)
  wire [7:0] _0175_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:4292" *)
  wire [7:0] _0176_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:7110" *)
  wire [7:0] _0177_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:4302" *)
  wire [7:0] _0178_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:7120" *)
  wire [7:0] _0179_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:4312" *)
  wire [7:0] _0180_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:7130" *)
  wire [7:0] _0181_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:4322" *)
  wire [7:0] _0182_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:7140" *)
  wire [7:0] _0183_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:4332" *)
  wire [7:0] _0184_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:7150" *)
  wire [7:0] _0185_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:4342" *)
  wire [7:0] _0186_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:7160" *)
  wire [7:0] _0187_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:3712" *)
  wire [7:0] _0188_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:6530" *)
  wire [7:0] _0189_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:4352" *)
  wire [7:0] _0190_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:7170" *)
  wire [7:0] _0191_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:4362" *)
  wire [7:0] _0192_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:7180" *)
  wire [7:0] _0193_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:4372" *)
  wire [7:0] _0194_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:7190" *)
  wire [7:0] _0195_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:4382" *)
  wire [7:0] _0196_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:7200" *)
  wire [7:0] _0197_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:4392" *)
  wire [7:0] _0198_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:7210" *)
  wire [7:0] _0199_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:4402" *)
  wire [7:0] _0200_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:7220" *)
  wire [7:0] _0201_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:4412" *)
  wire [7:0] _0202_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:7230" *)
  wire [7:0] _0203_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:4422" *)
  wire [7:0] _0204_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:7240" *)
  wire [7:0] _0205_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:4432" *)
  wire [7:0] _0206_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:7250" *)
  wire [7:0] _0207_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:4442" *)
  wire [7:0] _0208_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:7260" *)
  wire [7:0] _0209_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:3722" *)
  wire [7:0] _0210_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:6540" *)
  wire [7:0] _0211_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:4452" *)
  wire [7:0] _0212_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:7270" *)
  wire [7:0] _0213_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:4462" *)
  wire [7:0] _0214_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:7280" *)
  wire [7:0] _0215_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:4472" *)
  wire [7:0] _0216_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:7290" *)
  wire [7:0] _0217_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:4482" *)
  wire [7:0] _0218_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:7300" *)
  wire [7:0] _0219_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:4492" *)
  wire [7:0] _0220_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:7310" *)
  wire [7:0] _0221_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:4502" *)
  wire [7:0] _0222_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:7320" *)
  wire [7:0] _0223_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:4512" *)
  wire [7:0] _0224_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:7330" *)
  wire [7:0] _0225_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:4522" *)
  wire [7:0] _0226_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:7340" *)
  wire [7:0] _0227_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:4532" *)
  wire [7:0] _0228_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:7350" *)
  wire [7:0] _0229_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:4542" *)
  wire [7:0] _0230_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:7360" *)
  wire [7:0] _0231_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:3732" *)
  wire [7:0] _0232_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:6550" *)
  wire [7:0] _0233_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:4552" *)
  wire [7:0] _0234_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:7370" *)
  wire [7:0] _0235_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:4562" *)
  wire [7:0] _0236_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:7380" *)
  wire [7:0] _0237_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:4572" *)
  wire [7:0] _0238_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:7390" *)
  wire [7:0] _0239_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:4582" *)
  wire [7:0] _0240_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:7400" *)
  wire [7:0] _0241_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:4592" *)
  wire [7:0] _0242_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:7410" *)
  wire [7:0] _0243_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:4602" *)
  wire [7:0] _0244_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:7420" *)
  wire [7:0] _0245_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:4612" *)
  wire [7:0] _0246_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:7430" *)
  wire [7:0] _0247_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:4622" *)
  wire [7:0] _0248_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:7440" *)
  wire [7:0] _0249_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:4632" *)
  wire [7:0] _0250_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:7450" *)
  wire [7:0] _0251_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:4642" *)
  wire [7:0] _0252_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:7460" *)
  wire [7:0] _0253_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:3742" *)
  wire [7:0] _0254_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:6560" *)
  wire [7:0] _0255_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:3591" *)
  wire [127:0] _0256_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:6409" *)
  wire [127:0] _0257_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:3530" *)
  wire [8:0] _0258_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:6348" *)
  wire [8:0] _0259_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:2243" *)
  wire [7:0] _0260_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:5061" *)
  wire [7:0] _0261_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:3243" *)
  wire [7:0] _0262_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:6061" *)
  wire [7:0] _0263_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:3253" *)
  wire [7:0] _0264_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:6071" *)
  wire [7:0] _0265_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:3263" *)
  wire [7:0] _0266_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:6081" *)
  wire [7:0] _0267_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:3273" *)
  wire [7:0] _0268_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:6091" *)
  wire [7:0] _0269_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:3283" *)
  wire [7:0] _0270_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:6101" *)
  wire [7:0] _0271_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:3293" *)
  wire [7:0] _0272_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:6111" *)
  wire [7:0] _0273_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:3303" *)
  wire [7:0] _0274_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:6121" *)
  wire [7:0] _0275_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:3313" *)
  wire [7:0] _0276_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:6131" *)
  wire [7:0] _0277_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:3323" *)
  wire [7:0] _0278_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:6141" *)
  wire [7:0] _0279_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:3333" *)
  wire [7:0] _0280_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:6151" *)
  wire [7:0] _0281_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:2343" *)
  wire [7:0] _0282_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:5161" *)
  wire [7:0] _0283_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:3343" *)
  wire [7:0] _0284_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:6161" *)
  wire [7:0] _0285_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:3353" *)
  wire [7:0] _0286_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:6171" *)
  wire [7:0] _0287_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:3363" *)
  wire [7:0] _0288_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:6181" *)
  wire [7:0] _0289_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:3373" *)
  wire [7:0] _0290_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:6191" *)
  wire [7:0] _0291_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:3383" *)
  wire [7:0] _0292_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:6201" *)
  wire [7:0] _0293_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:3393" *)
  wire [7:0] _0294_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:6211" *)
  wire [7:0] _0295_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:3403" *)
  wire [7:0] _0296_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:6221" *)
  wire [7:0] _0297_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:3413" *)
  wire [7:0] _0298_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:6231" *)
  wire [7:0] _0299_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:3423" *)
  wire [7:0] _0300_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:6241" *)
  wire [7:0] _0301_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:3433" *)
  wire [7:0] _0302_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:6251" *)
  wire [7:0] _0303_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:2353" *)
  wire [7:0] _0304_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:5171" *)
  wire [7:0] _0305_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:3443" *)
  wire [7:0] _0306_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:6261" *)
  wire [7:0] _0307_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:3453" *)
  wire [7:0] _0308_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:6271" *)
  wire [7:0] _0309_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:3463" *)
  wire [7:0] _0310_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:6281" *)
  wire [7:0] _0311_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:3473" *)
  wire [7:0] _0312_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:6291" *)
  wire [7:0] _0313_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:3483" *)
  wire [7:0] _0314_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:6301" *)
  wire [7:0] _0315_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:3493" *)
  wire [7:0] _0316_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:6311" *)
  wire [7:0] _0317_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:3503" *)
  wire [7:0] _0318_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:6321" *)
  wire [7:0] _0319_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:3513" *)
  wire [7:0] _0320_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:6331" *)
  wire [7:0] _0321_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:2363" *)
  wire [7:0] _0322_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:5181" *)
  wire [7:0] _0323_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:2373" *)
  wire [7:0] _0324_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:5191" *)
  wire [7:0] _0325_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:2383" *)
  wire [7:0] _0326_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:5201" *)
  wire [7:0] _0327_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:2393" *)
  wire [7:0] _0328_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:5211" *)
  wire [7:0] _0329_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:2403" *)
  wire [7:0] _0330_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:5221" *)
  wire [7:0] _0331_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:2413" *)
  wire [7:0] _0332_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:5231" *)
  wire [7:0] _0333_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:2423" *)
  wire [7:0] _0334_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:5241" *)
  wire [7:0] _0335_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:2433" *)
  wire [7:0] _0336_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:5251" *)
  wire [7:0] _0337_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:2253" *)
  wire [7:0] _0338_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:5071" *)
  wire [7:0] _0339_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:2443" *)
  wire [7:0] _0340_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:5261" *)
  wire [7:0] _0341_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:2453" *)
  wire [7:0] _0342_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:5271" *)
  wire [7:0] _0343_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:2463" *)
  wire [7:0] _0344_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:5281" *)
  wire [7:0] _0345_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:2473" *)
  wire [7:0] _0346_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:5291" *)
  wire [7:0] _0347_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:2483" *)
  wire [7:0] _0348_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:5301" *)
  wire [7:0] _0349_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:2493" *)
  wire [7:0] _0350_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:5311" *)
  wire [7:0] _0351_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:2503" *)
  wire [7:0] _0352_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:5321" *)
  wire [7:0] _0353_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:2513" *)
  wire [7:0] _0354_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:5331" *)
  wire [7:0] _0355_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:2523" *)
  wire [7:0] _0356_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:5341" *)
  wire [7:0] _0357_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:2533" *)
  wire [7:0] _0358_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:5351" *)
  wire [7:0] _0359_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:2263" *)
  wire [7:0] _0360_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:5081" *)
  wire [7:0] _0361_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:2543" *)
  wire [7:0] _0362_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:5361" *)
  wire [7:0] _0363_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:2553" *)
  wire [7:0] _0364_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:5371" *)
  wire [7:0] _0365_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:2563" *)
  wire [7:0] _0366_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:5381" *)
  wire [7:0] _0367_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:2573" *)
  wire [7:0] _0368_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:5391" *)
  wire [7:0] _0369_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:2583" *)
  wire [7:0] _0370_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:5401" *)
  wire [7:0] _0371_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:2593" *)
  wire [7:0] _0372_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:5411" *)
  wire [7:0] _0373_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:2603" *)
  wire [7:0] _0374_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:5421" *)
  wire [7:0] _0375_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:2613" *)
  wire [7:0] _0376_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:5431" *)
  wire [7:0] _0377_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:2623" *)
  wire [7:0] _0378_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:5441" *)
  wire [7:0] _0379_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:2633" *)
  wire [7:0] _0380_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:5451" *)
  wire [7:0] _0381_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:2273" *)
  wire [7:0] _0382_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:5091" *)
  wire [7:0] _0383_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:2643" *)
  wire [7:0] _0384_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:5461" *)
  wire [7:0] _0385_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:2653" *)
  wire [7:0] _0386_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:5471" *)
  wire [7:0] _0387_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:2663" *)
  wire [7:0] _0388_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:5481" *)
  wire [7:0] _0389_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:2673" *)
  wire [7:0] _0390_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:5491" *)
  wire [7:0] _0391_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:2683" *)
  wire [7:0] _0392_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:5501" *)
  wire [7:0] _0393_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:2693" *)
  wire [7:0] _0394_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:5511" *)
  wire [7:0] _0395_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:2703" *)
  wire [7:0] _0396_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:5521" *)
  wire [7:0] _0397_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:2713" *)
  wire [7:0] _0398_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:5531" *)
  wire [7:0] _0399_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:2723" *)
  wire [7:0] _0400_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:5541" *)
  wire [7:0] _0401_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:2733" *)
  wire [7:0] _0402_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:5551" *)
  wire [7:0] _0403_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:2283" *)
  wire [7:0] _0404_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:5101" *)
  wire [7:0] _0405_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:2743" *)
  wire [7:0] _0406_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:5561" *)
  wire [7:0] _0407_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:2753" *)
  wire [7:0] _0408_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:5571" *)
  wire [7:0] _0409_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:2763" *)
  wire [7:0] _0410_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:5581" *)
  wire [7:0] _0411_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:2773" *)
  wire [7:0] _0412_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:5591" *)
  wire [7:0] _0413_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:2783" *)
  wire [7:0] _0414_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:5601" *)
  wire [7:0] _0415_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:2793" *)
  wire [7:0] _0416_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:5611" *)
  wire [7:0] _0417_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:2803" *)
  wire [7:0] _0418_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:5621" *)
  wire [7:0] _0419_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:2813" *)
  wire [7:0] _0420_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:5631" *)
  wire [7:0] _0421_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:2823" *)
  wire [7:0] _0422_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:5641" *)
  wire [7:0] _0423_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:2833" *)
  wire [7:0] _0424_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:5651" *)
  wire [7:0] _0425_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:2293" *)
  wire [7:0] _0426_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:5111" *)
  wire [7:0] _0427_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:2843" *)
  wire [7:0] _0428_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:5661" *)
  wire [7:0] _0429_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:2853" *)
  wire [7:0] _0430_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:5671" *)
  wire [7:0] _0431_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:2863" *)
  wire [7:0] _0432_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:5681" *)
  wire [7:0] _0433_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:2873" *)
  wire [7:0] _0434_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:5691" *)
  wire [7:0] _0435_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:2883" *)
  wire [7:0] _0436_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:5701" *)
  wire [7:0] _0437_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:2893" *)
  wire [7:0] _0438_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:5711" *)
  wire [7:0] _0439_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:2903" *)
  wire [7:0] _0440_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:5721" *)
  wire [7:0] _0441_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:2913" *)
  wire [7:0] _0442_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:5731" *)
  wire [7:0] _0443_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:2923" *)
  wire [7:0] _0444_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:5741" *)
  wire [7:0] _0445_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:2933" *)
  wire [7:0] _0446_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:5751" *)
  wire [7:0] _0447_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:2303" *)
  wire [7:0] _0448_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:5121" *)
  wire [7:0] _0449_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:2943" *)
  wire [7:0] _0450_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:5761" *)
  wire [7:0] _0451_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:2953" *)
  wire [7:0] _0452_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:5771" *)
  wire [7:0] _0453_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:2963" *)
  wire [7:0] _0454_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:5781" *)
  wire [7:0] _0455_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:2973" *)
  wire [7:0] _0456_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:5791" *)
  wire [7:0] _0457_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:2983" *)
  wire [7:0] _0458_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:5801" *)
  wire [7:0] _0459_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:2993" *)
  wire [7:0] _0460_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:5811" *)
  wire [7:0] _0461_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:3003" *)
  wire [7:0] _0462_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:5821" *)
  wire [7:0] _0463_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:3013" *)
  wire [7:0] _0464_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:5831" *)
  wire [7:0] _0465_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:3023" *)
  wire [7:0] _0466_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:5841" *)
  wire [7:0] _0467_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:3033" *)
  wire [7:0] _0468_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:5851" *)
  wire [7:0] _0469_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:2313" *)
  wire [7:0] _0470_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:5131" *)
  wire [7:0] _0471_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:3043" *)
  wire [7:0] _0472_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:5861" *)
  wire [7:0] _0473_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:3053" *)
  wire [7:0] _0474_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:5871" *)
  wire [7:0] _0475_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:3063" *)
  wire [7:0] _0476_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:5881" *)
  wire [7:0] _0477_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:3073" *)
  wire [7:0] _0478_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:5891" *)
  wire [7:0] _0479_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:3083" *)
  wire [7:0] _0480_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:5901" *)
  wire [7:0] _0481_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:3093" *)
  wire [7:0] _0482_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:5911" *)
  wire [7:0] _0483_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:3103" *)
  wire [7:0] _0484_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:5921" *)
  wire [7:0] _0485_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:3113" *)
  wire [7:0] _0486_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:5931" *)
  wire [7:0] _0487_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:3123" *)
  wire [7:0] _0488_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:5941" *)
  wire [7:0] _0489_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:3133" *)
  wire [7:0] _0490_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:5951" *)
  wire [7:0] _0491_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:2323" *)
  wire [7:0] _0492_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:5141" *)
  wire [7:0] _0493_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:3143" *)
  wire [7:0] _0494_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:5961" *)
  wire [7:0] _0495_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:3153" *)
  wire [7:0] _0496_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:5971" *)
  wire [7:0] _0497_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:3163" *)
  wire [7:0] _0498_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:5981" *)
  wire [7:0] _0499_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:3173" *)
  wire [7:0] _0500_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:5991" *)
  wire [7:0] _0501_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:3183" *)
  wire [7:0] _0502_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:6001" *)
  wire [7:0] _0503_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:3193" *)
  wire [7:0] _0504_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:6011" *)
  wire [7:0] _0505_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:3203" *)
  wire [7:0] _0506_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:6021" *)
  wire [7:0] _0507_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:3213" *)
  wire [7:0] _0508_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:6031" *)
  wire [7:0] _0509_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:3223" *)
  wire [7:0] _0510_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:6041" *)
  wire [7:0] _0511_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:3233" *)
  wire [7:0] _0512_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:6051" *)
  wire [7:0] _0513_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:2333" *)
  wire [7:0] _0514_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:5151" *)
  wire [7:0] _0515_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:2182" *)
  wire [127:0] _0516_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:5000" *)
  wire [127:0] _0517_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:2121" *)
  wire [7:0] _0518_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:4939" *)
  wire [7:0] _0519_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:2125" *)
  wire _0520_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:3534" *)
  wire _0521_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:4943" *)
  wire _0522_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:6352" *)
  wire _0523_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:540" *)
  input nvdla_core_clk;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:541" *)
  input nvdla_core_rstn;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1066" *)
  wire [7:0] sc2mac_dat_data0_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1328" *)
  reg [7:0] sc2mac_dat_data0_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1329" *)
  reg [7:0] sc2mac_dat_data0_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1067" *)
  wire [7:0] sc2mac_dat_data100_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1330" *)
  reg [7:0] sc2mac_dat_data100_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1331" *)
  reg [7:0] sc2mac_dat_data100_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1068" *)
  wire [7:0] sc2mac_dat_data101_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1332" *)
  reg [7:0] sc2mac_dat_data101_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1333" *)
  reg [7:0] sc2mac_dat_data101_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1069" *)
  wire [7:0] sc2mac_dat_data102_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1334" *)
  reg [7:0] sc2mac_dat_data102_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1335" *)
  reg [7:0] sc2mac_dat_data102_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1070" *)
  wire [7:0] sc2mac_dat_data103_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1336" *)
  reg [7:0] sc2mac_dat_data103_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1337" *)
  reg [7:0] sc2mac_dat_data103_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1071" *)
  wire [7:0] sc2mac_dat_data104_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1338" *)
  reg [7:0] sc2mac_dat_data104_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1339" *)
  reg [7:0] sc2mac_dat_data104_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1072" *)
  wire [7:0] sc2mac_dat_data105_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1340" *)
  reg [7:0] sc2mac_dat_data105_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1341" *)
  reg [7:0] sc2mac_dat_data105_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1073" *)
  wire [7:0] sc2mac_dat_data106_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1342" *)
  reg [7:0] sc2mac_dat_data106_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1343" *)
  reg [7:0] sc2mac_dat_data106_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1074" *)
  wire [7:0] sc2mac_dat_data107_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1344" *)
  reg [7:0] sc2mac_dat_data107_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1345" *)
  reg [7:0] sc2mac_dat_data107_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1075" *)
  wire [7:0] sc2mac_dat_data108_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1346" *)
  reg [7:0] sc2mac_dat_data108_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1347" *)
  reg [7:0] sc2mac_dat_data108_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1076" *)
  wire [7:0] sc2mac_dat_data109_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1348" *)
  reg [7:0] sc2mac_dat_data109_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1349" *)
  reg [7:0] sc2mac_dat_data109_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1077" *)
  wire [7:0] sc2mac_dat_data10_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1350" *)
  reg [7:0] sc2mac_dat_data10_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1351" *)
  reg [7:0] sc2mac_dat_data10_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1078" *)
  wire [7:0] sc2mac_dat_data110_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1352" *)
  reg [7:0] sc2mac_dat_data110_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1353" *)
  reg [7:0] sc2mac_dat_data110_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1079" *)
  wire [7:0] sc2mac_dat_data111_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1354" *)
  reg [7:0] sc2mac_dat_data111_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1355" *)
  reg [7:0] sc2mac_dat_data111_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1080" *)
  wire [7:0] sc2mac_dat_data112_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1356" *)
  reg [7:0] sc2mac_dat_data112_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1357" *)
  reg [7:0] sc2mac_dat_data112_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1081" *)
  wire [7:0] sc2mac_dat_data113_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1358" *)
  reg [7:0] sc2mac_dat_data113_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1359" *)
  reg [7:0] sc2mac_dat_data113_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1082" *)
  wire [7:0] sc2mac_dat_data114_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1360" *)
  reg [7:0] sc2mac_dat_data114_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1361" *)
  reg [7:0] sc2mac_dat_data114_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1083" *)
  wire [7:0] sc2mac_dat_data115_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1362" *)
  reg [7:0] sc2mac_dat_data115_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1363" *)
  reg [7:0] sc2mac_dat_data115_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1084" *)
  wire [7:0] sc2mac_dat_data116_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1364" *)
  reg [7:0] sc2mac_dat_data116_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1365" *)
  reg [7:0] sc2mac_dat_data116_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1085" *)
  wire [7:0] sc2mac_dat_data117_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1366" *)
  reg [7:0] sc2mac_dat_data117_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1367" *)
  reg [7:0] sc2mac_dat_data117_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1086" *)
  wire [7:0] sc2mac_dat_data118_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1368" *)
  reg [7:0] sc2mac_dat_data118_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1369" *)
  reg [7:0] sc2mac_dat_data118_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1087" *)
  wire [7:0] sc2mac_dat_data119_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1370" *)
  reg [7:0] sc2mac_dat_data119_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1371" *)
  reg [7:0] sc2mac_dat_data119_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1088" *)
  wire [7:0] sc2mac_dat_data11_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1372" *)
  reg [7:0] sc2mac_dat_data11_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1373" *)
  reg [7:0] sc2mac_dat_data11_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1089" *)
  wire [7:0] sc2mac_dat_data120_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1374" *)
  reg [7:0] sc2mac_dat_data120_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1375" *)
  reg [7:0] sc2mac_dat_data120_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1090" *)
  wire [7:0] sc2mac_dat_data121_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1376" *)
  reg [7:0] sc2mac_dat_data121_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1377" *)
  reg [7:0] sc2mac_dat_data121_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1091" *)
  wire [7:0] sc2mac_dat_data122_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1378" *)
  reg [7:0] sc2mac_dat_data122_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1379" *)
  reg [7:0] sc2mac_dat_data122_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1092" *)
  wire [7:0] sc2mac_dat_data123_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1380" *)
  reg [7:0] sc2mac_dat_data123_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1381" *)
  reg [7:0] sc2mac_dat_data123_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1093" *)
  wire [7:0] sc2mac_dat_data124_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1382" *)
  reg [7:0] sc2mac_dat_data124_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1383" *)
  reg [7:0] sc2mac_dat_data124_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1094" *)
  wire [7:0] sc2mac_dat_data125_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1384" *)
  reg [7:0] sc2mac_dat_data125_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1385" *)
  reg [7:0] sc2mac_dat_data125_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1095" *)
  wire [7:0] sc2mac_dat_data126_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1386" *)
  reg [7:0] sc2mac_dat_data126_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1387" *)
  reg [7:0] sc2mac_dat_data126_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1096" *)
  wire [7:0] sc2mac_dat_data127_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1388" *)
  reg [7:0] sc2mac_dat_data127_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1389" *)
  reg [7:0] sc2mac_dat_data127_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1097" *)
  wire [7:0] sc2mac_dat_data12_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1390" *)
  reg [7:0] sc2mac_dat_data12_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1391" *)
  reg [7:0] sc2mac_dat_data12_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1098" *)
  wire [7:0] sc2mac_dat_data13_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1392" *)
  reg [7:0] sc2mac_dat_data13_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1393" *)
  reg [7:0] sc2mac_dat_data13_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1099" *)
  wire [7:0] sc2mac_dat_data14_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1394" *)
  reg [7:0] sc2mac_dat_data14_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1395" *)
  reg [7:0] sc2mac_dat_data14_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1100" *)
  wire [7:0] sc2mac_dat_data15_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1396" *)
  reg [7:0] sc2mac_dat_data15_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1397" *)
  reg [7:0] sc2mac_dat_data15_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1101" *)
  wire [7:0] sc2mac_dat_data16_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1398" *)
  reg [7:0] sc2mac_dat_data16_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1399" *)
  reg [7:0] sc2mac_dat_data16_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1102" *)
  wire [7:0] sc2mac_dat_data17_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1400" *)
  reg [7:0] sc2mac_dat_data17_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1401" *)
  reg [7:0] sc2mac_dat_data17_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1103" *)
  wire [7:0] sc2mac_dat_data18_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1402" *)
  reg [7:0] sc2mac_dat_data18_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1403" *)
  reg [7:0] sc2mac_dat_data18_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1104" *)
  wire [7:0] sc2mac_dat_data19_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1404" *)
  reg [7:0] sc2mac_dat_data19_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1405" *)
  reg [7:0] sc2mac_dat_data19_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1105" *)
  wire [7:0] sc2mac_dat_data1_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1406" *)
  reg [7:0] sc2mac_dat_data1_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1407" *)
  reg [7:0] sc2mac_dat_data1_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1106" *)
  wire [7:0] sc2mac_dat_data20_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1408" *)
  reg [7:0] sc2mac_dat_data20_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1409" *)
  reg [7:0] sc2mac_dat_data20_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1107" *)
  wire [7:0] sc2mac_dat_data21_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1410" *)
  reg [7:0] sc2mac_dat_data21_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1411" *)
  reg [7:0] sc2mac_dat_data21_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1108" *)
  wire [7:0] sc2mac_dat_data22_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1412" *)
  reg [7:0] sc2mac_dat_data22_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1413" *)
  reg [7:0] sc2mac_dat_data22_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1109" *)
  wire [7:0] sc2mac_dat_data23_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1414" *)
  reg [7:0] sc2mac_dat_data23_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1415" *)
  reg [7:0] sc2mac_dat_data23_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1110" *)
  wire [7:0] sc2mac_dat_data24_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1416" *)
  reg [7:0] sc2mac_dat_data24_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1417" *)
  reg [7:0] sc2mac_dat_data24_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1111" *)
  wire [7:0] sc2mac_dat_data25_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1418" *)
  reg [7:0] sc2mac_dat_data25_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1419" *)
  reg [7:0] sc2mac_dat_data25_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1112" *)
  wire [7:0] sc2mac_dat_data26_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1420" *)
  reg [7:0] sc2mac_dat_data26_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1421" *)
  reg [7:0] sc2mac_dat_data26_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1113" *)
  wire [7:0] sc2mac_dat_data27_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1422" *)
  reg [7:0] sc2mac_dat_data27_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1423" *)
  reg [7:0] sc2mac_dat_data27_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1114" *)
  wire [7:0] sc2mac_dat_data28_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1424" *)
  reg [7:0] sc2mac_dat_data28_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1425" *)
  reg [7:0] sc2mac_dat_data28_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1115" *)
  wire [7:0] sc2mac_dat_data29_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1426" *)
  reg [7:0] sc2mac_dat_data29_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1427" *)
  reg [7:0] sc2mac_dat_data29_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1116" *)
  wire [7:0] sc2mac_dat_data2_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1428" *)
  reg [7:0] sc2mac_dat_data2_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1429" *)
  reg [7:0] sc2mac_dat_data2_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1117" *)
  wire [7:0] sc2mac_dat_data30_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1430" *)
  reg [7:0] sc2mac_dat_data30_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1431" *)
  reg [7:0] sc2mac_dat_data30_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1118" *)
  wire [7:0] sc2mac_dat_data31_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1432" *)
  reg [7:0] sc2mac_dat_data31_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1433" *)
  reg [7:0] sc2mac_dat_data31_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1119" *)
  wire [7:0] sc2mac_dat_data32_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1434" *)
  reg [7:0] sc2mac_dat_data32_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1435" *)
  reg [7:0] sc2mac_dat_data32_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1120" *)
  wire [7:0] sc2mac_dat_data33_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1436" *)
  reg [7:0] sc2mac_dat_data33_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1437" *)
  reg [7:0] sc2mac_dat_data33_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1121" *)
  wire [7:0] sc2mac_dat_data34_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1438" *)
  reg [7:0] sc2mac_dat_data34_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1439" *)
  reg [7:0] sc2mac_dat_data34_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1122" *)
  wire [7:0] sc2mac_dat_data35_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1440" *)
  reg [7:0] sc2mac_dat_data35_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1441" *)
  reg [7:0] sc2mac_dat_data35_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1123" *)
  wire [7:0] sc2mac_dat_data36_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1442" *)
  reg [7:0] sc2mac_dat_data36_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1443" *)
  reg [7:0] sc2mac_dat_data36_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1124" *)
  wire [7:0] sc2mac_dat_data37_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1444" *)
  reg [7:0] sc2mac_dat_data37_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1445" *)
  reg [7:0] sc2mac_dat_data37_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1125" *)
  wire [7:0] sc2mac_dat_data38_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1446" *)
  reg [7:0] sc2mac_dat_data38_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1447" *)
  reg [7:0] sc2mac_dat_data38_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1126" *)
  wire [7:0] sc2mac_dat_data39_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1448" *)
  reg [7:0] sc2mac_dat_data39_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1449" *)
  reg [7:0] sc2mac_dat_data39_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1127" *)
  wire [7:0] sc2mac_dat_data3_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1450" *)
  reg [7:0] sc2mac_dat_data3_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1451" *)
  reg [7:0] sc2mac_dat_data3_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1128" *)
  wire [7:0] sc2mac_dat_data40_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1452" *)
  reg [7:0] sc2mac_dat_data40_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1453" *)
  reg [7:0] sc2mac_dat_data40_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1129" *)
  wire [7:0] sc2mac_dat_data41_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1454" *)
  reg [7:0] sc2mac_dat_data41_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1455" *)
  reg [7:0] sc2mac_dat_data41_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1130" *)
  wire [7:0] sc2mac_dat_data42_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1456" *)
  reg [7:0] sc2mac_dat_data42_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1457" *)
  reg [7:0] sc2mac_dat_data42_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1131" *)
  wire [7:0] sc2mac_dat_data43_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1458" *)
  reg [7:0] sc2mac_dat_data43_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1459" *)
  reg [7:0] sc2mac_dat_data43_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1132" *)
  wire [7:0] sc2mac_dat_data44_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1460" *)
  reg [7:0] sc2mac_dat_data44_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1461" *)
  reg [7:0] sc2mac_dat_data44_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1133" *)
  wire [7:0] sc2mac_dat_data45_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1462" *)
  reg [7:0] sc2mac_dat_data45_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1463" *)
  reg [7:0] sc2mac_dat_data45_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1134" *)
  wire [7:0] sc2mac_dat_data46_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1464" *)
  reg [7:0] sc2mac_dat_data46_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1465" *)
  reg [7:0] sc2mac_dat_data46_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1135" *)
  wire [7:0] sc2mac_dat_data47_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1466" *)
  reg [7:0] sc2mac_dat_data47_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1467" *)
  reg [7:0] sc2mac_dat_data47_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1136" *)
  wire [7:0] sc2mac_dat_data48_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1468" *)
  reg [7:0] sc2mac_dat_data48_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1469" *)
  reg [7:0] sc2mac_dat_data48_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1137" *)
  wire [7:0] sc2mac_dat_data49_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1470" *)
  reg [7:0] sc2mac_dat_data49_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1471" *)
  reg [7:0] sc2mac_dat_data49_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1138" *)
  wire [7:0] sc2mac_dat_data4_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1472" *)
  reg [7:0] sc2mac_dat_data4_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1473" *)
  reg [7:0] sc2mac_dat_data4_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1139" *)
  wire [7:0] sc2mac_dat_data50_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1474" *)
  reg [7:0] sc2mac_dat_data50_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1475" *)
  reg [7:0] sc2mac_dat_data50_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1140" *)
  wire [7:0] sc2mac_dat_data51_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1476" *)
  reg [7:0] sc2mac_dat_data51_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1477" *)
  reg [7:0] sc2mac_dat_data51_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1141" *)
  wire [7:0] sc2mac_dat_data52_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1478" *)
  reg [7:0] sc2mac_dat_data52_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1479" *)
  reg [7:0] sc2mac_dat_data52_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1142" *)
  wire [7:0] sc2mac_dat_data53_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1480" *)
  reg [7:0] sc2mac_dat_data53_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1481" *)
  reg [7:0] sc2mac_dat_data53_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1143" *)
  wire [7:0] sc2mac_dat_data54_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1482" *)
  reg [7:0] sc2mac_dat_data54_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1483" *)
  reg [7:0] sc2mac_dat_data54_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1144" *)
  wire [7:0] sc2mac_dat_data55_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1484" *)
  reg [7:0] sc2mac_dat_data55_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1485" *)
  reg [7:0] sc2mac_dat_data55_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1145" *)
  wire [7:0] sc2mac_dat_data56_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1486" *)
  reg [7:0] sc2mac_dat_data56_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1487" *)
  reg [7:0] sc2mac_dat_data56_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1146" *)
  wire [7:0] sc2mac_dat_data57_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1488" *)
  reg [7:0] sc2mac_dat_data57_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1489" *)
  reg [7:0] sc2mac_dat_data57_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1147" *)
  wire [7:0] sc2mac_dat_data58_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1490" *)
  reg [7:0] sc2mac_dat_data58_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1491" *)
  reg [7:0] sc2mac_dat_data58_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1148" *)
  wire [7:0] sc2mac_dat_data59_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1492" *)
  reg [7:0] sc2mac_dat_data59_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1493" *)
  reg [7:0] sc2mac_dat_data59_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1149" *)
  wire [7:0] sc2mac_dat_data5_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1494" *)
  reg [7:0] sc2mac_dat_data5_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1495" *)
  reg [7:0] sc2mac_dat_data5_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1150" *)
  wire [7:0] sc2mac_dat_data60_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1496" *)
  reg [7:0] sc2mac_dat_data60_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1497" *)
  reg [7:0] sc2mac_dat_data60_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1151" *)
  wire [7:0] sc2mac_dat_data61_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1498" *)
  reg [7:0] sc2mac_dat_data61_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1499" *)
  reg [7:0] sc2mac_dat_data61_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1152" *)
  wire [7:0] sc2mac_dat_data62_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1500" *)
  reg [7:0] sc2mac_dat_data62_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1501" *)
  reg [7:0] sc2mac_dat_data62_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1153" *)
  wire [7:0] sc2mac_dat_data63_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1502" *)
  reg [7:0] sc2mac_dat_data63_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1503" *)
  reg [7:0] sc2mac_dat_data63_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1154" *)
  wire [7:0] sc2mac_dat_data64_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1504" *)
  reg [7:0] sc2mac_dat_data64_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1505" *)
  reg [7:0] sc2mac_dat_data64_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1155" *)
  wire [7:0] sc2mac_dat_data65_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1506" *)
  reg [7:0] sc2mac_dat_data65_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1507" *)
  reg [7:0] sc2mac_dat_data65_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1156" *)
  wire [7:0] sc2mac_dat_data66_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1508" *)
  reg [7:0] sc2mac_dat_data66_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1509" *)
  reg [7:0] sc2mac_dat_data66_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1157" *)
  wire [7:0] sc2mac_dat_data67_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1510" *)
  reg [7:0] sc2mac_dat_data67_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1511" *)
  reg [7:0] sc2mac_dat_data67_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1158" *)
  wire [7:0] sc2mac_dat_data68_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1512" *)
  reg [7:0] sc2mac_dat_data68_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1513" *)
  reg [7:0] sc2mac_dat_data68_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1159" *)
  wire [7:0] sc2mac_dat_data69_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1514" *)
  reg [7:0] sc2mac_dat_data69_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1515" *)
  reg [7:0] sc2mac_dat_data69_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1160" *)
  wire [7:0] sc2mac_dat_data6_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1516" *)
  reg [7:0] sc2mac_dat_data6_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1517" *)
  reg [7:0] sc2mac_dat_data6_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1161" *)
  wire [7:0] sc2mac_dat_data70_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1518" *)
  reg [7:0] sc2mac_dat_data70_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1519" *)
  reg [7:0] sc2mac_dat_data70_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1162" *)
  wire [7:0] sc2mac_dat_data71_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1520" *)
  reg [7:0] sc2mac_dat_data71_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1521" *)
  reg [7:0] sc2mac_dat_data71_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1163" *)
  wire [7:0] sc2mac_dat_data72_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1522" *)
  reg [7:0] sc2mac_dat_data72_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1523" *)
  reg [7:0] sc2mac_dat_data72_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1164" *)
  wire [7:0] sc2mac_dat_data73_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1524" *)
  reg [7:0] sc2mac_dat_data73_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1525" *)
  reg [7:0] sc2mac_dat_data73_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1165" *)
  wire [7:0] sc2mac_dat_data74_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1526" *)
  reg [7:0] sc2mac_dat_data74_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1527" *)
  reg [7:0] sc2mac_dat_data74_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1166" *)
  wire [7:0] sc2mac_dat_data75_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1528" *)
  reg [7:0] sc2mac_dat_data75_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1529" *)
  reg [7:0] sc2mac_dat_data75_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1167" *)
  wire [7:0] sc2mac_dat_data76_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1530" *)
  reg [7:0] sc2mac_dat_data76_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1531" *)
  reg [7:0] sc2mac_dat_data76_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1168" *)
  wire [7:0] sc2mac_dat_data77_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1532" *)
  reg [7:0] sc2mac_dat_data77_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1533" *)
  reg [7:0] sc2mac_dat_data77_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1169" *)
  wire [7:0] sc2mac_dat_data78_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1534" *)
  reg [7:0] sc2mac_dat_data78_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1535" *)
  reg [7:0] sc2mac_dat_data78_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1170" *)
  wire [7:0] sc2mac_dat_data79_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1536" *)
  reg [7:0] sc2mac_dat_data79_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1537" *)
  reg [7:0] sc2mac_dat_data79_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1171" *)
  wire [7:0] sc2mac_dat_data7_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1538" *)
  reg [7:0] sc2mac_dat_data7_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1539" *)
  reg [7:0] sc2mac_dat_data7_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1172" *)
  wire [7:0] sc2mac_dat_data80_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1540" *)
  reg [7:0] sc2mac_dat_data80_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1541" *)
  reg [7:0] sc2mac_dat_data80_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1173" *)
  wire [7:0] sc2mac_dat_data81_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1542" *)
  reg [7:0] sc2mac_dat_data81_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1543" *)
  reg [7:0] sc2mac_dat_data81_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1174" *)
  wire [7:0] sc2mac_dat_data82_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1544" *)
  reg [7:0] sc2mac_dat_data82_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1545" *)
  reg [7:0] sc2mac_dat_data82_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1175" *)
  wire [7:0] sc2mac_dat_data83_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1546" *)
  reg [7:0] sc2mac_dat_data83_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1547" *)
  reg [7:0] sc2mac_dat_data83_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1176" *)
  wire [7:0] sc2mac_dat_data84_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1548" *)
  reg [7:0] sc2mac_dat_data84_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1549" *)
  reg [7:0] sc2mac_dat_data84_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1177" *)
  wire [7:0] sc2mac_dat_data85_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1550" *)
  reg [7:0] sc2mac_dat_data85_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1551" *)
  reg [7:0] sc2mac_dat_data85_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1178" *)
  wire [7:0] sc2mac_dat_data86_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1552" *)
  reg [7:0] sc2mac_dat_data86_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1553" *)
  reg [7:0] sc2mac_dat_data86_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1179" *)
  wire [7:0] sc2mac_dat_data87_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1554" *)
  reg [7:0] sc2mac_dat_data87_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1555" *)
  reg [7:0] sc2mac_dat_data87_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1180" *)
  wire [7:0] sc2mac_dat_data88_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1556" *)
  reg [7:0] sc2mac_dat_data88_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1557" *)
  reg [7:0] sc2mac_dat_data88_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1181" *)
  wire [7:0] sc2mac_dat_data89_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1558" *)
  reg [7:0] sc2mac_dat_data89_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1559" *)
  reg [7:0] sc2mac_dat_data89_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1182" *)
  wire [7:0] sc2mac_dat_data8_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1560" *)
  reg [7:0] sc2mac_dat_data8_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1561" *)
  reg [7:0] sc2mac_dat_data8_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1183" *)
  wire [7:0] sc2mac_dat_data90_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1562" *)
  reg [7:0] sc2mac_dat_data90_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1563" *)
  reg [7:0] sc2mac_dat_data90_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1184" *)
  wire [7:0] sc2mac_dat_data91_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1564" *)
  reg [7:0] sc2mac_dat_data91_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1565" *)
  reg [7:0] sc2mac_dat_data91_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1185" *)
  wire [7:0] sc2mac_dat_data92_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1566" *)
  reg [7:0] sc2mac_dat_data92_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1567" *)
  reg [7:0] sc2mac_dat_data92_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1186" *)
  wire [7:0] sc2mac_dat_data93_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1568" *)
  reg [7:0] sc2mac_dat_data93_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1569" *)
  reg [7:0] sc2mac_dat_data93_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1187" *)
  wire [7:0] sc2mac_dat_data94_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1570" *)
  reg [7:0] sc2mac_dat_data94_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1571" *)
  reg [7:0] sc2mac_dat_data94_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1188" *)
  wire [7:0] sc2mac_dat_data95_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1572" *)
  reg [7:0] sc2mac_dat_data95_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1573" *)
  reg [7:0] sc2mac_dat_data95_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1189" *)
  wire [7:0] sc2mac_dat_data96_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1574" *)
  reg [7:0] sc2mac_dat_data96_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1575" *)
  reg [7:0] sc2mac_dat_data96_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1190" *)
  wire [7:0] sc2mac_dat_data97_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1576" *)
  reg [7:0] sc2mac_dat_data97_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1577" *)
  reg [7:0] sc2mac_dat_data97_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1191" *)
  wire [7:0] sc2mac_dat_data98_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1578" *)
  reg [7:0] sc2mac_dat_data98_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1579" *)
  reg [7:0] sc2mac_dat_data98_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1192" *)
  wire [7:0] sc2mac_dat_data99_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1580" *)
  reg [7:0] sc2mac_dat_data99_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1581" *)
  reg [7:0] sc2mac_dat_data99_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1193" *)
  wire [7:0] sc2mac_dat_data9_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1582" *)
  reg [7:0] sc2mac_dat_data9_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1583" *)
  reg [7:0] sc2mac_dat_data9_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:937" *)
  output [7:0] sc2mac_dat_dst_data0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:938" *)
  output [7:0] sc2mac_dat_dst_data1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:947" *)
  output [7:0] sc2mac_dat_dst_data10;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1037" *)
  output [7:0] sc2mac_dat_dst_data100;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1038" *)
  output [7:0] sc2mac_dat_dst_data101;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1039" *)
  output [7:0] sc2mac_dat_dst_data102;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1040" *)
  output [7:0] sc2mac_dat_dst_data103;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1041" *)
  output [7:0] sc2mac_dat_dst_data104;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1042" *)
  output [7:0] sc2mac_dat_dst_data105;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1043" *)
  output [7:0] sc2mac_dat_dst_data106;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1044" *)
  output [7:0] sc2mac_dat_dst_data107;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1045" *)
  output [7:0] sc2mac_dat_dst_data108;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1046" *)
  output [7:0] sc2mac_dat_dst_data109;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:948" *)
  output [7:0] sc2mac_dat_dst_data11;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1047" *)
  output [7:0] sc2mac_dat_dst_data110;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1048" *)
  output [7:0] sc2mac_dat_dst_data111;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1049" *)
  output [7:0] sc2mac_dat_dst_data112;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1050" *)
  output [7:0] sc2mac_dat_dst_data113;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1051" *)
  output [7:0] sc2mac_dat_dst_data114;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1052" *)
  output [7:0] sc2mac_dat_dst_data115;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1053" *)
  output [7:0] sc2mac_dat_dst_data116;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1054" *)
  output [7:0] sc2mac_dat_dst_data117;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1055" *)
  output [7:0] sc2mac_dat_dst_data118;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1056" *)
  output [7:0] sc2mac_dat_dst_data119;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:949" *)
  output [7:0] sc2mac_dat_dst_data12;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1057" *)
  output [7:0] sc2mac_dat_dst_data120;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1058" *)
  output [7:0] sc2mac_dat_dst_data121;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1059" *)
  output [7:0] sc2mac_dat_dst_data122;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1060" *)
  output [7:0] sc2mac_dat_dst_data123;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1061" *)
  output [7:0] sc2mac_dat_dst_data124;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1062" *)
  output [7:0] sc2mac_dat_dst_data125;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1063" *)
  output [7:0] sc2mac_dat_dst_data126;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1064" *)
  output [7:0] sc2mac_dat_dst_data127;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:950" *)
  output [7:0] sc2mac_dat_dst_data13;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:951" *)
  output [7:0] sc2mac_dat_dst_data14;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:952" *)
  output [7:0] sc2mac_dat_dst_data15;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:953" *)
  output [7:0] sc2mac_dat_dst_data16;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:954" *)
  output [7:0] sc2mac_dat_dst_data17;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:955" *)
  output [7:0] sc2mac_dat_dst_data18;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:956" *)
  output [7:0] sc2mac_dat_dst_data19;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:939" *)
  output [7:0] sc2mac_dat_dst_data2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:957" *)
  output [7:0] sc2mac_dat_dst_data20;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:958" *)
  output [7:0] sc2mac_dat_dst_data21;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:959" *)
  output [7:0] sc2mac_dat_dst_data22;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:960" *)
  output [7:0] sc2mac_dat_dst_data23;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:961" *)
  output [7:0] sc2mac_dat_dst_data24;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:962" *)
  output [7:0] sc2mac_dat_dst_data25;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:963" *)
  output [7:0] sc2mac_dat_dst_data26;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:964" *)
  output [7:0] sc2mac_dat_dst_data27;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:965" *)
  output [7:0] sc2mac_dat_dst_data28;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:966" *)
  output [7:0] sc2mac_dat_dst_data29;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:940" *)
  output [7:0] sc2mac_dat_dst_data3;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:967" *)
  output [7:0] sc2mac_dat_dst_data30;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:968" *)
  output [7:0] sc2mac_dat_dst_data31;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:969" *)
  output [7:0] sc2mac_dat_dst_data32;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:970" *)
  output [7:0] sc2mac_dat_dst_data33;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:971" *)
  output [7:0] sc2mac_dat_dst_data34;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:972" *)
  output [7:0] sc2mac_dat_dst_data35;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:973" *)
  output [7:0] sc2mac_dat_dst_data36;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:974" *)
  output [7:0] sc2mac_dat_dst_data37;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:975" *)
  output [7:0] sc2mac_dat_dst_data38;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:976" *)
  output [7:0] sc2mac_dat_dst_data39;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:941" *)
  output [7:0] sc2mac_dat_dst_data4;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:977" *)
  output [7:0] sc2mac_dat_dst_data40;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:978" *)
  output [7:0] sc2mac_dat_dst_data41;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:979" *)
  output [7:0] sc2mac_dat_dst_data42;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:980" *)
  output [7:0] sc2mac_dat_dst_data43;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:981" *)
  output [7:0] sc2mac_dat_dst_data44;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:982" *)
  output [7:0] sc2mac_dat_dst_data45;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:983" *)
  output [7:0] sc2mac_dat_dst_data46;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:984" *)
  output [7:0] sc2mac_dat_dst_data47;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:985" *)
  output [7:0] sc2mac_dat_dst_data48;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:986" *)
  output [7:0] sc2mac_dat_dst_data49;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:942" *)
  output [7:0] sc2mac_dat_dst_data5;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:987" *)
  output [7:0] sc2mac_dat_dst_data50;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:988" *)
  output [7:0] sc2mac_dat_dst_data51;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:989" *)
  output [7:0] sc2mac_dat_dst_data52;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:990" *)
  output [7:0] sc2mac_dat_dst_data53;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:991" *)
  output [7:0] sc2mac_dat_dst_data54;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:992" *)
  output [7:0] sc2mac_dat_dst_data55;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:993" *)
  output [7:0] sc2mac_dat_dst_data56;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:994" *)
  output [7:0] sc2mac_dat_dst_data57;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:995" *)
  output [7:0] sc2mac_dat_dst_data58;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:996" *)
  output [7:0] sc2mac_dat_dst_data59;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:943" *)
  output [7:0] sc2mac_dat_dst_data6;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:997" *)
  output [7:0] sc2mac_dat_dst_data60;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:998" *)
  output [7:0] sc2mac_dat_dst_data61;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:999" *)
  output [7:0] sc2mac_dat_dst_data62;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1000" *)
  output [7:0] sc2mac_dat_dst_data63;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1001" *)
  output [7:0] sc2mac_dat_dst_data64;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1002" *)
  output [7:0] sc2mac_dat_dst_data65;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1003" *)
  output [7:0] sc2mac_dat_dst_data66;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1004" *)
  output [7:0] sc2mac_dat_dst_data67;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1005" *)
  output [7:0] sc2mac_dat_dst_data68;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1006" *)
  output [7:0] sc2mac_dat_dst_data69;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:944" *)
  output [7:0] sc2mac_dat_dst_data7;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1007" *)
  output [7:0] sc2mac_dat_dst_data70;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1008" *)
  output [7:0] sc2mac_dat_dst_data71;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1009" *)
  output [7:0] sc2mac_dat_dst_data72;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1010" *)
  output [7:0] sc2mac_dat_dst_data73;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1011" *)
  output [7:0] sc2mac_dat_dst_data74;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1012" *)
  output [7:0] sc2mac_dat_dst_data75;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1013" *)
  output [7:0] sc2mac_dat_dst_data76;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1014" *)
  output [7:0] sc2mac_dat_dst_data77;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1015" *)
  output [7:0] sc2mac_dat_dst_data78;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1016" *)
  output [7:0] sc2mac_dat_dst_data79;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:945" *)
  output [7:0] sc2mac_dat_dst_data8;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1017" *)
  output [7:0] sc2mac_dat_dst_data80;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1018" *)
  output [7:0] sc2mac_dat_dst_data81;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1019" *)
  output [7:0] sc2mac_dat_dst_data82;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1020" *)
  output [7:0] sc2mac_dat_dst_data83;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1021" *)
  output [7:0] sc2mac_dat_dst_data84;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1022" *)
  output [7:0] sc2mac_dat_dst_data85;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1023" *)
  output [7:0] sc2mac_dat_dst_data86;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1024" *)
  output [7:0] sc2mac_dat_dst_data87;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1025" *)
  output [7:0] sc2mac_dat_dst_data88;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1026" *)
  output [7:0] sc2mac_dat_dst_data89;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:946" *)
  output [7:0] sc2mac_dat_dst_data9;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1027" *)
  output [7:0] sc2mac_dat_dst_data90;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1028" *)
  output [7:0] sc2mac_dat_dst_data91;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1029" *)
  output [7:0] sc2mac_dat_dst_data92;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1030" *)
  output [7:0] sc2mac_dat_dst_data93;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1031" *)
  output [7:0] sc2mac_dat_dst_data94;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1032" *)
  output [7:0] sc2mac_dat_dst_data95;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1033" *)
  output [7:0] sc2mac_dat_dst_data96;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1034" *)
  output [7:0] sc2mac_dat_dst_data97;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1035" *)
  output [7:0] sc2mac_dat_dst_data98;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1036" *)
  output [7:0] sc2mac_dat_dst_data99;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:936" *)
  output [127:0] sc2mac_dat_dst_mask;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1065" *)
  output [8:0] sc2mac_dat_dst_pd;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:935" *)
  output sc2mac_dat_dst_pvld;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1194" *)
  wire [127:0] sc2mac_dat_mask_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1584" *)
  reg [127:0] sc2mac_dat_mask_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1585" *)
  reg [127:0] sc2mac_dat_mask_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1195" *)
  wire [8:0] sc2mac_dat_pd_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1586" *)
  reg [8:0] sc2mac_dat_pd_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1587" *)
  reg [8:0] sc2mac_dat_pd_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1196" *)
  wire sc2mac_dat_pvld_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1588" *)
  reg sc2mac_dat_pvld_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1589" *)
  reg sc2mac_dat_pvld_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:675" *)
  input [7:0] sc2mac_dat_src_data0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:676" *)
  input [7:0] sc2mac_dat_src_data1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:685" *)
  input [7:0] sc2mac_dat_src_data10;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:775" *)
  input [7:0] sc2mac_dat_src_data100;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:776" *)
  input [7:0] sc2mac_dat_src_data101;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:777" *)
  input [7:0] sc2mac_dat_src_data102;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:778" *)
  input [7:0] sc2mac_dat_src_data103;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:779" *)
  input [7:0] sc2mac_dat_src_data104;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:780" *)
  input [7:0] sc2mac_dat_src_data105;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:781" *)
  input [7:0] sc2mac_dat_src_data106;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:782" *)
  input [7:0] sc2mac_dat_src_data107;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:783" *)
  input [7:0] sc2mac_dat_src_data108;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:784" *)
  input [7:0] sc2mac_dat_src_data109;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:686" *)
  input [7:0] sc2mac_dat_src_data11;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:785" *)
  input [7:0] sc2mac_dat_src_data110;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:786" *)
  input [7:0] sc2mac_dat_src_data111;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:787" *)
  input [7:0] sc2mac_dat_src_data112;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:788" *)
  input [7:0] sc2mac_dat_src_data113;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:789" *)
  input [7:0] sc2mac_dat_src_data114;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:790" *)
  input [7:0] sc2mac_dat_src_data115;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:791" *)
  input [7:0] sc2mac_dat_src_data116;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:792" *)
  input [7:0] sc2mac_dat_src_data117;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:793" *)
  input [7:0] sc2mac_dat_src_data118;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:794" *)
  input [7:0] sc2mac_dat_src_data119;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:687" *)
  input [7:0] sc2mac_dat_src_data12;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:795" *)
  input [7:0] sc2mac_dat_src_data120;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:796" *)
  input [7:0] sc2mac_dat_src_data121;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:797" *)
  input [7:0] sc2mac_dat_src_data122;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:798" *)
  input [7:0] sc2mac_dat_src_data123;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:799" *)
  input [7:0] sc2mac_dat_src_data124;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:800" *)
  input [7:0] sc2mac_dat_src_data125;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:801" *)
  input [7:0] sc2mac_dat_src_data126;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:802" *)
  input [7:0] sc2mac_dat_src_data127;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:688" *)
  input [7:0] sc2mac_dat_src_data13;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:689" *)
  input [7:0] sc2mac_dat_src_data14;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:690" *)
  input [7:0] sc2mac_dat_src_data15;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:691" *)
  input [7:0] sc2mac_dat_src_data16;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:692" *)
  input [7:0] sc2mac_dat_src_data17;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:693" *)
  input [7:0] sc2mac_dat_src_data18;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:694" *)
  input [7:0] sc2mac_dat_src_data19;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:677" *)
  input [7:0] sc2mac_dat_src_data2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:695" *)
  input [7:0] sc2mac_dat_src_data20;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:696" *)
  input [7:0] sc2mac_dat_src_data21;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:697" *)
  input [7:0] sc2mac_dat_src_data22;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:698" *)
  input [7:0] sc2mac_dat_src_data23;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:699" *)
  input [7:0] sc2mac_dat_src_data24;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:700" *)
  input [7:0] sc2mac_dat_src_data25;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:701" *)
  input [7:0] sc2mac_dat_src_data26;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:702" *)
  input [7:0] sc2mac_dat_src_data27;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:703" *)
  input [7:0] sc2mac_dat_src_data28;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:704" *)
  input [7:0] sc2mac_dat_src_data29;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:678" *)
  input [7:0] sc2mac_dat_src_data3;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:705" *)
  input [7:0] sc2mac_dat_src_data30;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:706" *)
  input [7:0] sc2mac_dat_src_data31;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:707" *)
  input [7:0] sc2mac_dat_src_data32;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:708" *)
  input [7:0] sc2mac_dat_src_data33;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:709" *)
  input [7:0] sc2mac_dat_src_data34;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:710" *)
  input [7:0] sc2mac_dat_src_data35;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:711" *)
  input [7:0] sc2mac_dat_src_data36;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:712" *)
  input [7:0] sc2mac_dat_src_data37;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:713" *)
  input [7:0] sc2mac_dat_src_data38;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:714" *)
  input [7:0] sc2mac_dat_src_data39;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:679" *)
  input [7:0] sc2mac_dat_src_data4;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:715" *)
  input [7:0] sc2mac_dat_src_data40;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:716" *)
  input [7:0] sc2mac_dat_src_data41;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:717" *)
  input [7:0] sc2mac_dat_src_data42;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:718" *)
  input [7:0] sc2mac_dat_src_data43;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:719" *)
  input [7:0] sc2mac_dat_src_data44;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:720" *)
  input [7:0] sc2mac_dat_src_data45;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:721" *)
  input [7:0] sc2mac_dat_src_data46;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:722" *)
  input [7:0] sc2mac_dat_src_data47;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:723" *)
  input [7:0] sc2mac_dat_src_data48;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:724" *)
  input [7:0] sc2mac_dat_src_data49;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:680" *)
  input [7:0] sc2mac_dat_src_data5;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:725" *)
  input [7:0] sc2mac_dat_src_data50;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:726" *)
  input [7:0] sc2mac_dat_src_data51;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:727" *)
  input [7:0] sc2mac_dat_src_data52;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:728" *)
  input [7:0] sc2mac_dat_src_data53;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:729" *)
  input [7:0] sc2mac_dat_src_data54;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:730" *)
  input [7:0] sc2mac_dat_src_data55;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:731" *)
  input [7:0] sc2mac_dat_src_data56;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:732" *)
  input [7:0] sc2mac_dat_src_data57;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:733" *)
  input [7:0] sc2mac_dat_src_data58;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:734" *)
  input [7:0] sc2mac_dat_src_data59;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:681" *)
  input [7:0] sc2mac_dat_src_data6;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:735" *)
  input [7:0] sc2mac_dat_src_data60;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:736" *)
  input [7:0] sc2mac_dat_src_data61;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:737" *)
  input [7:0] sc2mac_dat_src_data62;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:738" *)
  input [7:0] sc2mac_dat_src_data63;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:739" *)
  input [7:0] sc2mac_dat_src_data64;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:740" *)
  input [7:0] sc2mac_dat_src_data65;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:741" *)
  input [7:0] sc2mac_dat_src_data66;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:742" *)
  input [7:0] sc2mac_dat_src_data67;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:743" *)
  input [7:0] sc2mac_dat_src_data68;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:744" *)
  input [7:0] sc2mac_dat_src_data69;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:682" *)
  input [7:0] sc2mac_dat_src_data7;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:745" *)
  input [7:0] sc2mac_dat_src_data70;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:746" *)
  input [7:0] sc2mac_dat_src_data71;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:747" *)
  input [7:0] sc2mac_dat_src_data72;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:748" *)
  input [7:0] sc2mac_dat_src_data73;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:749" *)
  input [7:0] sc2mac_dat_src_data74;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:750" *)
  input [7:0] sc2mac_dat_src_data75;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:751" *)
  input [7:0] sc2mac_dat_src_data76;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:752" *)
  input [7:0] sc2mac_dat_src_data77;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:753" *)
  input [7:0] sc2mac_dat_src_data78;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:754" *)
  input [7:0] sc2mac_dat_src_data79;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:683" *)
  input [7:0] sc2mac_dat_src_data8;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:755" *)
  input [7:0] sc2mac_dat_src_data80;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:756" *)
  input [7:0] sc2mac_dat_src_data81;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:757" *)
  input [7:0] sc2mac_dat_src_data82;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:758" *)
  input [7:0] sc2mac_dat_src_data83;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:759" *)
  input [7:0] sc2mac_dat_src_data84;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:760" *)
  input [7:0] sc2mac_dat_src_data85;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:761" *)
  input [7:0] sc2mac_dat_src_data86;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:762" *)
  input [7:0] sc2mac_dat_src_data87;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:763" *)
  input [7:0] sc2mac_dat_src_data88;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:764" *)
  input [7:0] sc2mac_dat_src_data89;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:684" *)
  input [7:0] sc2mac_dat_src_data9;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:765" *)
  input [7:0] sc2mac_dat_src_data90;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:766" *)
  input [7:0] sc2mac_dat_src_data91;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:767" *)
  input [7:0] sc2mac_dat_src_data92;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:768" *)
  input [7:0] sc2mac_dat_src_data93;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:769" *)
  input [7:0] sc2mac_dat_src_data94;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:770" *)
  input [7:0] sc2mac_dat_src_data95;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:771" *)
  input [7:0] sc2mac_dat_src_data96;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:772" *)
  input [7:0] sc2mac_dat_src_data97;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:773" *)
  input [7:0] sc2mac_dat_src_data98;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:774" *)
  input [7:0] sc2mac_dat_src_data99;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:674" *)
  input [127:0] sc2mac_dat_src_mask;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:803" *)
  input [8:0] sc2mac_dat_src_pd;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:673" *)
  input sc2mac_dat_src_pvld;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1197" *)
  wire [7:0] sc2mac_wt_data0_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1590" *)
  reg [7:0] sc2mac_wt_data0_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1591" *)
  reg [7:0] sc2mac_wt_data0_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1198" *)
  wire [7:0] sc2mac_wt_data100_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1592" *)
  reg [7:0] sc2mac_wt_data100_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1593" *)
  reg [7:0] sc2mac_wt_data100_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1199" *)
  wire [7:0] sc2mac_wt_data101_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1594" *)
  reg [7:0] sc2mac_wt_data101_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1595" *)
  reg [7:0] sc2mac_wt_data101_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1200" *)
  wire [7:0] sc2mac_wt_data102_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1596" *)
  reg [7:0] sc2mac_wt_data102_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1597" *)
  reg [7:0] sc2mac_wt_data102_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1201" *)
  wire [7:0] sc2mac_wt_data103_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1598" *)
  reg [7:0] sc2mac_wt_data103_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1599" *)
  reg [7:0] sc2mac_wt_data103_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1202" *)
  wire [7:0] sc2mac_wt_data104_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1600" *)
  reg [7:0] sc2mac_wt_data104_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1601" *)
  reg [7:0] sc2mac_wt_data104_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1203" *)
  wire [7:0] sc2mac_wt_data105_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1602" *)
  reg [7:0] sc2mac_wt_data105_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1603" *)
  reg [7:0] sc2mac_wt_data105_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1204" *)
  wire [7:0] sc2mac_wt_data106_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1604" *)
  reg [7:0] sc2mac_wt_data106_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1605" *)
  reg [7:0] sc2mac_wt_data106_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1205" *)
  wire [7:0] sc2mac_wt_data107_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1606" *)
  reg [7:0] sc2mac_wt_data107_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1607" *)
  reg [7:0] sc2mac_wt_data107_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1206" *)
  wire [7:0] sc2mac_wt_data108_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1608" *)
  reg [7:0] sc2mac_wt_data108_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1609" *)
  reg [7:0] sc2mac_wt_data108_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1207" *)
  wire [7:0] sc2mac_wt_data109_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1610" *)
  reg [7:0] sc2mac_wt_data109_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1611" *)
  reg [7:0] sc2mac_wt_data109_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1208" *)
  wire [7:0] sc2mac_wt_data10_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1612" *)
  reg [7:0] sc2mac_wt_data10_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1613" *)
  reg [7:0] sc2mac_wt_data10_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1209" *)
  wire [7:0] sc2mac_wt_data110_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1614" *)
  reg [7:0] sc2mac_wt_data110_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1615" *)
  reg [7:0] sc2mac_wt_data110_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1210" *)
  wire [7:0] sc2mac_wt_data111_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1616" *)
  reg [7:0] sc2mac_wt_data111_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1617" *)
  reg [7:0] sc2mac_wt_data111_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1211" *)
  wire [7:0] sc2mac_wt_data112_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1618" *)
  reg [7:0] sc2mac_wt_data112_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1619" *)
  reg [7:0] sc2mac_wt_data112_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1212" *)
  wire [7:0] sc2mac_wt_data113_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1620" *)
  reg [7:0] sc2mac_wt_data113_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1621" *)
  reg [7:0] sc2mac_wt_data113_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1213" *)
  wire [7:0] sc2mac_wt_data114_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1622" *)
  reg [7:0] sc2mac_wt_data114_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1623" *)
  reg [7:0] sc2mac_wt_data114_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1214" *)
  wire [7:0] sc2mac_wt_data115_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1624" *)
  reg [7:0] sc2mac_wt_data115_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1625" *)
  reg [7:0] sc2mac_wt_data115_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1215" *)
  wire [7:0] sc2mac_wt_data116_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1626" *)
  reg [7:0] sc2mac_wt_data116_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1627" *)
  reg [7:0] sc2mac_wt_data116_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1216" *)
  wire [7:0] sc2mac_wt_data117_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1628" *)
  reg [7:0] sc2mac_wt_data117_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1629" *)
  reg [7:0] sc2mac_wt_data117_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1217" *)
  wire [7:0] sc2mac_wt_data118_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1630" *)
  reg [7:0] sc2mac_wt_data118_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1631" *)
  reg [7:0] sc2mac_wt_data118_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1218" *)
  wire [7:0] sc2mac_wt_data119_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1632" *)
  reg [7:0] sc2mac_wt_data119_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1633" *)
  reg [7:0] sc2mac_wt_data119_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1219" *)
  wire [7:0] sc2mac_wt_data11_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1634" *)
  reg [7:0] sc2mac_wt_data11_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1635" *)
  reg [7:0] sc2mac_wt_data11_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1220" *)
  wire [7:0] sc2mac_wt_data120_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1636" *)
  reg [7:0] sc2mac_wt_data120_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1637" *)
  reg [7:0] sc2mac_wt_data120_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1221" *)
  wire [7:0] sc2mac_wt_data121_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1638" *)
  reg [7:0] sc2mac_wt_data121_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1639" *)
  reg [7:0] sc2mac_wt_data121_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1222" *)
  wire [7:0] sc2mac_wt_data122_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1640" *)
  reg [7:0] sc2mac_wt_data122_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1641" *)
  reg [7:0] sc2mac_wt_data122_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1223" *)
  wire [7:0] sc2mac_wt_data123_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1642" *)
  reg [7:0] sc2mac_wt_data123_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1643" *)
  reg [7:0] sc2mac_wt_data123_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1224" *)
  wire [7:0] sc2mac_wt_data124_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1644" *)
  reg [7:0] sc2mac_wt_data124_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1645" *)
  reg [7:0] sc2mac_wt_data124_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1225" *)
  wire [7:0] sc2mac_wt_data125_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1646" *)
  reg [7:0] sc2mac_wt_data125_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1647" *)
  reg [7:0] sc2mac_wt_data125_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1226" *)
  wire [7:0] sc2mac_wt_data126_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1648" *)
  reg [7:0] sc2mac_wt_data126_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1649" *)
  reg [7:0] sc2mac_wt_data126_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1227" *)
  wire [7:0] sc2mac_wt_data127_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1650" *)
  reg [7:0] sc2mac_wt_data127_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1651" *)
  reg [7:0] sc2mac_wt_data127_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1228" *)
  wire [7:0] sc2mac_wt_data12_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1652" *)
  reg [7:0] sc2mac_wt_data12_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1653" *)
  reg [7:0] sc2mac_wt_data12_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1229" *)
  wire [7:0] sc2mac_wt_data13_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1654" *)
  reg [7:0] sc2mac_wt_data13_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1655" *)
  reg [7:0] sc2mac_wt_data13_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1230" *)
  wire [7:0] sc2mac_wt_data14_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1656" *)
  reg [7:0] sc2mac_wt_data14_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1657" *)
  reg [7:0] sc2mac_wt_data14_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1231" *)
  wire [7:0] sc2mac_wt_data15_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1658" *)
  reg [7:0] sc2mac_wt_data15_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1659" *)
  reg [7:0] sc2mac_wt_data15_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1232" *)
  wire [7:0] sc2mac_wt_data16_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1660" *)
  reg [7:0] sc2mac_wt_data16_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1661" *)
  reg [7:0] sc2mac_wt_data16_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1233" *)
  wire [7:0] sc2mac_wt_data17_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1662" *)
  reg [7:0] sc2mac_wt_data17_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1663" *)
  reg [7:0] sc2mac_wt_data17_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1234" *)
  wire [7:0] sc2mac_wt_data18_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1664" *)
  reg [7:0] sc2mac_wt_data18_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1665" *)
  reg [7:0] sc2mac_wt_data18_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1235" *)
  wire [7:0] sc2mac_wt_data19_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1666" *)
  reg [7:0] sc2mac_wt_data19_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1667" *)
  reg [7:0] sc2mac_wt_data19_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1236" *)
  wire [7:0] sc2mac_wt_data1_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1668" *)
  reg [7:0] sc2mac_wt_data1_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1669" *)
  reg [7:0] sc2mac_wt_data1_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1237" *)
  wire [7:0] sc2mac_wt_data20_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1670" *)
  reg [7:0] sc2mac_wt_data20_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1671" *)
  reg [7:0] sc2mac_wt_data20_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1238" *)
  wire [7:0] sc2mac_wt_data21_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1672" *)
  reg [7:0] sc2mac_wt_data21_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1673" *)
  reg [7:0] sc2mac_wt_data21_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1239" *)
  wire [7:0] sc2mac_wt_data22_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1674" *)
  reg [7:0] sc2mac_wt_data22_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1675" *)
  reg [7:0] sc2mac_wt_data22_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1240" *)
  wire [7:0] sc2mac_wt_data23_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1676" *)
  reg [7:0] sc2mac_wt_data23_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1677" *)
  reg [7:0] sc2mac_wt_data23_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1241" *)
  wire [7:0] sc2mac_wt_data24_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1678" *)
  reg [7:0] sc2mac_wt_data24_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1679" *)
  reg [7:0] sc2mac_wt_data24_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1242" *)
  wire [7:0] sc2mac_wt_data25_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1680" *)
  reg [7:0] sc2mac_wt_data25_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1681" *)
  reg [7:0] sc2mac_wt_data25_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1243" *)
  wire [7:0] sc2mac_wt_data26_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1682" *)
  reg [7:0] sc2mac_wt_data26_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1683" *)
  reg [7:0] sc2mac_wt_data26_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1244" *)
  wire [7:0] sc2mac_wt_data27_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1684" *)
  reg [7:0] sc2mac_wt_data27_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1685" *)
  reg [7:0] sc2mac_wt_data27_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1245" *)
  wire [7:0] sc2mac_wt_data28_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1686" *)
  reg [7:0] sc2mac_wt_data28_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1687" *)
  reg [7:0] sc2mac_wt_data28_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1246" *)
  wire [7:0] sc2mac_wt_data29_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1688" *)
  reg [7:0] sc2mac_wt_data29_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1689" *)
  reg [7:0] sc2mac_wt_data29_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1247" *)
  wire [7:0] sc2mac_wt_data2_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1690" *)
  reg [7:0] sc2mac_wt_data2_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1691" *)
  reg [7:0] sc2mac_wt_data2_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1248" *)
  wire [7:0] sc2mac_wt_data30_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1692" *)
  reg [7:0] sc2mac_wt_data30_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1693" *)
  reg [7:0] sc2mac_wt_data30_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1249" *)
  wire [7:0] sc2mac_wt_data31_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1694" *)
  reg [7:0] sc2mac_wt_data31_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1695" *)
  reg [7:0] sc2mac_wt_data31_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1250" *)
  wire [7:0] sc2mac_wt_data32_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1696" *)
  reg [7:0] sc2mac_wt_data32_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1697" *)
  reg [7:0] sc2mac_wt_data32_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1251" *)
  wire [7:0] sc2mac_wt_data33_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1698" *)
  reg [7:0] sc2mac_wt_data33_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1699" *)
  reg [7:0] sc2mac_wt_data33_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1252" *)
  wire [7:0] sc2mac_wt_data34_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1700" *)
  reg [7:0] sc2mac_wt_data34_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1701" *)
  reg [7:0] sc2mac_wt_data34_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1253" *)
  wire [7:0] sc2mac_wt_data35_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1702" *)
  reg [7:0] sc2mac_wt_data35_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1703" *)
  reg [7:0] sc2mac_wt_data35_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1254" *)
  wire [7:0] sc2mac_wt_data36_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1704" *)
  reg [7:0] sc2mac_wt_data36_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1705" *)
  reg [7:0] sc2mac_wt_data36_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1255" *)
  wire [7:0] sc2mac_wt_data37_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1706" *)
  reg [7:0] sc2mac_wt_data37_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1707" *)
  reg [7:0] sc2mac_wt_data37_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1256" *)
  wire [7:0] sc2mac_wt_data38_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1708" *)
  reg [7:0] sc2mac_wt_data38_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1709" *)
  reg [7:0] sc2mac_wt_data38_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1257" *)
  wire [7:0] sc2mac_wt_data39_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1710" *)
  reg [7:0] sc2mac_wt_data39_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1711" *)
  reg [7:0] sc2mac_wt_data39_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1258" *)
  wire [7:0] sc2mac_wt_data3_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1712" *)
  reg [7:0] sc2mac_wt_data3_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1713" *)
  reg [7:0] sc2mac_wt_data3_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1259" *)
  wire [7:0] sc2mac_wt_data40_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1714" *)
  reg [7:0] sc2mac_wt_data40_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1715" *)
  reg [7:0] sc2mac_wt_data40_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1260" *)
  wire [7:0] sc2mac_wt_data41_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1716" *)
  reg [7:0] sc2mac_wt_data41_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1717" *)
  reg [7:0] sc2mac_wt_data41_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1261" *)
  wire [7:0] sc2mac_wt_data42_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1718" *)
  reg [7:0] sc2mac_wt_data42_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1719" *)
  reg [7:0] sc2mac_wt_data42_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1262" *)
  wire [7:0] sc2mac_wt_data43_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1720" *)
  reg [7:0] sc2mac_wt_data43_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1721" *)
  reg [7:0] sc2mac_wt_data43_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1263" *)
  wire [7:0] sc2mac_wt_data44_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1722" *)
  reg [7:0] sc2mac_wt_data44_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1723" *)
  reg [7:0] sc2mac_wt_data44_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1264" *)
  wire [7:0] sc2mac_wt_data45_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1724" *)
  reg [7:0] sc2mac_wt_data45_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1725" *)
  reg [7:0] sc2mac_wt_data45_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1265" *)
  wire [7:0] sc2mac_wt_data46_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1726" *)
  reg [7:0] sc2mac_wt_data46_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1727" *)
  reg [7:0] sc2mac_wt_data46_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1266" *)
  wire [7:0] sc2mac_wt_data47_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1728" *)
  reg [7:0] sc2mac_wt_data47_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1729" *)
  reg [7:0] sc2mac_wt_data47_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1267" *)
  wire [7:0] sc2mac_wt_data48_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1730" *)
  reg [7:0] sc2mac_wt_data48_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1731" *)
  reg [7:0] sc2mac_wt_data48_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1268" *)
  wire [7:0] sc2mac_wt_data49_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1732" *)
  reg [7:0] sc2mac_wt_data49_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1733" *)
  reg [7:0] sc2mac_wt_data49_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1269" *)
  wire [7:0] sc2mac_wt_data4_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1734" *)
  reg [7:0] sc2mac_wt_data4_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1735" *)
  reg [7:0] sc2mac_wt_data4_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1270" *)
  wire [7:0] sc2mac_wt_data50_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1736" *)
  reg [7:0] sc2mac_wt_data50_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1737" *)
  reg [7:0] sc2mac_wt_data50_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1271" *)
  wire [7:0] sc2mac_wt_data51_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1738" *)
  reg [7:0] sc2mac_wt_data51_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1739" *)
  reg [7:0] sc2mac_wt_data51_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1272" *)
  wire [7:0] sc2mac_wt_data52_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1740" *)
  reg [7:0] sc2mac_wt_data52_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1741" *)
  reg [7:0] sc2mac_wt_data52_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1273" *)
  wire [7:0] sc2mac_wt_data53_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1742" *)
  reg [7:0] sc2mac_wt_data53_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1743" *)
  reg [7:0] sc2mac_wt_data53_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1274" *)
  wire [7:0] sc2mac_wt_data54_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1744" *)
  reg [7:0] sc2mac_wt_data54_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1745" *)
  reg [7:0] sc2mac_wt_data54_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1275" *)
  wire [7:0] sc2mac_wt_data55_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1746" *)
  reg [7:0] sc2mac_wt_data55_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1747" *)
  reg [7:0] sc2mac_wt_data55_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1276" *)
  wire [7:0] sc2mac_wt_data56_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1748" *)
  reg [7:0] sc2mac_wt_data56_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1749" *)
  reg [7:0] sc2mac_wt_data56_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1277" *)
  wire [7:0] sc2mac_wt_data57_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1750" *)
  reg [7:0] sc2mac_wt_data57_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1751" *)
  reg [7:0] sc2mac_wt_data57_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1278" *)
  wire [7:0] sc2mac_wt_data58_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1752" *)
  reg [7:0] sc2mac_wt_data58_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1753" *)
  reg [7:0] sc2mac_wt_data58_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1279" *)
  wire [7:0] sc2mac_wt_data59_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1754" *)
  reg [7:0] sc2mac_wt_data59_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1755" *)
  reg [7:0] sc2mac_wt_data59_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1280" *)
  wire [7:0] sc2mac_wt_data5_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1756" *)
  reg [7:0] sc2mac_wt_data5_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1757" *)
  reg [7:0] sc2mac_wt_data5_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1281" *)
  wire [7:0] sc2mac_wt_data60_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1758" *)
  reg [7:0] sc2mac_wt_data60_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1759" *)
  reg [7:0] sc2mac_wt_data60_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1282" *)
  wire [7:0] sc2mac_wt_data61_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1760" *)
  reg [7:0] sc2mac_wt_data61_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1761" *)
  reg [7:0] sc2mac_wt_data61_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1283" *)
  wire [7:0] sc2mac_wt_data62_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1762" *)
  reg [7:0] sc2mac_wt_data62_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1763" *)
  reg [7:0] sc2mac_wt_data62_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1284" *)
  wire [7:0] sc2mac_wt_data63_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1764" *)
  reg [7:0] sc2mac_wt_data63_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1765" *)
  reg [7:0] sc2mac_wt_data63_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1285" *)
  wire [7:0] sc2mac_wt_data64_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1766" *)
  reg [7:0] sc2mac_wt_data64_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1767" *)
  reg [7:0] sc2mac_wt_data64_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1286" *)
  wire [7:0] sc2mac_wt_data65_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1768" *)
  reg [7:0] sc2mac_wt_data65_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1769" *)
  reg [7:0] sc2mac_wt_data65_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1287" *)
  wire [7:0] sc2mac_wt_data66_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1770" *)
  reg [7:0] sc2mac_wt_data66_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1771" *)
  reg [7:0] sc2mac_wt_data66_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1288" *)
  wire [7:0] sc2mac_wt_data67_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1772" *)
  reg [7:0] sc2mac_wt_data67_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1773" *)
  reg [7:0] sc2mac_wt_data67_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1289" *)
  wire [7:0] sc2mac_wt_data68_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1774" *)
  reg [7:0] sc2mac_wt_data68_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1775" *)
  reg [7:0] sc2mac_wt_data68_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1290" *)
  wire [7:0] sc2mac_wt_data69_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1776" *)
  reg [7:0] sc2mac_wt_data69_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1777" *)
  reg [7:0] sc2mac_wt_data69_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1291" *)
  wire [7:0] sc2mac_wt_data6_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1778" *)
  reg [7:0] sc2mac_wt_data6_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1779" *)
  reg [7:0] sc2mac_wt_data6_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1292" *)
  wire [7:0] sc2mac_wt_data70_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1780" *)
  reg [7:0] sc2mac_wt_data70_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1781" *)
  reg [7:0] sc2mac_wt_data70_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1293" *)
  wire [7:0] sc2mac_wt_data71_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1782" *)
  reg [7:0] sc2mac_wt_data71_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1783" *)
  reg [7:0] sc2mac_wt_data71_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1294" *)
  wire [7:0] sc2mac_wt_data72_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1784" *)
  reg [7:0] sc2mac_wt_data72_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1785" *)
  reg [7:0] sc2mac_wt_data72_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1295" *)
  wire [7:0] sc2mac_wt_data73_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1786" *)
  reg [7:0] sc2mac_wt_data73_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1787" *)
  reg [7:0] sc2mac_wt_data73_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1296" *)
  wire [7:0] sc2mac_wt_data74_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1788" *)
  reg [7:0] sc2mac_wt_data74_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1789" *)
  reg [7:0] sc2mac_wt_data74_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1297" *)
  wire [7:0] sc2mac_wt_data75_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1790" *)
  reg [7:0] sc2mac_wt_data75_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1791" *)
  reg [7:0] sc2mac_wt_data75_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1298" *)
  wire [7:0] sc2mac_wt_data76_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1792" *)
  reg [7:0] sc2mac_wt_data76_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1793" *)
  reg [7:0] sc2mac_wt_data76_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1299" *)
  wire [7:0] sc2mac_wt_data77_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1794" *)
  reg [7:0] sc2mac_wt_data77_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1795" *)
  reg [7:0] sc2mac_wt_data77_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1300" *)
  wire [7:0] sc2mac_wt_data78_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1796" *)
  reg [7:0] sc2mac_wt_data78_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1797" *)
  reg [7:0] sc2mac_wt_data78_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1301" *)
  wire [7:0] sc2mac_wt_data79_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1798" *)
  reg [7:0] sc2mac_wt_data79_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1799" *)
  reg [7:0] sc2mac_wt_data79_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1302" *)
  wire [7:0] sc2mac_wt_data7_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1800" *)
  reg [7:0] sc2mac_wt_data7_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1801" *)
  reg [7:0] sc2mac_wt_data7_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1303" *)
  wire [7:0] sc2mac_wt_data80_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1802" *)
  reg [7:0] sc2mac_wt_data80_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1803" *)
  reg [7:0] sc2mac_wt_data80_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1304" *)
  wire [7:0] sc2mac_wt_data81_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1804" *)
  reg [7:0] sc2mac_wt_data81_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1805" *)
  reg [7:0] sc2mac_wt_data81_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1305" *)
  wire [7:0] sc2mac_wt_data82_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1806" *)
  reg [7:0] sc2mac_wt_data82_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1807" *)
  reg [7:0] sc2mac_wt_data82_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1306" *)
  wire [7:0] sc2mac_wt_data83_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1808" *)
  reg [7:0] sc2mac_wt_data83_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1809" *)
  reg [7:0] sc2mac_wt_data83_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1307" *)
  wire [7:0] sc2mac_wt_data84_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1810" *)
  reg [7:0] sc2mac_wt_data84_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1811" *)
  reg [7:0] sc2mac_wt_data84_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1308" *)
  wire [7:0] sc2mac_wt_data85_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1812" *)
  reg [7:0] sc2mac_wt_data85_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1813" *)
  reg [7:0] sc2mac_wt_data85_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1309" *)
  wire [7:0] sc2mac_wt_data86_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1814" *)
  reg [7:0] sc2mac_wt_data86_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1815" *)
  reg [7:0] sc2mac_wt_data86_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1310" *)
  wire [7:0] sc2mac_wt_data87_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1816" *)
  reg [7:0] sc2mac_wt_data87_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1817" *)
  reg [7:0] sc2mac_wt_data87_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1311" *)
  wire [7:0] sc2mac_wt_data88_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1818" *)
  reg [7:0] sc2mac_wt_data88_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1819" *)
  reg [7:0] sc2mac_wt_data88_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1312" *)
  wire [7:0] sc2mac_wt_data89_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1820" *)
  reg [7:0] sc2mac_wt_data89_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1821" *)
  reg [7:0] sc2mac_wt_data89_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1313" *)
  wire [7:0] sc2mac_wt_data8_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1822" *)
  reg [7:0] sc2mac_wt_data8_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1823" *)
  reg [7:0] sc2mac_wt_data8_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1314" *)
  wire [7:0] sc2mac_wt_data90_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1824" *)
  reg [7:0] sc2mac_wt_data90_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1825" *)
  reg [7:0] sc2mac_wt_data90_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1315" *)
  wire [7:0] sc2mac_wt_data91_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1826" *)
  reg [7:0] sc2mac_wt_data91_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1827" *)
  reg [7:0] sc2mac_wt_data91_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1316" *)
  wire [7:0] sc2mac_wt_data92_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1828" *)
  reg [7:0] sc2mac_wt_data92_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1829" *)
  reg [7:0] sc2mac_wt_data92_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1317" *)
  wire [7:0] sc2mac_wt_data93_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1830" *)
  reg [7:0] sc2mac_wt_data93_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1831" *)
  reg [7:0] sc2mac_wt_data93_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1318" *)
  wire [7:0] sc2mac_wt_data94_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1832" *)
  reg [7:0] sc2mac_wt_data94_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1833" *)
  reg [7:0] sc2mac_wt_data94_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1319" *)
  wire [7:0] sc2mac_wt_data95_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1834" *)
  reg [7:0] sc2mac_wt_data95_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1835" *)
  reg [7:0] sc2mac_wt_data95_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1320" *)
  wire [7:0] sc2mac_wt_data96_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1836" *)
  reg [7:0] sc2mac_wt_data96_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1837" *)
  reg [7:0] sc2mac_wt_data96_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1321" *)
  wire [7:0] sc2mac_wt_data97_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1838" *)
  reg [7:0] sc2mac_wt_data97_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1839" *)
  reg [7:0] sc2mac_wt_data97_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1322" *)
  wire [7:0] sc2mac_wt_data98_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1840" *)
  reg [7:0] sc2mac_wt_data98_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1841" *)
  reg [7:0] sc2mac_wt_data98_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1323" *)
  wire [7:0] sc2mac_wt_data99_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1842" *)
  reg [7:0] sc2mac_wt_data99_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1843" *)
  reg [7:0] sc2mac_wt_data99_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1324" *)
  wire [7:0] sc2mac_wt_data9_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1844" *)
  reg [7:0] sc2mac_wt_data9_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1845" *)
  reg [7:0] sc2mac_wt_data9_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:806" *)
  output [7:0] sc2mac_wt_dst_data0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:807" *)
  output [7:0] sc2mac_wt_dst_data1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:816" *)
  output [7:0] sc2mac_wt_dst_data10;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:906" *)
  output [7:0] sc2mac_wt_dst_data100;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:907" *)
  output [7:0] sc2mac_wt_dst_data101;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:908" *)
  output [7:0] sc2mac_wt_dst_data102;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:909" *)
  output [7:0] sc2mac_wt_dst_data103;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:910" *)
  output [7:0] sc2mac_wt_dst_data104;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:911" *)
  output [7:0] sc2mac_wt_dst_data105;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:912" *)
  output [7:0] sc2mac_wt_dst_data106;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:913" *)
  output [7:0] sc2mac_wt_dst_data107;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:914" *)
  output [7:0] sc2mac_wt_dst_data108;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:915" *)
  output [7:0] sc2mac_wt_dst_data109;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:817" *)
  output [7:0] sc2mac_wt_dst_data11;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:916" *)
  output [7:0] sc2mac_wt_dst_data110;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:917" *)
  output [7:0] sc2mac_wt_dst_data111;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:918" *)
  output [7:0] sc2mac_wt_dst_data112;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:919" *)
  output [7:0] sc2mac_wt_dst_data113;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:920" *)
  output [7:0] sc2mac_wt_dst_data114;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:921" *)
  output [7:0] sc2mac_wt_dst_data115;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:922" *)
  output [7:0] sc2mac_wt_dst_data116;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:923" *)
  output [7:0] sc2mac_wt_dst_data117;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:924" *)
  output [7:0] sc2mac_wt_dst_data118;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:925" *)
  output [7:0] sc2mac_wt_dst_data119;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:818" *)
  output [7:0] sc2mac_wt_dst_data12;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:926" *)
  output [7:0] sc2mac_wt_dst_data120;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:927" *)
  output [7:0] sc2mac_wt_dst_data121;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:928" *)
  output [7:0] sc2mac_wt_dst_data122;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:929" *)
  output [7:0] sc2mac_wt_dst_data123;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:930" *)
  output [7:0] sc2mac_wt_dst_data124;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:931" *)
  output [7:0] sc2mac_wt_dst_data125;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:932" *)
  output [7:0] sc2mac_wt_dst_data126;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:933" *)
  output [7:0] sc2mac_wt_dst_data127;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:819" *)
  output [7:0] sc2mac_wt_dst_data13;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:820" *)
  output [7:0] sc2mac_wt_dst_data14;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:821" *)
  output [7:0] sc2mac_wt_dst_data15;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:822" *)
  output [7:0] sc2mac_wt_dst_data16;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:823" *)
  output [7:0] sc2mac_wt_dst_data17;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:824" *)
  output [7:0] sc2mac_wt_dst_data18;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:825" *)
  output [7:0] sc2mac_wt_dst_data19;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:808" *)
  output [7:0] sc2mac_wt_dst_data2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:826" *)
  output [7:0] sc2mac_wt_dst_data20;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:827" *)
  output [7:0] sc2mac_wt_dst_data21;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:828" *)
  output [7:0] sc2mac_wt_dst_data22;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:829" *)
  output [7:0] sc2mac_wt_dst_data23;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:830" *)
  output [7:0] sc2mac_wt_dst_data24;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:831" *)
  output [7:0] sc2mac_wt_dst_data25;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:832" *)
  output [7:0] sc2mac_wt_dst_data26;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:833" *)
  output [7:0] sc2mac_wt_dst_data27;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:834" *)
  output [7:0] sc2mac_wt_dst_data28;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:835" *)
  output [7:0] sc2mac_wt_dst_data29;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:809" *)
  output [7:0] sc2mac_wt_dst_data3;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:836" *)
  output [7:0] sc2mac_wt_dst_data30;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:837" *)
  output [7:0] sc2mac_wt_dst_data31;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:838" *)
  output [7:0] sc2mac_wt_dst_data32;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:839" *)
  output [7:0] sc2mac_wt_dst_data33;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:840" *)
  output [7:0] sc2mac_wt_dst_data34;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:841" *)
  output [7:0] sc2mac_wt_dst_data35;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:842" *)
  output [7:0] sc2mac_wt_dst_data36;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:843" *)
  output [7:0] sc2mac_wt_dst_data37;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:844" *)
  output [7:0] sc2mac_wt_dst_data38;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:845" *)
  output [7:0] sc2mac_wt_dst_data39;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:810" *)
  output [7:0] sc2mac_wt_dst_data4;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:846" *)
  output [7:0] sc2mac_wt_dst_data40;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:847" *)
  output [7:0] sc2mac_wt_dst_data41;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:848" *)
  output [7:0] sc2mac_wt_dst_data42;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:849" *)
  output [7:0] sc2mac_wt_dst_data43;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:850" *)
  output [7:0] sc2mac_wt_dst_data44;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:851" *)
  output [7:0] sc2mac_wt_dst_data45;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:852" *)
  output [7:0] sc2mac_wt_dst_data46;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:853" *)
  output [7:0] sc2mac_wt_dst_data47;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:854" *)
  output [7:0] sc2mac_wt_dst_data48;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:855" *)
  output [7:0] sc2mac_wt_dst_data49;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:811" *)
  output [7:0] sc2mac_wt_dst_data5;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:856" *)
  output [7:0] sc2mac_wt_dst_data50;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:857" *)
  output [7:0] sc2mac_wt_dst_data51;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:858" *)
  output [7:0] sc2mac_wt_dst_data52;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:859" *)
  output [7:0] sc2mac_wt_dst_data53;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:860" *)
  output [7:0] sc2mac_wt_dst_data54;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:861" *)
  output [7:0] sc2mac_wt_dst_data55;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:862" *)
  output [7:0] sc2mac_wt_dst_data56;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:863" *)
  output [7:0] sc2mac_wt_dst_data57;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:864" *)
  output [7:0] sc2mac_wt_dst_data58;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:865" *)
  output [7:0] sc2mac_wt_dst_data59;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:812" *)
  output [7:0] sc2mac_wt_dst_data6;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:866" *)
  output [7:0] sc2mac_wt_dst_data60;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:867" *)
  output [7:0] sc2mac_wt_dst_data61;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:868" *)
  output [7:0] sc2mac_wt_dst_data62;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:869" *)
  output [7:0] sc2mac_wt_dst_data63;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:870" *)
  output [7:0] sc2mac_wt_dst_data64;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:871" *)
  output [7:0] sc2mac_wt_dst_data65;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:872" *)
  output [7:0] sc2mac_wt_dst_data66;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:873" *)
  output [7:0] sc2mac_wt_dst_data67;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:874" *)
  output [7:0] sc2mac_wt_dst_data68;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:875" *)
  output [7:0] sc2mac_wt_dst_data69;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:813" *)
  output [7:0] sc2mac_wt_dst_data7;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:876" *)
  output [7:0] sc2mac_wt_dst_data70;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:877" *)
  output [7:0] sc2mac_wt_dst_data71;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:878" *)
  output [7:0] sc2mac_wt_dst_data72;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:879" *)
  output [7:0] sc2mac_wt_dst_data73;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:880" *)
  output [7:0] sc2mac_wt_dst_data74;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:881" *)
  output [7:0] sc2mac_wt_dst_data75;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:882" *)
  output [7:0] sc2mac_wt_dst_data76;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:883" *)
  output [7:0] sc2mac_wt_dst_data77;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:884" *)
  output [7:0] sc2mac_wt_dst_data78;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:885" *)
  output [7:0] sc2mac_wt_dst_data79;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:814" *)
  output [7:0] sc2mac_wt_dst_data8;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:886" *)
  output [7:0] sc2mac_wt_dst_data80;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:887" *)
  output [7:0] sc2mac_wt_dst_data81;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:888" *)
  output [7:0] sc2mac_wt_dst_data82;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:889" *)
  output [7:0] sc2mac_wt_dst_data83;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:890" *)
  output [7:0] sc2mac_wt_dst_data84;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:891" *)
  output [7:0] sc2mac_wt_dst_data85;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:892" *)
  output [7:0] sc2mac_wt_dst_data86;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:893" *)
  output [7:0] sc2mac_wt_dst_data87;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:894" *)
  output [7:0] sc2mac_wt_dst_data88;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:895" *)
  output [7:0] sc2mac_wt_dst_data89;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:815" *)
  output [7:0] sc2mac_wt_dst_data9;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:896" *)
  output [7:0] sc2mac_wt_dst_data90;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:897" *)
  output [7:0] sc2mac_wt_dst_data91;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:898" *)
  output [7:0] sc2mac_wt_dst_data92;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:899" *)
  output [7:0] sc2mac_wt_dst_data93;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:900" *)
  output [7:0] sc2mac_wt_dst_data94;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:901" *)
  output [7:0] sc2mac_wt_dst_data95;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:902" *)
  output [7:0] sc2mac_wt_dst_data96;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:903" *)
  output [7:0] sc2mac_wt_dst_data97;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:904" *)
  output [7:0] sc2mac_wt_dst_data98;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:905" *)
  output [7:0] sc2mac_wt_dst_data99;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:805" *)
  output [127:0] sc2mac_wt_dst_mask;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:804" *)
  output sc2mac_wt_dst_pvld;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:934" *)
  output [7:0] sc2mac_wt_dst_sel;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1325" *)
  wire [127:0] sc2mac_wt_mask_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1846" *)
  reg [127:0] sc2mac_wt_mask_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1847" *)
  reg [127:0] sc2mac_wt_mask_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1326" *)
  wire sc2mac_wt_pvld_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1848" *)
  reg sc2mac_wt_pvld_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1849" *)
  reg sc2mac_wt_pvld_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1327" *)
  wire [7:0] sc2mac_wt_sel_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1850" *)
  reg [7:0] sc2mac_wt_sel_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:1851" *)
  reg [7:0] sc2mac_wt_sel_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:544" *)
  input [7:0] sc2mac_wt_src_data0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:545" *)
  input [7:0] sc2mac_wt_src_data1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:554" *)
  input [7:0] sc2mac_wt_src_data10;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:644" *)
  input [7:0] sc2mac_wt_src_data100;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:645" *)
  input [7:0] sc2mac_wt_src_data101;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:646" *)
  input [7:0] sc2mac_wt_src_data102;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:647" *)
  input [7:0] sc2mac_wt_src_data103;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:648" *)
  input [7:0] sc2mac_wt_src_data104;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:649" *)
  input [7:0] sc2mac_wt_src_data105;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:650" *)
  input [7:0] sc2mac_wt_src_data106;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:651" *)
  input [7:0] sc2mac_wt_src_data107;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:652" *)
  input [7:0] sc2mac_wt_src_data108;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:653" *)
  input [7:0] sc2mac_wt_src_data109;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:555" *)
  input [7:0] sc2mac_wt_src_data11;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:654" *)
  input [7:0] sc2mac_wt_src_data110;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:655" *)
  input [7:0] sc2mac_wt_src_data111;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:656" *)
  input [7:0] sc2mac_wt_src_data112;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:657" *)
  input [7:0] sc2mac_wt_src_data113;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:658" *)
  input [7:0] sc2mac_wt_src_data114;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:659" *)
  input [7:0] sc2mac_wt_src_data115;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:660" *)
  input [7:0] sc2mac_wt_src_data116;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:661" *)
  input [7:0] sc2mac_wt_src_data117;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:662" *)
  input [7:0] sc2mac_wt_src_data118;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:663" *)
  input [7:0] sc2mac_wt_src_data119;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:556" *)
  input [7:0] sc2mac_wt_src_data12;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:664" *)
  input [7:0] sc2mac_wt_src_data120;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:665" *)
  input [7:0] sc2mac_wt_src_data121;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:666" *)
  input [7:0] sc2mac_wt_src_data122;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:667" *)
  input [7:0] sc2mac_wt_src_data123;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:668" *)
  input [7:0] sc2mac_wt_src_data124;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:669" *)
  input [7:0] sc2mac_wt_src_data125;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:670" *)
  input [7:0] sc2mac_wt_src_data126;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:671" *)
  input [7:0] sc2mac_wt_src_data127;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:557" *)
  input [7:0] sc2mac_wt_src_data13;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:558" *)
  input [7:0] sc2mac_wt_src_data14;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:559" *)
  input [7:0] sc2mac_wt_src_data15;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:560" *)
  input [7:0] sc2mac_wt_src_data16;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:561" *)
  input [7:0] sc2mac_wt_src_data17;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:562" *)
  input [7:0] sc2mac_wt_src_data18;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:563" *)
  input [7:0] sc2mac_wt_src_data19;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:546" *)
  input [7:0] sc2mac_wt_src_data2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:564" *)
  input [7:0] sc2mac_wt_src_data20;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:565" *)
  input [7:0] sc2mac_wt_src_data21;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:566" *)
  input [7:0] sc2mac_wt_src_data22;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:567" *)
  input [7:0] sc2mac_wt_src_data23;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:568" *)
  input [7:0] sc2mac_wt_src_data24;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:569" *)
  input [7:0] sc2mac_wt_src_data25;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:570" *)
  input [7:0] sc2mac_wt_src_data26;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:571" *)
  input [7:0] sc2mac_wt_src_data27;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:572" *)
  input [7:0] sc2mac_wt_src_data28;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:573" *)
  input [7:0] sc2mac_wt_src_data29;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:547" *)
  input [7:0] sc2mac_wt_src_data3;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:574" *)
  input [7:0] sc2mac_wt_src_data30;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:575" *)
  input [7:0] sc2mac_wt_src_data31;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:576" *)
  input [7:0] sc2mac_wt_src_data32;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:577" *)
  input [7:0] sc2mac_wt_src_data33;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:578" *)
  input [7:0] sc2mac_wt_src_data34;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:579" *)
  input [7:0] sc2mac_wt_src_data35;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:580" *)
  input [7:0] sc2mac_wt_src_data36;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:581" *)
  input [7:0] sc2mac_wt_src_data37;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:582" *)
  input [7:0] sc2mac_wt_src_data38;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:583" *)
  input [7:0] sc2mac_wt_src_data39;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:548" *)
  input [7:0] sc2mac_wt_src_data4;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:584" *)
  input [7:0] sc2mac_wt_src_data40;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:585" *)
  input [7:0] sc2mac_wt_src_data41;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:586" *)
  input [7:0] sc2mac_wt_src_data42;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:587" *)
  input [7:0] sc2mac_wt_src_data43;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:588" *)
  input [7:0] sc2mac_wt_src_data44;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:589" *)
  input [7:0] sc2mac_wt_src_data45;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:590" *)
  input [7:0] sc2mac_wt_src_data46;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:591" *)
  input [7:0] sc2mac_wt_src_data47;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:592" *)
  input [7:0] sc2mac_wt_src_data48;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:593" *)
  input [7:0] sc2mac_wt_src_data49;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:549" *)
  input [7:0] sc2mac_wt_src_data5;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:594" *)
  input [7:0] sc2mac_wt_src_data50;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:595" *)
  input [7:0] sc2mac_wt_src_data51;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:596" *)
  input [7:0] sc2mac_wt_src_data52;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:597" *)
  input [7:0] sc2mac_wt_src_data53;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:598" *)
  input [7:0] sc2mac_wt_src_data54;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:599" *)
  input [7:0] sc2mac_wt_src_data55;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:600" *)
  input [7:0] sc2mac_wt_src_data56;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:601" *)
  input [7:0] sc2mac_wt_src_data57;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:602" *)
  input [7:0] sc2mac_wt_src_data58;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:603" *)
  input [7:0] sc2mac_wt_src_data59;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:550" *)
  input [7:0] sc2mac_wt_src_data6;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:604" *)
  input [7:0] sc2mac_wt_src_data60;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:605" *)
  input [7:0] sc2mac_wt_src_data61;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:606" *)
  input [7:0] sc2mac_wt_src_data62;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:607" *)
  input [7:0] sc2mac_wt_src_data63;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:608" *)
  input [7:0] sc2mac_wt_src_data64;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:609" *)
  input [7:0] sc2mac_wt_src_data65;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:610" *)
  input [7:0] sc2mac_wt_src_data66;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:611" *)
  input [7:0] sc2mac_wt_src_data67;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:612" *)
  input [7:0] sc2mac_wt_src_data68;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:613" *)
  input [7:0] sc2mac_wt_src_data69;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:551" *)
  input [7:0] sc2mac_wt_src_data7;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:614" *)
  input [7:0] sc2mac_wt_src_data70;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:615" *)
  input [7:0] sc2mac_wt_src_data71;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:616" *)
  input [7:0] sc2mac_wt_src_data72;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:617" *)
  input [7:0] sc2mac_wt_src_data73;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:618" *)
  input [7:0] sc2mac_wt_src_data74;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:619" *)
  input [7:0] sc2mac_wt_src_data75;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:620" *)
  input [7:0] sc2mac_wt_src_data76;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:621" *)
  input [7:0] sc2mac_wt_src_data77;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:622" *)
  input [7:0] sc2mac_wt_src_data78;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:623" *)
  input [7:0] sc2mac_wt_src_data79;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:552" *)
  input [7:0] sc2mac_wt_src_data8;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:624" *)
  input [7:0] sc2mac_wt_src_data80;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:625" *)
  input [7:0] sc2mac_wt_src_data81;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:626" *)
  input [7:0] sc2mac_wt_src_data82;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:627" *)
  input [7:0] sc2mac_wt_src_data83;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:628" *)
  input [7:0] sc2mac_wt_src_data84;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:629" *)
  input [7:0] sc2mac_wt_src_data85;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:630" *)
  input [7:0] sc2mac_wt_src_data86;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:631" *)
  input [7:0] sc2mac_wt_src_data87;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:632" *)
  input [7:0] sc2mac_wt_src_data88;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:633" *)
  input [7:0] sc2mac_wt_src_data89;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:553" *)
  input [7:0] sc2mac_wt_src_data9;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:634" *)
  input [7:0] sc2mac_wt_src_data90;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:635" *)
  input [7:0] sc2mac_wt_src_data91;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:636" *)
  input [7:0] sc2mac_wt_src_data92;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:637" *)
  input [7:0] sc2mac_wt_src_data93;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:638" *)
  input [7:0] sc2mac_wt_src_data94;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:639" *)
  input [7:0] sc2mac_wt_src_data95;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:640" *)
  input [7:0] sc2mac_wt_src_data96;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:641" *)
  input [7:0] sc2mac_wt_src_data97;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:642" *)
  input [7:0] sc2mac_wt_src_data98;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:643" *)
  input [7:0] sc2mac_wt_src_data99;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:543" *)
  input [127:0] sc2mac_wt_src_mask;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:542" *)
  input sc2mac_wt_src_pvld;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:672" *)
  input [7:0] sc2mac_wt_src_sel;
  assign _0520_ = sc2mac_wt_src_pvld | (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:2125" *) sc2mac_wt_pvld_d1;
  assign _0521_ = sc2mac_dat_src_pvld | (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:3534" *) sc2mac_dat_pvld_d1;
  assign _0522_ = sc2mac_wt_pvld_d1 | (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:4943" *) sc2mac_wt_pvld_d2;
  assign _0523_ = sc2mac_dat_pvld_d1 | (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:6352" *) sc2mac_dat_pvld_d2;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data127_d2 <= _0061_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data126_d2 <= _0059_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data125_d2 <= _0057_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data124_d2 <= _0055_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data123_d2 <= _0053_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data122_d2 <= _0051_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data121_d2 <= _0049_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data120_d2 <= _0047_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data119_d2 <= _0043_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data118_d2 <= _0041_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data117_d2 <= _0039_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data116_d2 <= _0037_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data115_d2 <= _0035_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data114_d2 <= _0033_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data113_d2 <= _0031_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data112_d2 <= _0029_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data111_d2 <= _0027_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data110_d2 <= _0025_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data109_d2 <= _0021_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data108_d2 <= _0019_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data107_d2 <= _0017_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data106_d2 <= _0015_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data105_d2 <= _0013_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data104_d2 <= _0011_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data103_d2 <= _0009_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data102_d2 <= _0007_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data101_d2 <= _0005_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data100_d2 <= _0003_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data99_d2 <= _0253_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data98_d2 <= _0251_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data97_d2 <= _0249_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data96_d2 <= _0247_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data95_d2 <= _0245_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data94_d2 <= _0243_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data93_d2 <= _0241_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data92_d2 <= _0239_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data91_d2 <= _0237_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data90_d2 <= _0235_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data89_d2 <= _0231_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data88_d2 <= _0229_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data87_d2 <= _0227_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data86_d2 <= _0225_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data85_d2 <= _0223_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data84_d2 <= _0221_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data83_d2 <= _0219_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data82_d2 <= _0217_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data81_d2 <= _0215_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data80_d2 <= _0213_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data79_d2 <= _0209_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data78_d2 <= _0207_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data77_d2 <= _0205_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data76_d2 <= _0203_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data75_d2 <= _0201_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data74_d2 <= _0199_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data73_d2 <= _0197_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data72_d2 <= _0195_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data71_d2 <= _0193_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data70_d2 <= _0191_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data69_d2 <= _0187_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data68_d2 <= _0185_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data67_d2 <= _0183_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data66_d2 <= _0181_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data65_d2 <= _0179_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data64_d2 <= _0177_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data63_d2 <= _0175_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data62_d2 <= _0173_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data61_d2 <= _0171_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data60_d2 <= _0169_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data59_d2 <= _0165_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data58_d2 <= _0163_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data57_d2 <= _0161_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data56_d2 <= _0159_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data55_d2 <= _0157_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data54_d2 <= _0155_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data53_d2 <= _0153_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data52_d2 <= _0151_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data51_d2 <= _0149_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data50_d2 <= _0147_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data49_d2 <= _0143_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data48_d2 <= _0141_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data47_d2 <= _0139_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data46_d2 <= _0137_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data45_d2 <= _0135_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data44_d2 <= _0133_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data43_d2 <= _0131_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data42_d2 <= _0129_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data41_d2 <= _0127_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data40_d2 <= _0125_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data39_d2 <= _0121_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data38_d2 <= _0119_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data37_d2 <= _0117_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data36_d2 <= _0115_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data35_d2 <= _0113_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data34_d2 <= _0111_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data33_d2 <= _0109_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data32_d2 <= _0107_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data31_d2 <= _0105_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data30_d2 <= _0103_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data29_d2 <= _0099_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data28_d2 <= _0097_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data27_d2 <= _0095_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data26_d2 <= _0093_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data25_d2 <= _0091_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data24_d2 <= _0089_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data23_d2 <= _0087_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data22_d2 <= _0085_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data21_d2 <= _0083_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data20_d2 <= _0081_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data19_d2 <= _0077_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data18_d2 <= _0075_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data17_d2 <= _0073_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data16_d2 <= _0071_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data15_d2 <= _0069_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data14_d2 <= _0067_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data13_d2 <= _0065_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data12_d2 <= _0063_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data11_d2 <= _0045_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data10_d2 <= _0023_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data9_d2 <= _0255_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data8_d2 <= _0233_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data7_d2 <= _0211_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data6_d2 <= _0189_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data5_d2 <= _0167_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data4_d2 <= _0145_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data3_d2 <= _0123_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data2_d2 <= _0101_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data1_d2 <= _0079_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data0_d2 <= _0001_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      sc2mac_dat_mask_d2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    else
      sc2mac_dat_mask_d2 <= _0257_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      sc2mac_dat_pd_d2 <= 9'b000000000;
    else
      sc2mac_dat_pd_d2 <= _0259_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      sc2mac_dat_pvld_d2 <= 1'b0;
    else
      sc2mac_dat_pvld_d2 <= sc2mac_dat_pvld_d1;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data127_d2 <= _0321_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data126_d2 <= _0319_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data125_d2 <= _0317_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data124_d2 <= _0315_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data123_d2 <= _0313_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data122_d2 <= _0311_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data121_d2 <= _0309_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data120_d2 <= _0307_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data119_d2 <= _0303_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data118_d2 <= _0301_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data117_d2 <= _0299_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data116_d2 <= _0297_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data115_d2 <= _0295_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data114_d2 <= _0293_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data113_d2 <= _0291_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data112_d2 <= _0289_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data111_d2 <= _0287_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data110_d2 <= _0285_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data109_d2 <= _0281_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data108_d2 <= _0279_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data107_d2 <= _0277_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data106_d2 <= _0275_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data105_d2 <= _0273_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data104_d2 <= _0271_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data103_d2 <= _0269_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data102_d2 <= _0267_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data101_d2 <= _0265_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data100_d2 <= _0263_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data99_d2 <= _0513_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data98_d2 <= _0511_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data97_d2 <= _0509_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data96_d2 <= _0507_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data95_d2 <= _0505_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data94_d2 <= _0503_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data93_d2 <= _0501_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data92_d2 <= _0499_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data91_d2 <= _0497_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data90_d2 <= _0495_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data89_d2 <= _0491_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data88_d2 <= _0489_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data87_d2 <= _0487_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data86_d2 <= _0485_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data85_d2 <= _0483_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data84_d2 <= _0481_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data83_d2 <= _0479_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data82_d2 <= _0477_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data81_d2 <= _0475_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data80_d2 <= _0473_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data79_d2 <= _0469_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data78_d2 <= _0467_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data77_d2 <= _0465_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data76_d2 <= _0463_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data75_d2 <= _0461_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data74_d2 <= _0459_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data73_d2 <= _0457_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data72_d2 <= _0455_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data71_d2 <= _0453_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data70_d2 <= _0451_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data69_d2 <= _0447_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data68_d2 <= _0445_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data67_d2 <= _0443_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data66_d2 <= _0441_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data65_d2 <= _0439_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data64_d2 <= _0437_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data63_d2 <= _0435_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data62_d2 <= _0433_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data61_d2 <= _0431_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data60_d2 <= _0429_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data59_d2 <= _0425_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data58_d2 <= _0423_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data57_d2 <= _0421_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data56_d2 <= _0419_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data55_d2 <= _0417_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data54_d2 <= _0415_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data53_d2 <= _0413_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data52_d2 <= _0411_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data51_d2 <= _0409_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data50_d2 <= _0407_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data49_d2 <= _0403_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data48_d2 <= _0401_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data47_d2 <= _0399_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data46_d2 <= _0397_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data45_d2 <= _0395_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data44_d2 <= _0393_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data43_d2 <= _0391_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data42_d2 <= _0389_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data41_d2 <= _0387_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data40_d2 <= _0385_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data39_d2 <= _0381_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data38_d2 <= _0379_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data37_d2 <= _0377_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data36_d2 <= _0375_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data35_d2 <= _0373_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data34_d2 <= _0371_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data33_d2 <= _0369_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data32_d2 <= _0367_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data31_d2 <= _0365_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data30_d2 <= _0363_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data29_d2 <= _0359_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data28_d2 <= _0357_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data27_d2 <= _0355_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data26_d2 <= _0353_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data25_d2 <= _0351_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data24_d2 <= _0349_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data23_d2 <= _0347_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data22_d2 <= _0345_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data21_d2 <= _0343_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data20_d2 <= _0341_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data19_d2 <= _0337_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data18_d2 <= _0335_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data17_d2 <= _0333_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data16_d2 <= _0331_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data15_d2 <= _0329_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data14_d2 <= _0327_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data13_d2 <= _0325_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data12_d2 <= _0323_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data11_d2 <= _0305_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data10_d2 <= _0283_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data9_d2 <= _0515_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data8_d2 <= _0493_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data7_d2 <= _0471_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data6_d2 <= _0449_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data5_d2 <= _0427_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data4_d2 <= _0405_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data3_d2 <= _0383_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data2_d2 <= _0361_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data1_d2 <= _0339_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data0_d2 <= _0261_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      sc2mac_wt_mask_d2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    else
      sc2mac_wt_mask_d2 <= _0517_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      sc2mac_wt_sel_d2 <= 8'b00000000;
    else
      sc2mac_wt_sel_d2 <= _0519_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      sc2mac_wt_pvld_d2 <= 1'b0;
    else
      sc2mac_wt_pvld_d2 <= sc2mac_wt_pvld_d1;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data127_d1 <= _0060_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data126_d1 <= _0058_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data125_d1 <= _0056_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data124_d1 <= _0054_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data123_d1 <= _0052_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data122_d1 <= _0050_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data121_d1 <= _0048_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data120_d1 <= _0046_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data119_d1 <= _0042_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data118_d1 <= _0040_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data117_d1 <= _0038_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data116_d1 <= _0036_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data115_d1 <= _0034_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data114_d1 <= _0032_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data113_d1 <= _0030_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data112_d1 <= _0028_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data111_d1 <= _0026_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data110_d1 <= _0024_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data109_d1 <= _0020_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data108_d1 <= _0018_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data107_d1 <= _0016_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data106_d1 <= _0014_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data105_d1 <= _0012_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data104_d1 <= _0010_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data103_d1 <= _0008_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data102_d1 <= _0006_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data101_d1 <= _0004_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data100_d1 <= _0002_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data99_d1 <= _0252_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data98_d1 <= _0250_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data97_d1 <= _0248_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data96_d1 <= _0246_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data95_d1 <= _0244_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data94_d1 <= _0242_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data93_d1 <= _0240_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data92_d1 <= _0238_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data91_d1 <= _0236_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data90_d1 <= _0234_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data89_d1 <= _0230_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data88_d1 <= _0228_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data87_d1 <= _0226_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data86_d1 <= _0224_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data85_d1 <= _0222_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data84_d1 <= _0220_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data83_d1 <= _0218_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data82_d1 <= _0216_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data81_d1 <= _0214_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data80_d1 <= _0212_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data79_d1 <= _0208_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data78_d1 <= _0206_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data77_d1 <= _0204_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data76_d1 <= _0202_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data75_d1 <= _0200_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data74_d1 <= _0198_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data73_d1 <= _0196_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data72_d1 <= _0194_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data71_d1 <= _0192_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data70_d1 <= _0190_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data69_d1 <= _0186_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data68_d1 <= _0184_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data67_d1 <= _0182_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data66_d1 <= _0180_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data65_d1 <= _0178_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data64_d1 <= _0176_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data63_d1 <= _0174_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data62_d1 <= _0172_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data61_d1 <= _0170_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data60_d1 <= _0168_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data59_d1 <= _0164_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data58_d1 <= _0162_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data57_d1 <= _0160_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data56_d1 <= _0158_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data55_d1 <= _0156_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data54_d1 <= _0154_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data53_d1 <= _0152_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data52_d1 <= _0150_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data51_d1 <= _0148_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data50_d1 <= _0146_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data49_d1 <= _0142_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data48_d1 <= _0140_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data47_d1 <= _0138_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data46_d1 <= _0136_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data45_d1 <= _0134_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data44_d1 <= _0132_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data43_d1 <= _0130_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data42_d1 <= _0128_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data41_d1 <= _0126_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data40_d1 <= _0124_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data39_d1 <= _0120_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data38_d1 <= _0118_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data37_d1 <= _0116_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data36_d1 <= _0114_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data35_d1 <= _0112_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data34_d1 <= _0110_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data33_d1 <= _0108_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data32_d1 <= _0106_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data31_d1 <= _0104_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data30_d1 <= _0102_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data29_d1 <= _0098_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data28_d1 <= _0096_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data27_d1 <= _0094_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data26_d1 <= _0092_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data25_d1 <= _0090_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data24_d1 <= _0088_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data23_d1 <= _0086_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data22_d1 <= _0084_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data21_d1 <= _0082_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data20_d1 <= _0080_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data19_d1 <= _0076_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data18_d1 <= _0074_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data17_d1 <= _0072_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data16_d1 <= _0070_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data15_d1 <= _0068_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data14_d1 <= _0066_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data13_d1 <= _0064_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data12_d1 <= _0062_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data11_d1 <= _0044_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data10_d1 <= _0022_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data9_d1 <= _0254_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data8_d1 <= _0232_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data7_d1 <= _0210_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data6_d1 <= _0188_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data5_d1 <= _0166_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data4_d1 <= _0144_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data3_d1 <= _0122_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data2_d1 <= _0100_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data1_d1 <= _0078_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data0_d1 <= _0000_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      sc2mac_dat_mask_d1 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    else
      sc2mac_dat_mask_d1 <= _0256_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      sc2mac_dat_pd_d1 <= 9'b000000000;
    else
      sc2mac_dat_pd_d1 <= _0258_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      sc2mac_dat_pvld_d1 <= 1'b0;
    else
      sc2mac_dat_pvld_d1 <= sc2mac_dat_src_pvld;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data127_d1 <= _0320_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data126_d1 <= _0318_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data125_d1 <= _0316_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data124_d1 <= _0314_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data123_d1 <= _0312_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data122_d1 <= _0310_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data121_d1 <= _0308_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data120_d1 <= _0306_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data119_d1 <= _0302_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data118_d1 <= _0300_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data117_d1 <= _0298_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data116_d1 <= _0296_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data115_d1 <= _0294_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data114_d1 <= _0292_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data113_d1 <= _0290_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data112_d1 <= _0288_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data111_d1 <= _0286_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data110_d1 <= _0284_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data109_d1 <= _0280_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data108_d1 <= _0278_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data107_d1 <= _0276_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data106_d1 <= _0274_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data105_d1 <= _0272_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data104_d1 <= _0270_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data103_d1 <= _0268_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data102_d1 <= _0266_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data101_d1 <= _0264_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data100_d1 <= _0262_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data99_d1 <= _0512_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data98_d1 <= _0510_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data97_d1 <= _0508_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data96_d1 <= _0506_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data95_d1 <= _0504_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data94_d1 <= _0502_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data93_d1 <= _0500_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data92_d1 <= _0498_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data91_d1 <= _0496_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data90_d1 <= _0494_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data89_d1 <= _0490_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data88_d1 <= _0488_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data87_d1 <= _0486_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data86_d1 <= _0484_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data85_d1 <= _0482_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data84_d1 <= _0480_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data83_d1 <= _0478_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data82_d1 <= _0476_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data81_d1 <= _0474_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data80_d1 <= _0472_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data79_d1 <= _0468_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data78_d1 <= _0466_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data77_d1 <= _0464_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data76_d1 <= _0462_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data75_d1 <= _0460_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data74_d1 <= _0458_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data73_d1 <= _0456_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data72_d1 <= _0454_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data71_d1 <= _0452_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data70_d1 <= _0450_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data69_d1 <= _0446_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data68_d1 <= _0444_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data67_d1 <= _0442_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data66_d1 <= _0440_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data65_d1 <= _0438_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data64_d1 <= _0436_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data63_d1 <= _0434_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data62_d1 <= _0432_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data61_d1 <= _0430_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data60_d1 <= _0428_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data59_d1 <= _0424_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data58_d1 <= _0422_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data57_d1 <= _0420_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data56_d1 <= _0418_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data55_d1 <= _0416_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data54_d1 <= _0414_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data53_d1 <= _0412_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data52_d1 <= _0410_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data51_d1 <= _0408_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data50_d1 <= _0406_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data49_d1 <= _0402_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data48_d1 <= _0400_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data47_d1 <= _0398_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data46_d1 <= _0396_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data45_d1 <= _0394_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data44_d1 <= _0392_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data43_d1 <= _0390_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data42_d1 <= _0388_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data41_d1 <= _0386_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data40_d1 <= _0384_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data39_d1 <= _0380_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data38_d1 <= _0378_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data37_d1 <= _0376_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data36_d1 <= _0374_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data35_d1 <= _0372_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data34_d1 <= _0370_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data33_d1 <= _0368_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data32_d1 <= _0366_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data31_d1 <= _0364_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data30_d1 <= _0362_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data29_d1 <= _0358_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data28_d1 <= _0356_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data27_d1 <= _0354_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data26_d1 <= _0352_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data25_d1 <= _0350_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data24_d1 <= _0348_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data23_d1 <= _0346_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data22_d1 <= _0344_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data21_d1 <= _0342_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data20_d1 <= _0340_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data19_d1 <= _0336_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data18_d1 <= _0334_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data17_d1 <= _0332_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data16_d1 <= _0330_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data15_d1 <= _0328_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data14_d1 <= _0326_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data13_d1 <= _0324_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data12_d1 <= _0322_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data11_d1 <= _0304_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data10_d1 <= _0282_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data9_d1 <= _0514_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data8_d1 <= _0492_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data7_d1 <= _0470_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data6_d1 <= _0448_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data5_d1 <= _0426_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data4_d1 <= _0404_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data3_d1 <= _0382_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data2_d1 <= _0360_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data1_d1 <= _0338_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data0_d1 <= _0260_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      sc2mac_wt_mask_d1 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    else
      sc2mac_wt_mask_d1 <= _0516_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      sc2mac_wt_sel_d1 <= 8'b00000000;
    else
      sc2mac_wt_sel_d1 <= _0518_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      sc2mac_wt_pvld_d1 <= 1'b0;
    else
      sc2mac_wt_pvld_d1 <= sc2mac_wt_src_pvld;
  assign _0061_ = sc2mac_dat_mask_d1[127] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:7741" *) sc2mac_dat_data127_d1 : sc2mac_dat_data127_d2;
  assign _0059_ = sc2mac_dat_mask_d1[126] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:7731" *) sc2mac_dat_data126_d1 : sc2mac_dat_data126_d2;
  assign _0057_ = sc2mac_dat_mask_d1[125] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:7721" *) sc2mac_dat_data125_d1 : sc2mac_dat_data125_d2;
  assign _0055_ = sc2mac_dat_mask_d1[124] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:7711" *) sc2mac_dat_data124_d1 : sc2mac_dat_data124_d2;
  assign _0053_ = sc2mac_dat_mask_d1[123] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:7701" *) sc2mac_dat_data123_d1 : sc2mac_dat_data123_d2;
  assign _0051_ = sc2mac_dat_mask_d1[122] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:7691" *) sc2mac_dat_data122_d1 : sc2mac_dat_data122_d2;
  assign _0049_ = sc2mac_dat_mask_d1[121] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:7681" *) sc2mac_dat_data121_d1 : sc2mac_dat_data121_d2;
  assign _0047_ = sc2mac_dat_mask_d1[120] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:7671" *) sc2mac_dat_data120_d1 : sc2mac_dat_data120_d2;
  assign _0043_ = sc2mac_dat_mask_d1[119] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:7661" *) sc2mac_dat_data119_d1 : sc2mac_dat_data119_d2;
  assign _0041_ = sc2mac_dat_mask_d1[118] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:7651" *) sc2mac_dat_data118_d1 : sc2mac_dat_data118_d2;
  assign _0039_ = sc2mac_dat_mask_d1[117] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:7641" *) sc2mac_dat_data117_d1 : sc2mac_dat_data117_d2;
  assign _0037_ = sc2mac_dat_mask_d1[116] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:7631" *) sc2mac_dat_data116_d1 : sc2mac_dat_data116_d2;
  assign _0035_ = sc2mac_dat_mask_d1[115] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:7621" *) sc2mac_dat_data115_d1 : sc2mac_dat_data115_d2;
  assign _0033_ = sc2mac_dat_mask_d1[114] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:7611" *) sc2mac_dat_data114_d1 : sc2mac_dat_data114_d2;
  assign _0031_ = sc2mac_dat_mask_d1[113] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:7601" *) sc2mac_dat_data113_d1 : sc2mac_dat_data113_d2;
  assign _0029_ = sc2mac_dat_mask_d1[112] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:7591" *) sc2mac_dat_data112_d1 : sc2mac_dat_data112_d2;
  assign _0027_ = sc2mac_dat_mask_d1[111] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:7581" *) sc2mac_dat_data111_d1 : sc2mac_dat_data111_d2;
  assign _0025_ = sc2mac_dat_mask_d1[110] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:7571" *) sc2mac_dat_data110_d1 : sc2mac_dat_data110_d2;
  assign _0021_ = sc2mac_dat_mask_d1[109] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:7561" *) sc2mac_dat_data109_d1 : sc2mac_dat_data109_d2;
  assign _0019_ = sc2mac_dat_mask_d1[108] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:7551" *) sc2mac_dat_data108_d1 : sc2mac_dat_data108_d2;
  assign _0017_ = sc2mac_dat_mask_d1[107] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:7541" *) sc2mac_dat_data107_d1 : sc2mac_dat_data107_d2;
  assign _0015_ = sc2mac_dat_mask_d1[106] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:7531" *) sc2mac_dat_data106_d1 : sc2mac_dat_data106_d2;
  assign _0013_ = sc2mac_dat_mask_d1[105] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:7521" *) sc2mac_dat_data105_d1 : sc2mac_dat_data105_d2;
  assign _0011_ = sc2mac_dat_mask_d1[104] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:7511" *) sc2mac_dat_data104_d1 : sc2mac_dat_data104_d2;
  assign _0009_ = sc2mac_dat_mask_d1[103] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:7501" *) sc2mac_dat_data103_d1 : sc2mac_dat_data103_d2;
  assign _0007_ = sc2mac_dat_mask_d1[102] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:7491" *) sc2mac_dat_data102_d1 : sc2mac_dat_data102_d2;
  assign _0005_ = sc2mac_dat_mask_d1[101] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:7481" *) sc2mac_dat_data101_d1 : sc2mac_dat_data101_d2;
  assign _0003_ = sc2mac_dat_mask_d1[100] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:7471" *) sc2mac_dat_data100_d1 : sc2mac_dat_data100_d2;
  assign _0253_ = sc2mac_dat_mask_d1[99] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:7461" *) sc2mac_dat_data99_d1 : sc2mac_dat_data99_d2;
  assign _0251_ = sc2mac_dat_mask_d1[98] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:7451" *) sc2mac_dat_data98_d1 : sc2mac_dat_data98_d2;
  assign _0249_ = sc2mac_dat_mask_d1[97] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:7441" *) sc2mac_dat_data97_d1 : sc2mac_dat_data97_d2;
  assign _0247_ = sc2mac_dat_mask_d1[96] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:7431" *) sc2mac_dat_data96_d1 : sc2mac_dat_data96_d2;
  assign _0245_ = sc2mac_dat_mask_d1[95] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:7421" *) sc2mac_dat_data95_d1 : sc2mac_dat_data95_d2;
  assign _0243_ = sc2mac_dat_mask_d1[94] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:7411" *) sc2mac_dat_data94_d1 : sc2mac_dat_data94_d2;
  assign _0241_ = sc2mac_dat_mask_d1[93] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:7401" *) sc2mac_dat_data93_d1 : sc2mac_dat_data93_d2;
  assign _0239_ = sc2mac_dat_mask_d1[92] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:7391" *) sc2mac_dat_data92_d1 : sc2mac_dat_data92_d2;
  assign _0237_ = sc2mac_dat_mask_d1[91] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:7381" *) sc2mac_dat_data91_d1 : sc2mac_dat_data91_d2;
  assign _0235_ = sc2mac_dat_mask_d1[90] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:7371" *) sc2mac_dat_data90_d1 : sc2mac_dat_data90_d2;
  assign _0231_ = sc2mac_dat_mask_d1[89] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:7361" *) sc2mac_dat_data89_d1 : sc2mac_dat_data89_d2;
  assign _0229_ = sc2mac_dat_mask_d1[88] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:7351" *) sc2mac_dat_data88_d1 : sc2mac_dat_data88_d2;
  assign _0227_ = sc2mac_dat_mask_d1[87] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:7341" *) sc2mac_dat_data87_d1 : sc2mac_dat_data87_d2;
  assign _0225_ = sc2mac_dat_mask_d1[86] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:7331" *) sc2mac_dat_data86_d1 : sc2mac_dat_data86_d2;
  assign _0223_ = sc2mac_dat_mask_d1[85] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:7321" *) sc2mac_dat_data85_d1 : sc2mac_dat_data85_d2;
  assign _0221_ = sc2mac_dat_mask_d1[84] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:7311" *) sc2mac_dat_data84_d1 : sc2mac_dat_data84_d2;
  assign _0219_ = sc2mac_dat_mask_d1[83] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:7301" *) sc2mac_dat_data83_d1 : sc2mac_dat_data83_d2;
  assign _0217_ = sc2mac_dat_mask_d1[82] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:7291" *) sc2mac_dat_data82_d1 : sc2mac_dat_data82_d2;
  assign _0215_ = sc2mac_dat_mask_d1[81] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:7281" *) sc2mac_dat_data81_d1 : sc2mac_dat_data81_d2;
  assign _0213_ = sc2mac_dat_mask_d1[80] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:7271" *) sc2mac_dat_data80_d1 : sc2mac_dat_data80_d2;
  assign _0209_ = sc2mac_dat_mask_d1[79] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:7261" *) sc2mac_dat_data79_d1 : sc2mac_dat_data79_d2;
  assign _0207_ = sc2mac_dat_mask_d1[78] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:7251" *) sc2mac_dat_data78_d1 : sc2mac_dat_data78_d2;
  assign _0205_ = sc2mac_dat_mask_d1[77] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:7241" *) sc2mac_dat_data77_d1 : sc2mac_dat_data77_d2;
  assign _0203_ = sc2mac_dat_mask_d1[76] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:7231" *) sc2mac_dat_data76_d1 : sc2mac_dat_data76_d2;
  assign _0201_ = sc2mac_dat_mask_d1[75] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:7221" *) sc2mac_dat_data75_d1 : sc2mac_dat_data75_d2;
  assign _0199_ = sc2mac_dat_mask_d1[74] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:7211" *) sc2mac_dat_data74_d1 : sc2mac_dat_data74_d2;
  assign _0197_ = sc2mac_dat_mask_d1[73] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:7201" *) sc2mac_dat_data73_d1 : sc2mac_dat_data73_d2;
  assign _0195_ = sc2mac_dat_mask_d1[72] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:7191" *) sc2mac_dat_data72_d1 : sc2mac_dat_data72_d2;
  assign _0193_ = sc2mac_dat_mask_d1[71] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:7181" *) sc2mac_dat_data71_d1 : sc2mac_dat_data71_d2;
  assign _0191_ = sc2mac_dat_mask_d1[70] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:7171" *) sc2mac_dat_data70_d1 : sc2mac_dat_data70_d2;
  assign _0187_ = sc2mac_dat_mask_d1[69] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:7161" *) sc2mac_dat_data69_d1 : sc2mac_dat_data69_d2;
  assign _0185_ = sc2mac_dat_mask_d1[68] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:7151" *) sc2mac_dat_data68_d1 : sc2mac_dat_data68_d2;
  assign _0183_ = sc2mac_dat_mask_d1[67] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:7141" *) sc2mac_dat_data67_d1 : sc2mac_dat_data67_d2;
  assign _0181_ = sc2mac_dat_mask_d1[66] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:7131" *) sc2mac_dat_data66_d1 : sc2mac_dat_data66_d2;
  assign _0179_ = sc2mac_dat_mask_d1[65] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:7121" *) sc2mac_dat_data65_d1 : sc2mac_dat_data65_d2;
  assign _0177_ = sc2mac_dat_mask_d1[64] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:7111" *) sc2mac_dat_data64_d1 : sc2mac_dat_data64_d2;
  assign _0175_ = sc2mac_dat_mask_d1[63] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:7101" *) sc2mac_dat_data63_d1 : sc2mac_dat_data63_d2;
  assign _0173_ = sc2mac_dat_mask_d1[62] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:7091" *) sc2mac_dat_data62_d1 : sc2mac_dat_data62_d2;
  assign _0171_ = sc2mac_dat_mask_d1[61] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:7081" *) sc2mac_dat_data61_d1 : sc2mac_dat_data61_d2;
  assign _0169_ = sc2mac_dat_mask_d1[60] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:7071" *) sc2mac_dat_data60_d1 : sc2mac_dat_data60_d2;
  assign _0165_ = sc2mac_dat_mask_d1[59] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:7061" *) sc2mac_dat_data59_d1 : sc2mac_dat_data59_d2;
  assign _0163_ = sc2mac_dat_mask_d1[58] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:7051" *) sc2mac_dat_data58_d1 : sc2mac_dat_data58_d2;
  assign _0161_ = sc2mac_dat_mask_d1[57] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:7041" *) sc2mac_dat_data57_d1 : sc2mac_dat_data57_d2;
  assign _0159_ = sc2mac_dat_mask_d1[56] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:7031" *) sc2mac_dat_data56_d1 : sc2mac_dat_data56_d2;
  assign _0157_ = sc2mac_dat_mask_d1[55] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:7021" *) sc2mac_dat_data55_d1 : sc2mac_dat_data55_d2;
  assign _0155_ = sc2mac_dat_mask_d1[54] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:7011" *) sc2mac_dat_data54_d1 : sc2mac_dat_data54_d2;
  assign _0153_ = sc2mac_dat_mask_d1[53] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:7001" *) sc2mac_dat_data53_d1 : sc2mac_dat_data53_d2;
  assign _0151_ = sc2mac_dat_mask_d1[52] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:6991" *) sc2mac_dat_data52_d1 : sc2mac_dat_data52_d2;
  assign _0149_ = sc2mac_dat_mask_d1[51] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:6981" *) sc2mac_dat_data51_d1 : sc2mac_dat_data51_d2;
  assign _0147_ = sc2mac_dat_mask_d1[50] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:6971" *) sc2mac_dat_data50_d1 : sc2mac_dat_data50_d2;
  assign _0143_ = sc2mac_dat_mask_d1[49] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:6961" *) sc2mac_dat_data49_d1 : sc2mac_dat_data49_d2;
  assign _0141_ = sc2mac_dat_mask_d1[48] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:6951" *) sc2mac_dat_data48_d1 : sc2mac_dat_data48_d2;
  assign _0139_ = sc2mac_dat_mask_d1[47] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:6941" *) sc2mac_dat_data47_d1 : sc2mac_dat_data47_d2;
  assign _0137_ = sc2mac_dat_mask_d1[46] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:6931" *) sc2mac_dat_data46_d1 : sc2mac_dat_data46_d2;
  assign _0135_ = sc2mac_dat_mask_d1[45] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:6921" *) sc2mac_dat_data45_d1 : sc2mac_dat_data45_d2;
  assign _0133_ = sc2mac_dat_mask_d1[44] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:6911" *) sc2mac_dat_data44_d1 : sc2mac_dat_data44_d2;
  assign _0131_ = sc2mac_dat_mask_d1[43] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:6901" *) sc2mac_dat_data43_d1 : sc2mac_dat_data43_d2;
  assign _0129_ = sc2mac_dat_mask_d1[42] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:6891" *) sc2mac_dat_data42_d1 : sc2mac_dat_data42_d2;
  assign _0127_ = sc2mac_dat_mask_d1[41] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:6881" *) sc2mac_dat_data41_d1 : sc2mac_dat_data41_d2;
  assign _0125_ = sc2mac_dat_mask_d1[40] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:6871" *) sc2mac_dat_data40_d1 : sc2mac_dat_data40_d2;
  assign _0121_ = sc2mac_dat_mask_d1[39] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:6861" *) sc2mac_dat_data39_d1 : sc2mac_dat_data39_d2;
  assign _0119_ = sc2mac_dat_mask_d1[38] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:6851" *) sc2mac_dat_data38_d1 : sc2mac_dat_data38_d2;
  assign _0117_ = sc2mac_dat_mask_d1[37] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:6841" *) sc2mac_dat_data37_d1 : sc2mac_dat_data37_d2;
  assign _0115_ = sc2mac_dat_mask_d1[36] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:6831" *) sc2mac_dat_data36_d1 : sc2mac_dat_data36_d2;
  assign _0113_ = sc2mac_dat_mask_d1[35] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:6821" *) sc2mac_dat_data35_d1 : sc2mac_dat_data35_d2;
  assign _0111_ = sc2mac_dat_mask_d1[34] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:6811" *) sc2mac_dat_data34_d1 : sc2mac_dat_data34_d2;
  assign _0109_ = sc2mac_dat_mask_d1[33] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:6801" *) sc2mac_dat_data33_d1 : sc2mac_dat_data33_d2;
  assign _0107_ = sc2mac_dat_mask_d1[32] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:6791" *) sc2mac_dat_data32_d1 : sc2mac_dat_data32_d2;
  assign _0105_ = sc2mac_dat_mask_d1[31] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:6781" *) sc2mac_dat_data31_d1 : sc2mac_dat_data31_d2;
  assign _0103_ = sc2mac_dat_mask_d1[30] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:6771" *) sc2mac_dat_data30_d1 : sc2mac_dat_data30_d2;
  assign _0099_ = sc2mac_dat_mask_d1[29] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:6761" *) sc2mac_dat_data29_d1 : sc2mac_dat_data29_d2;
  assign _0097_ = sc2mac_dat_mask_d1[28] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:6751" *) sc2mac_dat_data28_d1 : sc2mac_dat_data28_d2;
  assign _0095_ = sc2mac_dat_mask_d1[27] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:6741" *) sc2mac_dat_data27_d1 : sc2mac_dat_data27_d2;
  assign _0093_ = sc2mac_dat_mask_d1[26] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:6731" *) sc2mac_dat_data26_d1 : sc2mac_dat_data26_d2;
  assign _0091_ = sc2mac_dat_mask_d1[25] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:6721" *) sc2mac_dat_data25_d1 : sc2mac_dat_data25_d2;
  assign _0089_ = sc2mac_dat_mask_d1[24] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:6711" *) sc2mac_dat_data24_d1 : sc2mac_dat_data24_d2;
  assign _0087_ = sc2mac_dat_mask_d1[23] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:6701" *) sc2mac_dat_data23_d1 : sc2mac_dat_data23_d2;
  assign _0085_ = sc2mac_dat_mask_d1[22] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:6691" *) sc2mac_dat_data22_d1 : sc2mac_dat_data22_d2;
  assign _0083_ = sc2mac_dat_mask_d1[21] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:6681" *) sc2mac_dat_data21_d1 : sc2mac_dat_data21_d2;
  assign _0081_ = sc2mac_dat_mask_d1[20] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:6671" *) sc2mac_dat_data20_d1 : sc2mac_dat_data20_d2;
  assign _0077_ = sc2mac_dat_mask_d1[19] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:6661" *) sc2mac_dat_data19_d1 : sc2mac_dat_data19_d2;
  assign _0075_ = sc2mac_dat_mask_d1[18] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:6651" *) sc2mac_dat_data18_d1 : sc2mac_dat_data18_d2;
  assign _0073_ = sc2mac_dat_mask_d1[17] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:6641" *) sc2mac_dat_data17_d1 : sc2mac_dat_data17_d2;
  assign _0071_ = sc2mac_dat_mask_d1[16] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:6631" *) sc2mac_dat_data16_d1 : sc2mac_dat_data16_d2;
  assign _0069_ = sc2mac_dat_mask_d1[15] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:6621" *) sc2mac_dat_data15_d1 : sc2mac_dat_data15_d2;
  assign _0067_ = sc2mac_dat_mask_d1[14] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:6611" *) sc2mac_dat_data14_d1 : sc2mac_dat_data14_d2;
  assign _0065_ = sc2mac_dat_mask_d1[13] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:6601" *) sc2mac_dat_data13_d1 : sc2mac_dat_data13_d2;
  assign _0063_ = sc2mac_dat_mask_d1[12] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:6591" *) sc2mac_dat_data12_d1 : sc2mac_dat_data12_d2;
  assign _0045_ = sc2mac_dat_mask_d1[11] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:6581" *) sc2mac_dat_data11_d1 : sc2mac_dat_data11_d2;
  assign _0023_ = sc2mac_dat_mask_d1[10] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:6571" *) sc2mac_dat_data10_d1 : sc2mac_dat_data10_d2;
  assign _0255_ = sc2mac_dat_mask_d1[9] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:6561" *) sc2mac_dat_data9_d1 : sc2mac_dat_data9_d2;
  assign _0233_ = sc2mac_dat_mask_d1[8] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:6551" *) sc2mac_dat_data8_d1 : sc2mac_dat_data8_d2;
  assign _0211_ = sc2mac_dat_mask_d1[7] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:6541" *) sc2mac_dat_data7_d1 : sc2mac_dat_data7_d2;
  assign _0189_ = sc2mac_dat_mask_d1[6] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:6531" *) sc2mac_dat_data6_d1 : sc2mac_dat_data6_d2;
  assign _0167_ = sc2mac_dat_mask_d1[5] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:6521" *) sc2mac_dat_data5_d1 : sc2mac_dat_data5_d2;
  assign _0145_ = sc2mac_dat_mask_d1[4] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:6511" *) sc2mac_dat_data4_d1 : sc2mac_dat_data4_d2;
  assign _0123_ = sc2mac_dat_mask_d1[3] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:6501" *) sc2mac_dat_data3_d1 : sc2mac_dat_data3_d2;
  assign _0101_ = sc2mac_dat_mask_d1[2] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:6491" *) sc2mac_dat_data2_d1 : sc2mac_dat_data2_d2;
  assign _0079_ = sc2mac_dat_mask_d1[1] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:6481" *) sc2mac_dat_data1_d1 : sc2mac_dat_data1_d2;
  assign _0001_ = sc2mac_dat_mask_d1[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:6471" *) sc2mac_dat_data0_d1 : sc2mac_dat_data0_d2;
  assign _0257_ = _0523_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:6413" *) sc2mac_dat_mask_d1 : sc2mac_dat_mask_d2;
  assign _0259_ = _0523_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:6352" *) sc2mac_dat_pd_d1 : sc2mac_dat_pd_d2;
  assign _0321_ = sc2mac_wt_mask_d1[127] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:6332" *) sc2mac_wt_data127_d1 : sc2mac_wt_data127_d2;
  assign _0319_ = sc2mac_wt_mask_d1[126] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:6322" *) sc2mac_wt_data126_d1 : sc2mac_wt_data126_d2;
  assign _0317_ = sc2mac_wt_mask_d1[125] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:6312" *) sc2mac_wt_data125_d1 : sc2mac_wt_data125_d2;
  assign _0315_ = sc2mac_wt_mask_d1[124] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:6302" *) sc2mac_wt_data124_d1 : sc2mac_wt_data124_d2;
  assign _0313_ = sc2mac_wt_mask_d1[123] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:6292" *) sc2mac_wt_data123_d1 : sc2mac_wt_data123_d2;
  assign _0311_ = sc2mac_wt_mask_d1[122] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:6282" *) sc2mac_wt_data122_d1 : sc2mac_wt_data122_d2;
  assign _0309_ = sc2mac_wt_mask_d1[121] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:6272" *) sc2mac_wt_data121_d1 : sc2mac_wt_data121_d2;
  assign _0307_ = sc2mac_wt_mask_d1[120] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:6262" *) sc2mac_wt_data120_d1 : sc2mac_wt_data120_d2;
  assign _0303_ = sc2mac_wt_mask_d1[119] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:6252" *) sc2mac_wt_data119_d1 : sc2mac_wt_data119_d2;
  assign _0301_ = sc2mac_wt_mask_d1[118] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:6242" *) sc2mac_wt_data118_d1 : sc2mac_wt_data118_d2;
  assign _0299_ = sc2mac_wt_mask_d1[117] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:6232" *) sc2mac_wt_data117_d1 : sc2mac_wt_data117_d2;
  assign _0297_ = sc2mac_wt_mask_d1[116] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:6222" *) sc2mac_wt_data116_d1 : sc2mac_wt_data116_d2;
  assign _0295_ = sc2mac_wt_mask_d1[115] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:6212" *) sc2mac_wt_data115_d1 : sc2mac_wt_data115_d2;
  assign _0293_ = sc2mac_wt_mask_d1[114] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:6202" *) sc2mac_wt_data114_d1 : sc2mac_wt_data114_d2;
  assign _0291_ = sc2mac_wt_mask_d1[113] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:6192" *) sc2mac_wt_data113_d1 : sc2mac_wt_data113_d2;
  assign _0289_ = sc2mac_wt_mask_d1[112] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:6182" *) sc2mac_wt_data112_d1 : sc2mac_wt_data112_d2;
  assign _0287_ = sc2mac_wt_mask_d1[111] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:6172" *) sc2mac_wt_data111_d1 : sc2mac_wt_data111_d2;
  assign _0285_ = sc2mac_wt_mask_d1[110] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:6162" *) sc2mac_wt_data110_d1 : sc2mac_wt_data110_d2;
  assign _0281_ = sc2mac_wt_mask_d1[109] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:6152" *) sc2mac_wt_data109_d1 : sc2mac_wt_data109_d2;
  assign _0279_ = sc2mac_wt_mask_d1[108] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:6142" *) sc2mac_wt_data108_d1 : sc2mac_wt_data108_d2;
  assign _0277_ = sc2mac_wt_mask_d1[107] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:6132" *) sc2mac_wt_data107_d1 : sc2mac_wt_data107_d2;
  assign _0275_ = sc2mac_wt_mask_d1[106] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:6122" *) sc2mac_wt_data106_d1 : sc2mac_wt_data106_d2;
  assign _0273_ = sc2mac_wt_mask_d1[105] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:6112" *) sc2mac_wt_data105_d1 : sc2mac_wt_data105_d2;
  assign _0271_ = sc2mac_wt_mask_d1[104] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:6102" *) sc2mac_wt_data104_d1 : sc2mac_wt_data104_d2;
  assign _0269_ = sc2mac_wt_mask_d1[103] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:6092" *) sc2mac_wt_data103_d1 : sc2mac_wt_data103_d2;
  assign _0267_ = sc2mac_wt_mask_d1[102] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:6082" *) sc2mac_wt_data102_d1 : sc2mac_wt_data102_d2;
  assign _0265_ = sc2mac_wt_mask_d1[101] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:6072" *) sc2mac_wt_data101_d1 : sc2mac_wt_data101_d2;
  assign _0263_ = sc2mac_wt_mask_d1[100] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:6062" *) sc2mac_wt_data100_d1 : sc2mac_wt_data100_d2;
  assign _0513_ = sc2mac_wt_mask_d1[99] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:6052" *) sc2mac_wt_data99_d1 : sc2mac_wt_data99_d2;
  assign _0511_ = sc2mac_wt_mask_d1[98] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:6042" *) sc2mac_wt_data98_d1 : sc2mac_wt_data98_d2;
  assign _0509_ = sc2mac_wt_mask_d1[97] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:6032" *) sc2mac_wt_data97_d1 : sc2mac_wt_data97_d2;
  assign _0507_ = sc2mac_wt_mask_d1[96] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:6022" *) sc2mac_wt_data96_d1 : sc2mac_wt_data96_d2;
  assign _0505_ = sc2mac_wt_mask_d1[95] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:6012" *) sc2mac_wt_data95_d1 : sc2mac_wt_data95_d2;
  assign _0503_ = sc2mac_wt_mask_d1[94] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:6002" *) sc2mac_wt_data94_d1 : sc2mac_wt_data94_d2;
  assign _0501_ = sc2mac_wt_mask_d1[93] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:5992" *) sc2mac_wt_data93_d1 : sc2mac_wt_data93_d2;
  assign _0499_ = sc2mac_wt_mask_d1[92] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:5982" *) sc2mac_wt_data92_d1 : sc2mac_wt_data92_d2;
  assign _0497_ = sc2mac_wt_mask_d1[91] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:5972" *) sc2mac_wt_data91_d1 : sc2mac_wt_data91_d2;
  assign _0495_ = sc2mac_wt_mask_d1[90] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:5962" *) sc2mac_wt_data90_d1 : sc2mac_wt_data90_d2;
  assign _0491_ = sc2mac_wt_mask_d1[89] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:5952" *) sc2mac_wt_data89_d1 : sc2mac_wt_data89_d2;
  assign _0489_ = sc2mac_wt_mask_d1[88] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:5942" *) sc2mac_wt_data88_d1 : sc2mac_wt_data88_d2;
  assign _0487_ = sc2mac_wt_mask_d1[87] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:5932" *) sc2mac_wt_data87_d1 : sc2mac_wt_data87_d2;
  assign _0485_ = sc2mac_wt_mask_d1[86] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:5922" *) sc2mac_wt_data86_d1 : sc2mac_wt_data86_d2;
  assign _0483_ = sc2mac_wt_mask_d1[85] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:5912" *) sc2mac_wt_data85_d1 : sc2mac_wt_data85_d2;
  assign _0481_ = sc2mac_wt_mask_d1[84] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:5902" *) sc2mac_wt_data84_d1 : sc2mac_wt_data84_d2;
  assign _0479_ = sc2mac_wt_mask_d1[83] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:5892" *) sc2mac_wt_data83_d1 : sc2mac_wt_data83_d2;
  assign _0477_ = sc2mac_wt_mask_d1[82] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:5882" *) sc2mac_wt_data82_d1 : sc2mac_wt_data82_d2;
  assign _0475_ = sc2mac_wt_mask_d1[81] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:5872" *) sc2mac_wt_data81_d1 : sc2mac_wt_data81_d2;
  assign _0473_ = sc2mac_wt_mask_d1[80] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:5862" *) sc2mac_wt_data80_d1 : sc2mac_wt_data80_d2;
  assign _0469_ = sc2mac_wt_mask_d1[79] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:5852" *) sc2mac_wt_data79_d1 : sc2mac_wt_data79_d2;
  assign _0467_ = sc2mac_wt_mask_d1[78] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:5842" *) sc2mac_wt_data78_d1 : sc2mac_wt_data78_d2;
  assign _0465_ = sc2mac_wt_mask_d1[77] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:5832" *) sc2mac_wt_data77_d1 : sc2mac_wt_data77_d2;
  assign _0463_ = sc2mac_wt_mask_d1[76] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:5822" *) sc2mac_wt_data76_d1 : sc2mac_wt_data76_d2;
  assign _0461_ = sc2mac_wt_mask_d1[75] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:5812" *) sc2mac_wt_data75_d1 : sc2mac_wt_data75_d2;
  assign _0459_ = sc2mac_wt_mask_d1[74] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:5802" *) sc2mac_wt_data74_d1 : sc2mac_wt_data74_d2;
  assign _0457_ = sc2mac_wt_mask_d1[73] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:5792" *) sc2mac_wt_data73_d1 : sc2mac_wt_data73_d2;
  assign _0455_ = sc2mac_wt_mask_d1[72] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:5782" *) sc2mac_wt_data72_d1 : sc2mac_wt_data72_d2;
  assign _0453_ = sc2mac_wt_mask_d1[71] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:5772" *) sc2mac_wt_data71_d1 : sc2mac_wt_data71_d2;
  assign _0451_ = sc2mac_wt_mask_d1[70] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:5762" *) sc2mac_wt_data70_d1 : sc2mac_wt_data70_d2;
  assign _0447_ = sc2mac_wt_mask_d1[69] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:5752" *) sc2mac_wt_data69_d1 : sc2mac_wt_data69_d2;
  assign _0445_ = sc2mac_wt_mask_d1[68] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:5742" *) sc2mac_wt_data68_d1 : sc2mac_wt_data68_d2;
  assign _0443_ = sc2mac_wt_mask_d1[67] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:5732" *) sc2mac_wt_data67_d1 : sc2mac_wt_data67_d2;
  assign _0441_ = sc2mac_wt_mask_d1[66] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:5722" *) sc2mac_wt_data66_d1 : sc2mac_wt_data66_d2;
  assign _0439_ = sc2mac_wt_mask_d1[65] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:5712" *) sc2mac_wt_data65_d1 : sc2mac_wt_data65_d2;
  assign _0437_ = sc2mac_wt_mask_d1[64] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:5702" *) sc2mac_wt_data64_d1 : sc2mac_wt_data64_d2;
  assign _0435_ = sc2mac_wt_mask_d1[63] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:5692" *) sc2mac_wt_data63_d1 : sc2mac_wt_data63_d2;
  assign _0433_ = sc2mac_wt_mask_d1[62] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:5682" *) sc2mac_wt_data62_d1 : sc2mac_wt_data62_d2;
  assign _0431_ = sc2mac_wt_mask_d1[61] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:5672" *) sc2mac_wt_data61_d1 : sc2mac_wt_data61_d2;
  assign _0429_ = sc2mac_wt_mask_d1[60] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:5662" *) sc2mac_wt_data60_d1 : sc2mac_wt_data60_d2;
  assign _0425_ = sc2mac_wt_mask_d1[59] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:5652" *) sc2mac_wt_data59_d1 : sc2mac_wt_data59_d2;
  assign _0423_ = sc2mac_wt_mask_d1[58] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:5642" *) sc2mac_wt_data58_d1 : sc2mac_wt_data58_d2;
  assign _0421_ = sc2mac_wt_mask_d1[57] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:5632" *) sc2mac_wt_data57_d1 : sc2mac_wt_data57_d2;
  assign _0419_ = sc2mac_wt_mask_d1[56] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:5622" *) sc2mac_wt_data56_d1 : sc2mac_wt_data56_d2;
  assign _0417_ = sc2mac_wt_mask_d1[55] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:5612" *) sc2mac_wt_data55_d1 : sc2mac_wt_data55_d2;
  assign _0415_ = sc2mac_wt_mask_d1[54] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:5602" *) sc2mac_wt_data54_d1 : sc2mac_wt_data54_d2;
  assign _0413_ = sc2mac_wt_mask_d1[53] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:5592" *) sc2mac_wt_data53_d1 : sc2mac_wt_data53_d2;
  assign _0411_ = sc2mac_wt_mask_d1[52] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:5582" *) sc2mac_wt_data52_d1 : sc2mac_wt_data52_d2;
  assign _0409_ = sc2mac_wt_mask_d1[51] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:5572" *) sc2mac_wt_data51_d1 : sc2mac_wt_data51_d2;
  assign _0407_ = sc2mac_wt_mask_d1[50] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:5562" *) sc2mac_wt_data50_d1 : sc2mac_wt_data50_d2;
  assign _0403_ = sc2mac_wt_mask_d1[49] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:5552" *) sc2mac_wt_data49_d1 : sc2mac_wt_data49_d2;
  assign _0401_ = sc2mac_wt_mask_d1[48] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:5542" *) sc2mac_wt_data48_d1 : sc2mac_wt_data48_d2;
  assign _0399_ = sc2mac_wt_mask_d1[47] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:5532" *) sc2mac_wt_data47_d1 : sc2mac_wt_data47_d2;
  assign _0397_ = sc2mac_wt_mask_d1[46] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:5522" *) sc2mac_wt_data46_d1 : sc2mac_wt_data46_d2;
  assign _0395_ = sc2mac_wt_mask_d1[45] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:5512" *) sc2mac_wt_data45_d1 : sc2mac_wt_data45_d2;
  assign _0393_ = sc2mac_wt_mask_d1[44] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:5502" *) sc2mac_wt_data44_d1 : sc2mac_wt_data44_d2;
  assign _0391_ = sc2mac_wt_mask_d1[43] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:5492" *) sc2mac_wt_data43_d1 : sc2mac_wt_data43_d2;
  assign _0389_ = sc2mac_wt_mask_d1[42] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:5482" *) sc2mac_wt_data42_d1 : sc2mac_wt_data42_d2;
  assign _0387_ = sc2mac_wt_mask_d1[41] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:5472" *) sc2mac_wt_data41_d1 : sc2mac_wt_data41_d2;
  assign _0385_ = sc2mac_wt_mask_d1[40] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:5462" *) sc2mac_wt_data40_d1 : sc2mac_wt_data40_d2;
  assign _0381_ = sc2mac_wt_mask_d1[39] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:5452" *) sc2mac_wt_data39_d1 : sc2mac_wt_data39_d2;
  assign _0379_ = sc2mac_wt_mask_d1[38] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:5442" *) sc2mac_wt_data38_d1 : sc2mac_wt_data38_d2;
  assign _0377_ = sc2mac_wt_mask_d1[37] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:5432" *) sc2mac_wt_data37_d1 : sc2mac_wt_data37_d2;
  assign _0375_ = sc2mac_wt_mask_d1[36] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:5422" *) sc2mac_wt_data36_d1 : sc2mac_wt_data36_d2;
  assign _0373_ = sc2mac_wt_mask_d1[35] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:5412" *) sc2mac_wt_data35_d1 : sc2mac_wt_data35_d2;
  assign _0371_ = sc2mac_wt_mask_d1[34] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:5402" *) sc2mac_wt_data34_d1 : sc2mac_wt_data34_d2;
  assign _0369_ = sc2mac_wt_mask_d1[33] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:5392" *) sc2mac_wt_data33_d1 : sc2mac_wt_data33_d2;
  assign _0367_ = sc2mac_wt_mask_d1[32] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:5382" *) sc2mac_wt_data32_d1 : sc2mac_wt_data32_d2;
  assign _0365_ = sc2mac_wt_mask_d1[31] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:5372" *) sc2mac_wt_data31_d1 : sc2mac_wt_data31_d2;
  assign _0363_ = sc2mac_wt_mask_d1[30] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:5362" *) sc2mac_wt_data30_d1 : sc2mac_wt_data30_d2;
  assign _0359_ = sc2mac_wt_mask_d1[29] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:5352" *) sc2mac_wt_data29_d1 : sc2mac_wt_data29_d2;
  assign _0357_ = sc2mac_wt_mask_d1[28] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:5342" *) sc2mac_wt_data28_d1 : sc2mac_wt_data28_d2;
  assign _0355_ = sc2mac_wt_mask_d1[27] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:5332" *) sc2mac_wt_data27_d1 : sc2mac_wt_data27_d2;
  assign _0353_ = sc2mac_wt_mask_d1[26] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:5322" *) sc2mac_wt_data26_d1 : sc2mac_wt_data26_d2;
  assign _0351_ = sc2mac_wt_mask_d1[25] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:5312" *) sc2mac_wt_data25_d1 : sc2mac_wt_data25_d2;
  assign _0349_ = sc2mac_wt_mask_d1[24] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:5302" *) sc2mac_wt_data24_d1 : sc2mac_wt_data24_d2;
  assign _0347_ = sc2mac_wt_mask_d1[23] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:5292" *) sc2mac_wt_data23_d1 : sc2mac_wt_data23_d2;
  assign _0345_ = sc2mac_wt_mask_d1[22] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:5282" *) sc2mac_wt_data22_d1 : sc2mac_wt_data22_d2;
  assign _0343_ = sc2mac_wt_mask_d1[21] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:5272" *) sc2mac_wt_data21_d1 : sc2mac_wt_data21_d2;
  assign _0341_ = sc2mac_wt_mask_d1[20] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:5262" *) sc2mac_wt_data20_d1 : sc2mac_wt_data20_d2;
  assign _0337_ = sc2mac_wt_mask_d1[19] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:5252" *) sc2mac_wt_data19_d1 : sc2mac_wt_data19_d2;
  assign _0335_ = sc2mac_wt_mask_d1[18] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:5242" *) sc2mac_wt_data18_d1 : sc2mac_wt_data18_d2;
  assign _0333_ = sc2mac_wt_mask_d1[17] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:5232" *) sc2mac_wt_data17_d1 : sc2mac_wt_data17_d2;
  assign _0331_ = sc2mac_wt_mask_d1[16] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:5222" *) sc2mac_wt_data16_d1 : sc2mac_wt_data16_d2;
  assign _0329_ = sc2mac_wt_mask_d1[15] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:5212" *) sc2mac_wt_data15_d1 : sc2mac_wt_data15_d2;
  assign _0327_ = sc2mac_wt_mask_d1[14] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:5202" *) sc2mac_wt_data14_d1 : sc2mac_wt_data14_d2;
  assign _0325_ = sc2mac_wt_mask_d1[13] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:5192" *) sc2mac_wt_data13_d1 : sc2mac_wt_data13_d2;
  assign _0323_ = sc2mac_wt_mask_d1[12] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:5182" *) sc2mac_wt_data12_d1 : sc2mac_wt_data12_d2;
  assign _0305_ = sc2mac_wt_mask_d1[11] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:5172" *) sc2mac_wt_data11_d1 : sc2mac_wt_data11_d2;
  assign _0283_ = sc2mac_wt_mask_d1[10] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:5162" *) sc2mac_wt_data10_d1 : sc2mac_wt_data10_d2;
  assign _0515_ = sc2mac_wt_mask_d1[9] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:5152" *) sc2mac_wt_data9_d1 : sc2mac_wt_data9_d2;
  assign _0493_ = sc2mac_wt_mask_d1[8] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:5142" *) sc2mac_wt_data8_d1 : sc2mac_wt_data8_d2;
  assign _0471_ = sc2mac_wt_mask_d1[7] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:5132" *) sc2mac_wt_data7_d1 : sc2mac_wt_data7_d2;
  assign _0449_ = sc2mac_wt_mask_d1[6] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:5122" *) sc2mac_wt_data6_d1 : sc2mac_wt_data6_d2;
  assign _0427_ = sc2mac_wt_mask_d1[5] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:5112" *) sc2mac_wt_data5_d1 : sc2mac_wt_data5_d2;
  assign _0405_ = sc2mac_wt_mask_d1[4] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:5102" *) sc2mac_wt_data4_d1 : sc2mac_wt_data4_d2;
  assign _0383_ = sc2mac_wt_mask_d1[3] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:5092" *) sc2mac_wt_data3_d1 : sc2mac_wt_data3_d2;
  assign _0361_ = sc2mac_wt_mask_d1[2] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:5082" *) sc2mac_wt_data2_d1 : sc2mac_wt_data2_d2;
  assign _0339_ = sc2mac_wt_mask_d1[1] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:5072" *) sc2mac_wt_data1_d1 : sc2mac_wt_data1_d2;
  assign _0261_ = sc2mac_wt_mask_d1[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:5062" *) sc2mac_wt_data0_d1 : sc2mac_wt_data0_d2;
  assign _0517_ = _0522_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:5004" *) sc2mac_wt_mask_d1 : sc2mac_wt_mask_d2;
  assign _0519_ = _0522_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:4943" *) sc2mac_wt_sel_d1 : sc2mac_wt_sel_d2;
  assign _0060_ = sc2mac_dat_src_mask[127] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:4923" *) sc2mac_dat_src_data127 : sc2mac_dat_data127_d1;
  assign _0058_ = sc2mac_dat_src_mask[126] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:4913" *) sc2mac_dat_src_data126 : sc2mac_dat_data126_d1;
  assign _0056_ = sc2mac_dat_src_mask[125] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:4903" *) sc2mac_dat_src_data125 : sc2mac_dat_data125_d1;
  assign _0054_ = sc2mac_dat_src_mask[124] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:4893" *) sc2mac_dat_src_data124 : sc2mac_dat_data124_d1;
  assign _0052_ = sc2mac_dat_src_mask[123] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:4883" *) sc2mac_dat_src_data123 : sc2mac_dat_data123_d1;
  assign _0050_ = sc2mac_dat_src_mask[122] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:4873" *) sc2mac_dat_src_data122 : sc2mac_dat_data122_d1;
  assign _0048_ = sc2mac_dat_src_mask[121] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:4863" *) sc2mac_dat_src_data121 : sc2mac_dat_data121_d1;
  assign _0046_ = sc2mac_dat_src_mask[120] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:4853" *) sc2mac_dat_src_data120 : sc2mac_dat_data120_d1;
  assign _0042_ = sc2mac_dat_src_mask[119] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:4843" *) sc2mac_dat_src_data119 : sc2mac_dat_data119_d1;
  assign _0040_ = sc2mac_dat_src_mask[118] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:4833" *) sc2mac_dat_src_data118 : sc2mac_dat_data118_d1;
  assign _0038_ = sc2mac_dat_src_mask[117] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:4823" *) sc2mac_dat_src_data117 : sc2mac_dat_data117_d1;
  assign _0036_ = sc2mac_dat_src_mask[116] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:4813" *) sc2mac_dat_src_data116 : sc2mac_dat_data116_d1;
  assign _0034_ = sc2mac_dat_src_mask[115] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:4803" *) sc2mac_dat_src_data115 : sc2mac_dat_data115_d1;
  assign _0032_ = sc2mac_dat_src_mask[114] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:4793" *) sc2mac_dat_src_data114 : sc2mac_dat_data114_d1;
  assign _0030_ = sc2mac_dat_src_mask[113] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:4783" *) sc2mac_dat_src_data113 : sc2mac_dat_data113_d1;
  assign _0028_ = sc2mac_dat_src_mask[112] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:4773" *) sc2mac_dat_src_data112 : sc2mac_dat_data112_d1;
  assign _0026_ = sc2mac_dat_src_mask[111] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:4763" *) sc2mac_dat_src_data111 : sc2mac_dat_data111_d1;
  assign _0024_ = sc2mac_dat_src_mask[110] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:4753" *) sc2mac_dat_src_data110 : sc2mac_dat_data110_d1;
  assign _0020_ = sc2mac_dat_src_mask[109] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:4743" *) sc2mac_dat_src_data109 : sc2mac_dat_data109_d1;
  assign _0018_ = sc2mac_dat_src_mask[108] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:4733" *) sc2mac_dat_src_data108 : sc2mac_dat_data108_d1;
  assign _0016_ = sc2mac_dat_src_mask[107] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:4723" *) sc2mac_dat_src_data107 : sc2mac_dat_data107_d1;
  assign _0014_ = sc2mac_dat_src_mask[106] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:4713" *) sc2mac_dat_src_data106 : sc2mac_dat_data106_d1;
  assign _0012_ = sc2mac_dat_src_mask[105] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:4703" *) sc2mac_dat_src_data105 : sc2mac_dat_data105_d1;
  assign _0010_ = sc2mac_dat_src_mask[104] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:4693" *) sc2mac_dat_src_data104 : sc2mac_dat_data104_d1;
  assign _0008_ = sc2mac_dat_src_mask[103] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:4683" *) sc2mac_dat_src_data103 : sc2mac_dat_data103_d1;
  assign _0006_ = sc2mac_dat_src_mask[102] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:4673" *) sc2mac_dat_src_data102 : sc2mac_dat_data102_d1;
  assign _0004_ = sc2mac_dat_src_mask[101] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:4663" *) sc2mac_dat_src_data101 : sc2mac_dat_data101_d1;
  assign _0002_ = sc2mac_dat_src_mask[100] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:4653" *) sc2mac_dat_src_data100 : sc2mac_dat_data100_d1;
  assign _0252_ = sc2mac_dat_src_mask[99] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:4643" *) sc2mac_dat_src_data99 : sc2mac_dat_data99_d1;
  assign _0250_ = sc2mac_dat_src_mask[98] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:4633" *) sc2mac_dat_src_data98 : sc2mac_dat_data98_d1;
  assign _0248_ = sc2mac_dat_src_mask[97] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:4623" *) sc2mac_dat_src_data97 : sc2mac_dat_data97_d1;
  assign _0246_ = sc2mac_dat_src_mask[96] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:4613" *) sc2mac_dat_src_data96 : sc2mac_dat_data96_d1;
  assign _0244_ = sc2mac_dat_src_mask[95] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:4603" *) sc2mac_dat_src_data95 : sc2mac_dat_data95_d1;
  assign _0242_ = sc2mac_dat_src_mask[94] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:4593" *) sc2mac_dat_src_data94 : sc2mac_dat_data94_d1;
  assign _0240_ = sc2mac_dat_src_mask[93] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:4583" *) sc2mac_dat_src_data93 : sc2mac_dat_data93_d1;
  assign _0238_ = sc2mac_dat_src_mask[92] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:4573" *) sc2mac_dat_src_data92 : sc2mac_dat_data92_d1;
  assign _0236_ = sc2mac_dat_src_mask[91] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:4563" *) sc2mac_dat_src_data91 : sc2mac_dat_data91_d1;
  assign _0234_ = sc2mac_dat_src_mask[90] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:4553" *) sc2mac_dat_src_data90 : sc2mac_dat_data90_d1;
  assign _0230_ = sc2mac_dat_src_mask[89] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:4543" *) sc2mac_dat_src_data89 : sc2mac_dat_data89_d1;
  assign _0228_ = sc2mac_dat_src_mask[88] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:4533" *) sc2mac_dat_src_data88 : sc2mac_dat_data88_d1;
  assign _0226_ = sc2mac_dat_src_mask[87] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:4523" *) sc2mac_dat_src_data87 : sc2mac_dat_data87_d1;
  assign _0224_ = sc2mac_dat_src_mask[86] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:4513" *) sc2mac_dat_src_data86 : sc2mac_dat_data86_d1;
  assign _0222_ = sc2mac_dat_src_mask[85] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:4503" *) sc2mac_dat_src_data85 : sc2mac_dat_data85_d1;
  assign _0220_ = sc2mac_dat_src_mask[84] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:4493" *) sc2mac_dat_src_data84 : sc2mac_dat_data84_d1;
  assign _0218_ = sc2mac_dat_src_mask[83] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:4483" *) sc2mac_dat_src_data83 : sc2mac_dat_data83_d1;
  assign _0216_ = sc2mac_dat_src_mask[82] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:4473" *) sc2mac_dat_src_data82 : sc2mac_dat_data82_d1;
  assign _0214_ = sc2mac_dat_src_mask[81] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:4463" *) sc2mac_dat_src_data81 : sc2mac_dat_data81_d1;
  assign _0212_ = sc2mac_dat_src_mask[80] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:4453" *) sc2mac_dat_src_data80 : sc2mac_dat_data80_d1;
  assign _0208_ = sc2mac_dat_src_mask[79] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:4443" *) sc2mac_dat_src_data79 : sc2mac_dat_data79_d1;
  assign _0206_ = sc2mac_dat_src_mask[78] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:4433" *) sc2mac_dat_src_data78 : sc2mac_dat_data78_d1;
  assign _0204_ = sc2mac_dat_src_mask[77] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:4423" *) sc2mac_dat_src_data77 : sc2mac_dat_data77_d1;
  assign _0202_ = sc2mac_dat_src_mask[76] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:4413" *) sc2mac_dat_src_data76 : sc2mac_dat_data76_d1;
  assign _0200_ = sc2mac_dat_src_mask[75] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:4403" *) sc2mac_dat_src_data75 : sc2mac_dat_data75_d1;
  assign _0198_ = sc2mac_dat_src_mask[74] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:4393" *) sc2mac_dat_src_data74 : sc2mac_dat_data74_d1;
  assign _0196_ = sc2mac_dat_src_mask[73] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:4383" *) sc2mac_dat_src_data73 : sc2mac_dat_data73_d1;
  assign _0194_ = sc2mac_dat_src_mask[72] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:4373" *) sc2mac_dat_src_data72 : sc2mac_dat_data72_d1;
  assign _0192_ = sc2mac_dat_src_mask[71] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:4363" *) sc2mac_dat_src_data71 : sc2mac_dat_data71_d1;
  assign _0190_ = sc2mac_dat_src_mask[70] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:4353" *) sc2mac_dat_src_data70 : sc2mac_dat_data70_d1;
  assign _0186_ = sc2mac_dat_src_mask[69] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:4343" *) sc2mac_dat_src_data69 : sc2mac_dat_data69_d1;
  assign _0184_ = sc2mac_dat_src_mask[68] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:4333" *) sc2mac_dat_src_data68 : sc2mac_dat_data68_d1;
  assign _0182_ = sc2mac_dat_src_mask[67] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:4323" *) sc2mac_dat_src_data67 : sc2mac_dat_data67_d1;
  assign _0180_ = sc2mac_dat_src_mask[66] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:4313" *) sc2mac_dat_src_data66 : sc2mac_dat_data66_d1;
  assign _0178_ = sc2mac_dat_src_mask[65] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:4303" *) sc2mac_dat_src_data65 : sc2mac_dat_data65_d1;
  assign _0176_ = sc2mac_dat_src_mask[64] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:4293" *) sc2mac_dat_src_data64 : sc2mac_dat_data64_d1;
  assign _0174_ = sc2mac_dat_src_mask[63] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:4283" *) sc2mac_dat_src_data63 : sc2mac_dat_data63_d1;
  assign _0172_ = sc2mac_dat_src_mask[62] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:4273" *) sc2mac_dat_src_data62 : sc2mac_dat_data62_d1;
  assign _0170_ = sc2mac_dat_src_mask[61] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:4263" *) sc2mac_dat_src_data61 : sc2mac_dat_data61_d1;
  assign _0168_ = sc2mac_dat_src_mask[60] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:4253" *) sc2mac_dat_src_data60 : sc2mac_dat_data60_d1;
  assign _0164_ = sc2mac_dat_src_mask[59] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:4243" *) sc2mac_dat_src_data59 : sc2mac_dat_data59_d1;
  assign _0162_ = sc2mac_dat_src_mask[58] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:4233" *) sc2mac_dat_src_data58 : sc2mac_dat_data58_d1;
  assign _0160_ = sc2mac_dat_src_mask[57] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:4223" *) sc2mac_dat_src_data57 : sc2mac_dat_data57_d1;
  assign _0158_ = sc2mac_dat_src_mask[56] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:4213" *) sc2mac_dat_src_data56 : sc2mac_dat_data56_d1;
  assign _0156_ = sc2mac_dat_src_mask[55] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:4203" *) sc2mac_dat_src_data55 : sc2mac_dat_data55_d1;
  assign _0154_ = sc2mac_dat_src_mask[54] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:4193" *) sc2mac_dat_src_data54 : sc2mac_dat_data54_d1;
  assign _0152_ = sc2mac_dat_src_mask[53] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:4183" *) sc2mac_dat_src_data53 : sc2mac_dat_data53_d1;
  assign _0150_ = sc2mac_dat_src_mask[52] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:4173" *) sc2mac_dat_src_data52 : sc2mac_dat_data52_d1;
  assign _0148_ = sc2mac_dat_src_mask[51] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:4163" *) sc2mac_dat_src_data51 : sc2mac_dat_data51_d1;
  assign _0146_ = sc2mac_dat_src_mask[50] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:4153" *) sc2mac_dat_src_data50 : sc2mac_dat_data50_d1;
  assign _0142_ = sc2mac_dat_src_mask[49] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:4143" *) sc2mac_dat_src_data49 : sc2mac_dat_data49_d1;
  assign _0140_ = sc2mac_dat_src_mask[48] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:4133" *) sc2mac_dat_src_data48 : sc2mac_dat_data48_d1;
  assign _0138_ = sc2mac_dat_src_mask[47] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:4123" *) sc2mac_dat_src_data47 : sc2mac_dat_data47_d1;
  assign _0136_ = sc2mac_dat_src_mask[46] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:4113" *) sc2mac_dat_src_data46 : sc2mac_dat_data46_d1;
  assign _0134_ = sc2mac_dat_src_mask[45] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:4103" *) sc2mac_dat_src_data45 : sc2mac_dat_data45_d1;
  assign _0132_ = sc2mac_dat_src_mask[44] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:4093" *) sc2mac_dat_src_data44 : sc2mac_dat_data44_d1;
  assign _0130_ = sc2mac_dat_src_mask[43] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:4083" *) sc2mac_dat_src_data43 : sc2mac_dat_data43_d1;
  assign _0128_ = sc2mac_dat_src_mask[42] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:4073" *) sc2mac_dat_src_data42 : sc2mac_dat_data42_d1;
  assign _0126_ = sc2mac_dat_src_mask[41] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:4063" *) sc2mac_dat_src_data41 : sc2mac_dat_data41_d1;
  assign _0124_ = sc2mac_dat_src_mask[40] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:4053" *) sc2mac_dat_src_data40 : sc2mac_dat_data40_d1;
  assign _0120_ = sc2mac_dat_src_mask[39] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:4043" *) sc2mac_dat_src_data39 : sc2mac_dat_data39_d1;
  assign _0118_ = sc2mac_dat_src_mask[38] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:4033" *) sc2mac_dat_src_data38 : sc2mac_dat_data38_d1;
  assign _0116_ = sc2mac_dat_src_mask[37] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:4023" *) sc2mac_dat_src_data37 : sc2mac_dat_data37_d1;
  assign _0114_ = sc2mac_dat_src_mask[36] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:4013" *) sc2mac_dat_src_data36 : sc2mac_dat_data36_d1;
  assign _0112_ = sc2mac_dat_src_mask[35] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:4003" *) sc2mac_dat_src_data35 : sc2mac_dat_data35_d1;
  assign _0110_ = sc2mac_dat_src_mask[34] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:3993" *) sc2mac_dat_src_data34 : sc2mac_dat_data34_d1;
  assign _0108_ = sc2mac_dat_src_mask[33] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:3983" *) sc2mac_dat_src_data33 : sc2mac_dat_data33_d1;
  assign _0106_ = sc2mac_dat_src_mask[32] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:3973" *) sc2mac_dat_src_data32 : sc2mac_dat_data32_d1;
  assign _0104_ = sc2mac_dat_src_mask[31] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:3963" *) sc2mac_dat_src_data31 : sc2mac_dat_data31_d1;
  assign _0102_ = sc2mac_dat_src_mask[30] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:3953" *) sc2mac_dat_src_data30 : sc2mac_dat_data30_d1;
  assign _0098_ = sc2mac_dat_src_mask[29] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:3943" *) sc2mac_dat_src_data29 : sc2mac_dat_data29_d1;
  assign _0096_ = sc2mac_dat_src_mask[28] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:3933" *) sc2mac_dat_src_data28 : sc2mac_dat_data28_d1;
  assign _0094_ = sc2mac_dat_src_mask[27] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:3923" *) sc2mac_dat_src_data27 : sc2mac_dat_data27_d1;
  assign _0092_ = sc2mac_dat_src_mask[26] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:3913" *) sc2mac_dat_src_data26 : sc2mac_dat_data26_d1;
  assign _0090_ = sc2mac_dat_src_mask[25] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:3903" *) sc2mac_dat_src_data25 : sc2mac_dat_data25_d1;
  assign _0088_ = sc2mac_dat_src_mask[24] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:3893" *) sc2mac_dat_src_data24 : sc2mac_dat_data24_d1;
  assign _0086_ = sc2mac_dat_src_mask[23] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:3883" *) sc2mac_dat_src_data23 : sc2mac_dat_data23_d1;
  assign _0084_ = sc2mac_dat_src_mask[22] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:3873" *) sc2mac_dat_src_data22 : sc2mac_dat_data22_d1;
  assign _0082_ = sc2mac_dat_src_mask[21] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:3863" *) sc2mac_dat_src_data21 : sc2mac_dat_data21_d1;
  assign _0080_ = sc2mac_dat_src_mask[20] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:3853" *) sc2mac_dat_src_data20 : sc2mac_dat_data20_d1;
  assign _0076_ = sc2mac_dat_src_mask[19] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:3843" *) sc2mac_dat_src_data19 : sc2mac_dat_data19_d1;
  assign _0074_ = sc2mac_dat_src_mask[18] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:3833" *) sc2mac_dat_src_data18 : sc2mac_dat_data18_d1;
  assign _0072_ = sc2mac_dat_src_mask[17] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:3823" *) sc2mac_dat_src_data17 : sc2mac_dat_data17_d1;
  assign _0070_ = sc2mac_dat_src_mask[16] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:3813" *) sc2mac_dat_src_data16 : sc2mac_dat_data16_d1;
  assign _0068_ = sc2mac_dat_src_mask[15] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:3803" *) sc2mac_dat_src_data15 : sc2mac_dat_data15_d1;
  assign _0066_ = sc2mac_dat_src_mask[14] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:3793" *) sc2mac_dat_src_data14 : sc2mac_dat_data14_d1;
  assign _0064_ = sc2mac_dat_src_mask[13] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:3783" *) sc2mac_dat_src_data13 : sc2mac_dat_data13_d1;
  assign _0062_ = sc2mac_dat_src_mask[12] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:3773" *) sc2mac_dat_src_data12 : sc2mac_dat_data12_d1;
  assign _0044_ = sc2mac_dat_src_mask[11] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:3763" *) sc2mac_dat_src_data11 : sc2mac_dat_data11_d1;
  assign _0022_ = sc2mac_dat_src_mask[10] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:3753" *) sc2mac_dat_src_data10 : sc2mac_dat_data10_d1;
  assign _0254_ = sc2mac_dat_src_mask[9] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:3743" *) sc2mac_dat_src_data9 : sc2mac_dat_data9_d1;
  assign _0232_ = sc2mac_dat_src_mask[8] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:3733" *) sc2mac_dat_src_data8 : sc2mac_dat_data8_d1;
  assign _0210_ = sc2mac_dat_src_mask[7] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:3723" *) sc2mac_dat_src_data7 : sc2mac_dat_data7_d1;
  assign _0188_ = sc2mac_dat_src_mask[6] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:3713" *) sc2mac_dat_src_data6 : sc2mac_dat_data6_d1;
  assign _0166_ = sc2mac_dat_src_mask[5] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:3703" *) sc2mac_dat_src_data5 : sc2mac_dat_data5_d1;
  assign _0144_ = sc2mac_dat_src_mask[4] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:3693" *) sc2mac_dat_src_data4 : sc2mac_dat_data4_d1;
  assign _0122_ = sc2mac_dat_src_mask[3] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:3683" *) sc2mac_dat_src_data3 : sc2mac_dat_data3_d1;
  assign _0100_ = sc2mac_dat_src_mask[2] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:3673" *) sc2mac_dat_src_data2 : sc2mac_dat_data2_d1;
  assign _0078_ = sc2mac_dat_src_mask[1] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:3663" *) sc2mac_dat_src_data1 : sc2mac_dat_data1_d1;
  assign _0000_ = sc2mac_dat_src_mask[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:3653" *) sc2mac_dat_src_data0 : sc2mac_dat_data0_d1;
  assign _0256_ = _0521_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:3595" *) sc2mac_dat_src_mask : sc2mac_dat_mask_d1;
  assign _0258_ = _0521_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:3534" *) sc2mac_dat_src_pd : sc2mac_dat_pd_d1;
  assign _0320_ = sc2mac_wt_src_mask[127] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:3514" *) sc2mac_wt_src_data127 : sc2mac_wt_data127_d1;
  assign _0318_ = sc2mac_wt_src_mask[126] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:3504" *) sc2mac_wt_src_data126 : sc2mac_wt_data126_d1;
  assign _0316_ = sc2mac_wt_src_mask[125] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:3494" *) sc2mac_wt_src_data125 : sc2mac_wt_data125_d1;
  assign _0314_ = sc2mac_wt_src_mask[124] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:3484" *) sc2mac_wt_src_data124 : sc2mac_wt_data124_d1;
  assign _0312_ = sc2mac_wt_src_mask[123] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:3474" *) sc2mac_wt_src_data123 : sc2mac_wt_data123_d1;
  assign _0310_ = sc2mac_wt_src_mask[122] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:3464" *) sc2mac_wt_src_data122 : sc2mac_wt_data122_d1;
  assign _0308_ = sc2mac_wt_src_mask[121] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:3454" *) sc2mac_wt_src_data121 : sc2mac_wt_data121_d1;
  assign _0306_ = sc2mac_wt_src_mask[120] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:3444" *) sc2mac_wt_src_data120 : sc2mac_wt_data120_d1;
  assign _0302_ = sc2mac_wt_src_mask[119] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:3434" *) sc2mac_wt_src_data119 : sc2mac_wt_data119_d1;
  assign _0300_ = sc2mac_wt_src_mask[118] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:3424" *) sc2mac_wt_src_data118 : sc2mac_wt_data118_d1;
  assign _0298_ = sc2mac_wt_src_mask[117] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:3414" *) sc2mac_wt_src_data117 : sc2mac_wt_data117_d1;
  assign _0296_ = sc2mac_wt_src_mask[116] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:3404" *) sc2mac_wt_src_data116 : sc2mac_wt_data116_d1;
  assign _0294_ = sc2mac_wt_src_mask[115] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:3394" *) sc2mac_wt_src_data115 : sc2mac_wt_data115_d1;
  assign _0292_ = sc2mac_wt_src_mask[114] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:3384" *) sc2mac_wt_src_data114 : sc2mac_wt_data114_d1;
  assign _0290_ = sc2mac_wt_src_mask[113] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:3374" *) sc2mac_wt_src_data113 : sc2mac_wt_data113_d1;
  assign _0288_ = sc2mac_wt_src_mask[112] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:3364" *) sc2mac_wt_src_data112 : sc2mac_wt_data112_d1;
  assign _0286_ = sc2mac_wt_src_mask[111] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:3354" *) sc2mac_wt_src_data111 : sc2mac_wt_data111_d1;
  assign _0284_ = sc2mac_wt_src_mask[110] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:3344" *) sc2mac_wt_src_data110 : sc2mac_wt_data110_d1;
  assign _0280_ = sc2mac_wt_src_mask[109] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:3334" *) sc2mac_wt_src_data109 : sc2mac_wt_data109_d1;
  assign _0278_ = sc2mac_wt_src_mask[108] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:3324" *) sc2mac_wt_src_data108 : sc2mac_wt_data108_d1;
  assign _0276_ = sc2mac_wt_src_mask[107] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:3314" *) sc2mac_wt_src_data107 : sc2mac_wt_data107_d1;
  assign _0274_ = sc2mac_wt_src_mask[106] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:3304" *) sc2mac_wt_src_data106 : sc2mac_wt_data106_d1;
  assign _0272_ = sc2mac_wt_src_mask[105] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:3294" *) sc2mac_wt_src_data105 : sc2mac_wt_data105_d1;
  assign _0270_ = sc2mac_wt_src_mask[104] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:3284" *) sc2mac_wt_src_data104 : sc2mac_wt_data104_d1;
  assign _0268_ = sc2mac_wt_src_mask[103] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:3274" *) sc2mac_wt_src_data103 : sc2mac_wt_data103_d1;
  assign _0266_ = sc2mac_wt_src_mask[102] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:3264" *) sc2mac_wt_src_data102 : sc2mac_wt_data102_d1;
  assign _0264_ = sc2mac_wt_src_mask[101] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:3254" *) sc2mac_wt_src_data101 : sc2mac_wt_data101_d1;
  assign _0262_ = sc2mac_wt_src_mask[100] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:3244" *) sc2mac_wt_src_data100 : sc2mac_wt_data100_d1;
  assign _0512_ = sc2mac_wt_src_mask[99] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:3234" *) sc2mac_wt_src_data99 : sc2mac_wt_data99_d1;
  assign _0510_ = sc2mac_wt_src_mask[98] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:3224" *) sc2mac_wt_src_data98 : sc2mac_wt_data98_d1;
  assign _0508_ = sc2mac_wt_src_mask[97] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:3214" *) sc2mac_wt_src_data97 : sc2mac_wt_data97_d1;
  assign _0506_ = sc2mac_wt_src_mask[96] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:3204" *) sc2mac_wt_src_data96 : sc2mac_wt_data96_d1;
  assign _0504_ = sc2mac_wt_src_mask[95] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:3194" *) sc2mac_wt_src_data95 : sc2mac_wt_data95_d1;
  assign _0502_ = sc2mac_wt_src_mask[94] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:3184" *) sc2mac_wt_src_data94 : sc2mac_wt_data94_d1;
  assign _0500_ = sc2mac_wt_src_mask[93] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:3174" *) sc2mac_wt_src_data93 : sc2mac_wt_data93_d1;
  assign _0498_ = sc2mac_wt_src_mask[92] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:3164" *) sc2mac_wt_src_data92 : sc2mac_wt_data92_d1;
  assign _0496_ = sc2mac_wt_src_mask[91] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:3154" *) sc2mac_wt_src_data91 : sc2mac_wt_data91_d1;
  assign _0494_ = sc2mac_wt_src_mask[90] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:3144" *) sc2mac_wt_src_data90 : sc2mac_wt_data90_d1;
  assign _0490_ = sc2mac_wt_src_mask[89] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:3134" *) sc2mac_wt_src_data89 : sc2mac_wt_data89_d1;
  assign _0488_ = sc2mac_wt_src_mask[88] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:3124" *) sc2mac_wt_src_data88 : sc2mac_wt_data88_d1;
  assign _0486_ = sc2mac_wt_src_mask[87] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:3114" *) sc2mac_wt_src_data87 : sc2mac_wt_data87_d1;
  assign _0484_ = sc2mac_wt_src_mask[86] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:3104" *) sc2mac_wt_src_data86 : sc2mac_wt_data86_d1;
  assign _0482_ = sc2mac_wt_src_mask[85] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:3094" *) sc2mac_wt_src_data85 : sc2mac_wt_data85_d1;
  assign _0480_ = sc2mac_wt_src_mask[84] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:3084" *) sc2mac_wt_src_data84 : sc2mac_wt_data84_d1;
  assign _0478_ = sc2mac_wt_src_mask[83] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:3074" *) sc2mac_wt_src_data83 : sc2mac_wt_data83_d1;
  assign _0476_ = sc2mac_wt_src_mask[82] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:3064" *) sc2mac_wt_src_data82 : sc2mac_wt_data82_d1;
  assign _0474_ = sc2mac_wt_src_mask[81] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:3054" *) sc2mac_wt_src_data81 : sc2mac_wt_data81_d1;
  assign _0472_ = sc2mac_wt_src_mask[80] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:3044" *) sc2mac_wt_src_data80 : sc2mac_wt_data80_d1;
  assign _0468_ = sc2mac_wt_src_mask[79] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:3034" *) sc2mac_wt_src_data79 : sc2mac_wt_data79_d1;
  assign _0466_ = sc2mac_wt_src_mask[78] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:3024" *) sc2mac_wt_src_data78 : sc2mac_wt_data78_d1;
  assign _0464_ = sc2mac_wt_src_mask[77] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:3014" *) sc2mac_wt_src_data77 : sc2mac_wt_data77_d1;
  assign _0462_ = sc2mac_wt_src_mask[76] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:3004" *) sc2mac_wt_src_data76 : sc2mac_wt_data76_d1;
  assign _0460_ = sc2mac_wt_src_mask[75] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:2994" *) sc2mac_wt_src_data75 : sc2mac_wt_data75_d1;
  assign _0458_ = sc2mac_wt_src_mask[74] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:2984" *) sc2mac_wt_src_data74 : sc2mac_wt_data74_d1;
  assign _0456_ = sc2mac_wt_src_mask[73] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:2974" *) sc2mac_wt_src_data73 : sc2mac_wt_data73_d1;
  assign _0454_ = sc2mac_wt_src_mask[72] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:2964" *) sc2mac_wt_src_data72 : sc2mac_wt_data72_d1;
  assign _0452_ = sc2mac_wt_src_mask[71] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:2954" *) sc2mac_wt_src_data71 : sc2mac_wt_data71_d1;
  assign _0450_ = sc2mac_wt_src_mask[70] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:2944" *) sc2mac_wt_src_data70 : sc2mac_wt_data70_d1;
  assign _0446_ = sc2mac_wt_src_mask[69] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:2934" *) sc2mac_wt_src_data69 : sc2mac_wt_data69_d1;
  assign _0444_ = sc2mac_wt_src_mask[68] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:2924" *) sc2mac_wt_src_data68 : sc2mac_wt_data68_d1;
  assign _0442_ = sc2mac_wt_src_mask[67] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:2914" *) sc2mac_wt_src_data67 : sc2mac_wt_data67_d1;
  assign _0440_ = sc2mac_wt_src_mask[66] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:2904" *) sc2mac_wt_src_data66 : sc2mac_wt_data66_d1;
  assign _0438_ = sc2mac_wt_src_mask[65] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:2894" *) sc2mac_wt_src_data65 : sc2mac_wt_data65_d1;
  assign _0436_ = sc2mac_wt_src_mask[64] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:2884" *) sc2mac_wt_src_data64 : sc2mac_wt_data64_d1;
  assign _0434_ = sc2mac_wt_src_mask[63] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:2874" *) sc2mac_wt_src_data63 : sc2mac_wt_data63_d1;
  assign _0432_ = sc2mac_wt_src_mask[62] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:2864" *) sc2mac_wt_src_data62 : sc2mac_wt_data62_d1;
  assign _0430_ = sc2mac_wt_src_mask[61] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:2854" *) sc2mac_wt_src_data61 : sc2mac_wt_data61_d1;
  assign _0428_ = sc2mac_wt_src_mask[60] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:2844" *) sc2mac_wt_src_data60 : sc2mac_wt_data60_d1;
  assign _0424_ = sc2mac_wt_src_mask[59] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:2834" *) sc2mac_wt_src_data59 : sc2mac_wt_data59_d1;
  assign _0422_ = sc2mac_wt_src_mask[58] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:2824" *) sc2mac_wt_src_data58 : sc2mac_wt_data58_d1;
  assign _0420_ = sc2mac_wt_src_mask[57] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:2814" *) sc2mac_wt_src_data57 : sc2mac_wt_data57_d1;
  assign _0418_ = sc2mac_wt_src_mask[56] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:2804" *) sc2mac_wt_src_data56 : sc2mac_wt_data56_d1;
  assign _0416_ = sc2mac_wt_src_mask[55] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:2794" *) sc2mac_wt_src_data55 : sc2mac_wt_data55_d1;
  assign _0414_ = sc2mac_wt_src_mask[54] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:2784" *) sc2mac_wt_src_data54 : sc2mac_wt_data54_d1;
  assign _0412_ = sc2mac_wt_src_mask[53] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:2774" *) sc2mac_wt_src_data53 : sc2mac_wt_data53_d1;
  assign _0410_ = sc2mac_wt_src_mask[52] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:2764" *) sc2mac_wt_src_data52 : sc2mac_wt_data52_d1;
  assign _0408_ = sc2mac_wt_src_mask[51] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:2754" *) sc2mac_wt_src_data51 : sc2mac_wt_data51_d1;
  assign _0406_ = sc2mac_wt_src_mask[50] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:2744" *) sc2mac_wt_src_data50 : sc2mac_wt_data50_d1;
  assign _0402_ = sc2mac_wt_src_mask[49] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:2734" *) sc2mac_wt_src_data49 : sc2mac_wt_data49_d1;
  assign _0400_ = sc2mac_wt_src_mask[48] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:2724" *) sc2mac_wt_src_data48 : sc2mac_wt_data48_d1;
  assign _0398_ = sc2mac_wt_src_mask[47] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:2714" *) sc2mac_wt_src_data47 : sc2mac_wt_data47_d1;
  assign _0396_ = sc2mac_wt_src_mask[46] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:2704" *) sc2mac_wt_src_data46 : sc2mac_wt_data46_d1;
  assign _0394_ = sc2mac_wt_src_mask[45] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:2694" *) sc2mac_wt_src_data45 : sc2mac_wt_data45_d1;
  assign _0392_ = sc2mac_wt_src_mask[44] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:2684" *) sc2mac_wt_src_data44 : sc2mac_wt_data44_d1;
  assign _0390_ = sc2mac_wt_src_mask[43] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:2674" *) sc2mac_wt_src_data43 : sc2mac_wt_data43_d1;
  assign _0388_ = sc2mac_wt_src_mask[42] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:2664" *) sc2mac_wt_src_data42 : sc2mac_wt_data42_d1;
  assign _0386_ = sc2mac_wt_src_mask[41] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:2654" *) sc2mac_wt_src_data41 : sc2mac_wt_data41_d1;
  assign _0384_ = sc2mac_wt_src_mask[40] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:2644" *) sc2mac_wt_src_data40 : sc2mac_wt_data40_d1;
  assign _0380_ = sc2mac_wt_src_mask[39] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:2634" *) sc2mac_wt_src_data39 : sc2mac_wt_data39_d1;
  assign _0378_ = sc2mac_wt_src_mask[38] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:2624" *) sc2mac_wt_src_data38 : sc2mac_wt_data38_d1;
  assign _0376_ = sc2mac_wt_src_mask[37] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:2614" *) sc2mac_wt_src_data37 : sc2mac_wt_data37_d1;
  assign _0374_ = sc2mac_wt_src_mask[36] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:2604" *) sc2mac_wt_src_data36 : sc2mac_wt_data36_d1;
  assign _0372_ = sc2mac_wt_src_mask[35] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:2594" *) sc2mac_wt_src_data35 : sc2mac_wt_data35_d1;
  assign _0370_ = sc2mac_wt_src_mask[34] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:2584" *) sc2mac_wt_src_data34 : sc2mac_wt_data34_d1;
  assign _0368_ = sc2mac_wt_src_mask[33] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:2574" *) sc2mac_wt_src_data33 : sc2mac_wt_data33_d1;
  assign _0366_ = sc2mac_wt_src_mask[32] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:2564" *) sc2mac_wt_src_data32 : sc2mac_wt_data32_d1;
  assign _0364_ = sc2mac_wt_src_mask[31] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:2554" *) sc2mac_wt_src_data31 : sc2mac_wt_data31_d1;
  assign _0362_ = sc2mac_wt_src_mask[30] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:2544" *) sc2mac_wt_src_data30 : sc2mac_wt_data30_d1;
  assign _0358_ = sc2mac_wt_src_mask[29] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:2534" *) sc2mac_wt_src_data29 : sc2mac_wt_data29_d1;
  assign _0356_ = sc2mac_wt_src_mask[28] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:2524" *) sc2mac_wt_src_data28 : sc2mac_wt_data28_d1;
  assign _0354_ = sc2mac_wt_src_mask[27] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:2514" *) sc2mac_wt_src_data27 : sc2mac_wt_data27_d1;
  assign _0352_ = sc2mac_wt_src_mask[26] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:2504" *) sc2mac_wt_src_data26 : sc2mac_wt_data26_d1;
  assign _0350_ = sc2mac_wt_src_mask[25] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:2494" *) sc2mac_wt_src_data25 : sc2mac_wt_data25_d1;
  assign _0348_ = sc2mac_wt_src_mask[24] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:2484" *) sc2mac_wt_src_data24 : sc2mac_wt_data24_d1;
  assign _0346_ = sc2mac_wt_src_mask[23] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:2474" *) sc2mac_wt_src_data23 : sc2mac_wt_data23_d1;
  assign _0344_ = sc2mac_wt_src_mask[22] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:2464" *) sc2mac_wt_src_data22 : sc2mac_wt_data22_d1;
  assign _0342_ = sc2mac_wt_src_mask[21] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:2454" *) sc2mac_wt_src_data21 : sc2mac_wt_data21_d1;
  assign _0340_ = sc2mac_wt_src_mask[20] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:2444" *) sc2mac_wt_src_data20 : sc2mac_wt_data20_d1;
  assign _0336_ = sc2mac_wt_src_mask[19] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:2434" *) sc2mac_wt_src_data19 : sc2mac_wt_data19_d1;
  assign _0334_ = sc2mac_wt_src_mask[18] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:2424" *) sc2mac_wt_src_data18 : sc2mac_wt_data18_d1;
  assign _0332_ = sc2mac_wt_src_mask[17] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:2414" *) sc2mac_wt_src_data17 : sc2mac_wt_data17_d1;
  assign _0330_ = sc2mac_wt_src_mask[16] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:2404" *) sc2mac_wt_src_data16 : sc2mac_wt_data16_d1;
  assign _0328_ = sc2mac_wt_src_mask[15] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:2394" *) sc2mac_wt_src_data15 : sc2mac_wt_data15_d1;
  assign _0326_ = sc2mac_wt_src_mask[14] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:2384" *) sc2mac_wt_src_data14 : sc2mac_wt_data14_d1;
  assign _0324_ = sc2mac_wt_src_mask[13] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:2374" *) sc2mac_wt_src_data13 : sc2mac_wt_data13_d1;
  assign _0322_ = sc2mac_wt_src_mask[12] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:2364" *) sc2mac_wt_src_data12 : sc2mac_wt_data12_d1;
  assign _0304_ = sc2mac_wt_src_mask[11] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:2354" *) sc2mac_wt_src_data11 : sc2mac_wt_data11_d1;
  assign _0282_ = sc2mac_wt_src_mask[10] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:2344" *) sc2mac_wt_src_data10 : sc2mac_wt_data10_d1;
  assign _0514_ = sc2mac_wt_src_mask[9] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:2334" *) sc2mac_wt_src_data9 : sc2mac_wt_data9_d1;
  assign _0492_ = sc2mac_wt_src_mask[8] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:2324" *) sc2mac_wt_src_data8 : sc2mac_wt_data8_d1;
  assign _0470_ = sc2mac_wt_src_mask[7] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:2314" *) sc2mac_wt_src_data7 : sc2mac_wt_data7_d1;
  assign _0448_ = sc2mac_wt_src_mask[6] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:2304" *) sc2mac_wt_src_data6 : sc2mac_wt_data6_d1;
  assign _0426_ = sc2mac_wt_src_mask[5] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:2294" *) sc2mac_wt_src_data5 : sc2mac_wt_data5_d1;
  assign _0404_ = sc2mac_wt_src_mask[4] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:2284" *) sc2mac_wt_src_data4 : sc2mac_wt_data4_d1;
  assign _0382_ = sc2mac_wt_src_mask[3] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:2274" *) sc2mac_wt_src_data3 : sc2mac_wt_data3_d1;
  assign _0360_ = sc2mac_wt_src_mask[2] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:2264" *) sc2mac_wt_src_data2 : sc2mac_wt_data2_d1;
  assign _0338_ = sc2mac_wt_src_mask[1] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:2254" *) sc2mac_wt_src_data1 : sc2mac_wt_data1_d1;
  assign _0260_ = sc2mac_wt_src_mask[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:2244" *) sc2mac_wt_src_data0 : sc2mac_wt_data0_d1;
  assign _0516_ = _0520_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:2186" *) sc2mac_wt_src_mask : sc2mac_wt_mask_d1;
  assign _0518_ = _0520_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_a.v:2125" *) sc2mac_wt_src_sel : sc2mac_wt_sel_d1;
  assign sc2mac_dat_data0_d0 = sc2mac_dat_src_data0;
  assign sc2mac_dat_data100_d0 = sc2mac_dat_src_data100;
  assign sc2mac_dat_data101_d0 = sc2mac_dat_src_data101;
  assign sc2mac_dat_data102_d0 = sc2mac_dat_src_data102;
  assign sc2mac_dat_data103_d0 = sc2mac_dat_src_data103;
  assign sc2mac_dat_data104_d0 = sc2mac_dat_src_data104;
  assign sc2mac_dat_data105_d0 = sc2mac_dat_src_data105;
  assign sc2mac_dat_data106_d0 = sc2mac_dat_src_data106;
  assign sc2mac_dat_data107_d0 = sc2mac_dat_src_data107;
  assign sc2mac_dat_data108_d0 = sc2mac_dat_src_data108;
  assign sc2mac_dat_data109_d0 = sc2mac_dat_src_data109;
  assign sc2mac_dat_data10_d0 = sc2mac_dat_src_data10;
  assign sc2mac_dat_data110_d0 = sc2mac_dat_src_data110;
  assign sc2mac_dat_data111_d0 = sc2mac_dat_src_data111;
  assign sc2mac_dat_data112_d0 = sc2mac_dat_src_data112;
  assign sc2mac_dat_data113_d0 = sc2mac_dat_src_data113;
  assign sc2mac_dat_data114_d0 = sc2mac_dat_src_data114;
  assign sc2mac_dat_data115_d0 = sc2mac_dat_src_data115;
  assign sc2mac_dat_data116_d0 = sc2mac_dat_src_data116;
  assign sc2mac_dat_data117_d0 = sc2mac_dat_src_data117;
  assign sc2mac_dat_data118_d0 = sc2mac_dat_src_data118;
  assign sc2mac_dat_data119_d0 = sc2mac_dat_src_data119;
  assign sc2mac_dat_data11_d0 = sc2mac_dat_src_data11;
  assign sc2mac_dat_data120_d0 = sc2mac_dat_src_data120;
  assign sc2mac_dat_data121_d0 = sc2mac_dat_src_data121;
  assign sc2mac_dat_data122_d0 = sc2mac_dat_src_data122;
  assign sc2mac_dat_data123_d0 = sc2mac_dat_src_data123;
  assign sc2mac_dat_data124_d0 = sc2mac_dat_src_data124;
  assign sc2mac_dat_data125_d0 = sc2mac_dat_src_data125;
  assign sc2mac_dat_data126_d0 = sc2mac_dat_src_data126;
  assign sc2mac_dat_data127_d0 = sc2mac_dat_src_data127;
  assign sc2mac_dat_data12_d0 = sc2mac_dat_src_data12;
  assign sc2mac_dat_data13_d0 = sc2mac_dat_src_data13;
  assign sc2mac_dat_data14_d0 = sc2mac_dat_src_data14;
  assign sc2mac_dat_data15_d0 = sc2mac_dat_src_data15;
  assign sc2mac_dat_data16_d0 = sc2mac_dat_src_data16;
  assign sc2mac_dat_data17_d0 = sc2mac_dat_src_data17;
  assign sc2mac_dat_data18_d0 = sc2mac_dat_src_data18;
  assign sc2mac_dat_data19_d0 = sc2mac_dat_src_data19;
  assign sc2mac_dat_data1_d0 = sc2mac_dat_src_data1;
  assign sc2mac_dat_data20_d0 = sc2mac_dat_src_data20;
  assign sc2mac_dat_data21_d0 = sc2mac_dat_src_data21;
  assign sc2mac_dat_data22_d0 = sc2mac_dat_src_data22;
  assign sc2mac_dat_data23_d0 = sc2mac_dat_src_data23;
  assign sc2mac_dat_data24_d0 = sc2mac_dat_src_data24;
  assign sc2mac_dat_data25_d0 = sc2mac_dat_src_data25;
  assign sc2mac_dat_data26_d0 = sc2mac_dat_src_data26;
  assign sc2mac_dat_data27_d0 = sc2mac_dat_src_data27;
  assign sc2mac_dat_data28_d0 = sc2mac_dat_src_data28;
  assign sc2mac_dat_data29_d0 = sc2mac_dat_src_data29;
  assign sc2mac_dat_data2_d0 = sc2mac_dat_src_data2;
  assign sc2mac_dat_data30_d0 = sc2mac_dat_src_data30;
  assign sc2mac_dat_data31_d0 = sc2mac_dat_src_data31;
  assign sc2mac_dat_data32_d0 = sc2mac_dat_src_data32;
  assign sc2mac_dat_data33_d0 = sc2mac_dat_src_data33;
  assign sc2mac_dat_data34_d0 = sc2mac_dat_src_data34;
  assign sc2mac_dat_data35_d0 = sc2mac_dat_src_data35;
  assign sc2mac_dat_data36_d0 = sc2mac_dat_src_data36;
  assign sc2mac_dat_data37_d0 = sc2mac_dat_src_data37;
  assign sc2mac_dat_data38_d0 = sc2mac_dat_src_data38;
  assign sc2mac_dat_data39_d0 = sc2mac_dat_src_data39;
  assign sc2mac_dat_data3_d0 = sc2mac_dat_src_data3;
  assign sc2mac_dat_data40_d0 = sc2mac_dat_src_data40;
  assign sc2mac_dat_data41_d0 = sc2mac_dat_src_data41;
  assign sc2mac_dat_data42_d0 = sc2mac_dat_src_data42;
  assign sc2mac_dat_data43_d0 = sc2mac_dat_src_data43;
  assign sc2mac_dat_data44_d0 = sc2mac_dat_src_data44;
  assign sc2mac_dat_data45_d0 = sc2mac_dat_src_data45;
  assign sc2mac_dat_data46_d0 = sc2mac_dat_src_data46;
  assign sc2mac_dat_data47_d0 = sc2mac_dat_src_data47;
  assign sc2mac_dat_data48_d0 = sc2mac_dat_src_data48;
  assign sc2mac_dat_data49_d0 = sc2mac_dat_src_data49;
  assign sc2mac_dat_data4_d0 = sc2mac_dat_src_data4;
  assign sc2mac_dat_data50_d0 = sc2mac_dat_src_data50;
  assign sc2mac_dat_data51_d0 = sc2mac_dat_src_data51;
  assign sc2mac_dat_data52_d0 = sc2mac_dat_src_data52;
  assign sc2mac_dat_data53_d0 = sc2mac_dat_src_data53;
  assign sc2mac_dat_data54_d0 = sc2mac_dat_src_data54;
  assign sc2mac_dat_data55_d0 = sc2mac_dat_src_data55;
  assign sc2mac_dat_data56_d0 = sc2mac_dat_src_data56;
  assign sc2mac_dat_data57_d0 = sc2mac_dat_src_data57;
  assign sc2mac_dat_data58_d0 = sc2mac_dat_src_data58;
  assign sc2mac_dat_data59_d0 = sc2mac_dat_src_data59;
  assign sc2mac_dat_data5_d0 = sc2mac_dat_src_data5;
  assign sc2mac_dat_data60_d0 = sc2mac_dat_src_data60;
  assign sc2mac_dat_data61_d0 = sc2mac_dat_src_data61;
  assign sc2mac_dat_data62_d0 = sc2mac_dat_src_data62;
  assign sc2mac_dat_data63_d0 = sc2mac_dat_src_data63;
  assign sc2mac_dat_data64_d0 = sc2mac_dat_src_data64;
  assign sc2mac_dat_data65_d0 = sc2mac_dat_src_data65;
  assign sc2mac_dat_data66_d0 = sc2mac_dat_src_data66;
  assign sc2mac_dat_data67_d0 = sc2mac_dat_src_data67;
  assign sc2mac_dat_data68_d0 = sc2mac_dat_src_data68;
  assign sc2mac_dat_data69_d0 = sc2mac_dat_src_data69;
  assign sc2mac_dat_data6_d0 = sc2mac_dat_src_data6;
  assign sc2mac_dat_data70_d0 = sc2mac_dat_src_data70;
  assign sc2mac_dat_data71_d0 = sc2mac_dat_src_data71;
  assign sc2mac_dat_data72_d0 = sc2mac_dat_src_data72;
  assign sc2mac_dat_data73_d0 = sc2mac_dat_src_data73;
  assign sc2mac_dat_data74_d0 = sc2mac_dat_src_data74;
  assign sc2mac_dat_data75_d0 = sc2mac_dat_src_data75;
  assign sc2mac_dat_data76_d0 = sc2mac_dat_src_data76;
  assign sc2mac_dat_data77_d0 = sc2mac_dat_src_data77;
  assign sc2mac_dat_data78_d0 = sc2mac_dat_src_data78;
  assign sc2mac_dat_data79_d0 = sc2mac_dat_src_data79;
  assign sc2mac_dat_data7_d0 = sc2mac_dat_src_data7;
  assign sc2mac_dat_data80_d0 = sc2mac_dat_src_data80;
  assign sc2mac_dat_data81_d0 = sc2mac_dat_src_data81;
  assign sc2mac_dat_data82_d0 = sc2mac_dat_src_data82;
  assign sc2mac_dat_data83_d0 = sc2mac_dat_src_data83;
  assign sc2mac_dat_data84_d0 = sc2mac_dat_src_data84;
  assign sc2mac_dat_data85_d0 = sc2mac_dat_src_data85;
  assign sc2mac_dat_data86_d0 = sc2mac_dat_src_data86;
  assign sc2mac_dat_data87_d0 = sc2mac_dat_src_data87;
  assign sc2mac_dat_data88_d0 = sc2mac_dat_src_data88;
  assign sc2mac_dat_data89_d0 = sc2mac_dat_src_data89;
  assign sc2mac_dat_data8_d0 = sc2mac_dat_src_data8;
  assign sc2mac_dat_data90_d0 = sc2mac_dat_src_data90;
  assign sc2mac_dat_data91_d0 = sc2mac_dat_src_data91;
  assign sc2mac_dat_data92_d0 = sc2mac_dat_src_data92;
  assign sc2mac_dat_data93_d0 = sc2mac_dat_src_data93;
  assign sc2mac_dat_data94_d0 = sc2mac_dat_src_data94;
  assign sc2mac_dat_data95_d0 = sc2mac_dat_src_data95;
  assign sc2mac_dat_data96_d0 = sc2mac_dat_src_data96;
  assign sc2mac_dat_data97_d0 = sc2mac_dat_src_data97;
  assign sc2mac_dat_data98_d0 = sc2mac_dat_src_data98;
  assign sc2mac_dat_data99_d0 = sc2mac_dat_src_data99;
  assign sc2mac_dat_data9_d0 = sc2mac_dat_src_data9;
  assign sc2mac_dat_dst_data0 = sc2mac_dat_data0_d2;
  assign sc2mac_dat_dst_data1 = sc2mac_dat_data1_d2;
  assign sc2mac_dat_dst_data10 = sc2mac_dat_data10_d2;
  assign sc2mac_dat_dst_data100 = sc2mac_dat_data100_d2;
  assign sc2mac_dat_dst_data101 = sc2mac_dat_data101_d2;
  assign sc2mac_dat_dst_data102 = sc2mac_dat_data102_d2;
  assign sc2mac_dat_dst_data103 = sc2mac_dat_data103_d2;
  assign sc2mac_dat_dst_data104 = sc2mac_dat_data104_d2;
  assign sc2mac_dat_dst_data105 = sc2mac_dat_data105_d2;
  assign sc2mac_dat_dst_data106 = sc2mac_dat_data106_d2;
  assign sc2mac_dat_dst_data107 = sc2mac_dat_data107_d2;
  assign sc2mac_dat_dst_data108 = sc2mac_dat_data108_d2;
  assign sc2mac_dat_dst_data109 = sc2mac_dat_data109_d2;
  assign sc2mac_dat_dst_data11 = sc2mac_dat_data11_d2;
  assign sc2mac_dat_dst_data110 = sc2mac_dat_data110_d2;
  assign sc2mac_dat_dst_data111 = sc2mac_dat_data111_d2;
  assign sc2mac_dat_dst_data112 = sc2mac_dat_data112_d2;
  assign sc2mac_dat_dst_data113 = sc2mac_dat_data113_d2;
  assign sc2mac_dat_dst_data114 = sc2mac_dat_data114_d2;
  assign sc2mac_dat_dst_data115 = sc2mac_dat_data115_d2;
  assign sc2mac_dat_dst_data116 = sc2mac_dat_data116_d2;
  assign sc2mac_dat_dst_data117 = sc2mac_dat_data117_d2;
  assign sc2mac_dat_dst_data118 = sc2mac_dat_data118_d2;
  assign sc2mac_dat_dst_data119 = sc2mac_dat_data119_d2;
  assign sc2mac_dat_dst_data12 = sc2mac_dat_data12_d2;
  assign sc2mac_dat_dst_data120 = sc2mac_dat_data120_d2;
  assign sc2mac_dat_dst_data121 = sc2mac_dat_data121_d2;
  assign sc2mac_dat_dst_data122 = sc2mac_dat_data122_d2;
  assign sc2mac_dat_dst_data123 = sc2mac_dat_data123_d2;
  assign sc2mac_dat_dst_data124 = sc2mac_dat_data124_d2;
  assign sc2mac_dat_dst_data125 = sc2mac_dat_data125_d2;
  assign sc2mac_dat_dst_data126 = sc2mac_dat_data126_d2;
  assign sc2mac_dat_dst_data127 = sc2mac_dat_data127_d2;
  assign sc2mac_dat_dst_data13 = sc2mac_dat_data13_d2;
  assign sc2mac_dat_dst_data14 = sc2mac_dat_data14_d2;
  assign sc2mac_dat_dst_data15 = sc2mac_dat_data15_d2;
  assign sc2mac_dat_dst_data16 = sc2mac_dat_data16_d2;
  assign sc2mac_dat_dst_data17 = sc2mac_dat_data17_d2;
  assign sc2mac_dat_dst_data18 = sc2mac_dat_data18_d2;
  assign sc2mac_dat_dst_data19 = sc2mac_dat_data19_d2;
  assign sc2mac_dat_dst_data2 = sc2mac_dat_data2_d2;
  assign sc2mac_dat_dst_data20 = sc2mac_dat_data20_d2;
  assign sc2mac_dat_dst_data21 = sc2mac_dat_data21_d2;
  assign sc2mac_dat_dst_data22 = sc2mac_dat_data22_d2;
  assign sc2mac_dat_dst_data23 = sc2mac_dat_data23_d2;
  assign sc2mac_dat_dst_data24 = sc2mac_dat_data24_d2;
  assign sc2mac_dat_dst_data25 = sc2mac_dat_data25_d2;
  assign sc2mac_dat_dst_data26 = sc2mac_dat_data26_d2;
  assign sc2mac_dat_dst_data27 = sc2mac_dat_data27_d2;
  assign sc2mac_dat_dst_data28 = sc2mac_dat_data28_d2;
  assign sc2mac_dat_dst_data29 = sc2mac_dat_data29_d2;
  assign sc2mac_dat_dst_data3 = sc2mac_dat_data3_d2;
  assign sc2mac_dat_dst_data30 = sc2mac_dat_data30_d2;
  assign sc2mac_dat_dst_data31 = sc2mac_dat_data31_d2;
  assign sc2mac_dat_dst_data32 = sc2mac_dat_data32_d2;
  assign sc2mac_dat_dst_data33 = sc2mac_dat_data33_d2;
  assign sc2mac_dat_dst_data34 = sc2mac_dat_data34_d2;
  assign sc2mac_dat_dst_data35 = sc2mac_dat_data35_d2;
  assign sc2mac_dat_dst_data36 = sc2mac_dat_data36_d2;
  assign sc2mac_dat_dst_data37 = sc2mac_dat_data37_d2;
  assign sc2mac_dat_dst_data38 = sc2mac_dat_data38_d2;
  assign sc2mac_dat_dst_data39 = sc2mac_dat_data39_d2;
  assign sc2mac_dat_dst_data4 = sc2mac_dat_data4_d2;
  assign sc2mac_dat_dst_data40 = sc2mac_dat_data40_d2;
  assign sc2mac_dat_dst_data41 = sc2mac_dat_data41_d2;
  assign sc2mac_dat_dst_data42 = sc2mac_dat_data42_d2;
  assign sc2mac_dat_dst_data43 = sc2mac_dat_data43_d2;
  assign sc2mac_dat_dst_data44 = sc2mac_dat_data44_d2;
  assign sc2mac_dat_dst_data45 = sc2mac_dat_data45_d2;
  assign sc2mac_dat_dst_data46 = sc2mac_dat_data46_d2;
  assign sc2mac_dat_dst_data47 = sc2mac_dat_data47_d2;
  assign sc2mac_dat_dst_data48 = sc2mac_dat_data48_d2;
  assign sc2mac_dat_dst_data49 = sc2mac_dat_data49_d2;
  assign sc2mac_dat_dst_data5 = sc2mac_dat_data5_d2;
  assign sc2mac_dat_dst_data50 = sc2mac_dat_data50_d2;
  assign sc2mac_dat_dst_data51 = sc2mac_dat_data51_d2;
  assign sc2mac_dat_dst_data52 = sc2mac_dat_data52_d2;
  assign sc2mac_dat_dst_data53 = sc2mac_dat_data53_d2;
  assign sc2mac_dat_dst_data54 = sc2mac_dat_data54_d2;
  assign sc2mac_dat_dst_data55 = sc2mac_dat_data55_d2;
  assign sc2mac_dat_dst_data56 = sc2mac_dat_data56_d2;
  assign sc2mac_dat_dst_data57 = sc2mac_dat_data57_d2;
  assign sc2mac_dat_dst_data58 = sc2mac_dat_data58_d2;
  assign sc2mac_dat_dst_data59 = sc2mac_dat_data59_d2;
  assign sc2mac_dat_dst_data6 = sc2mac_dat_data6_d2;
  assign sc2mac_dat_dst_data60 = sc2mac_dat_data60_d2;
  assign sc2mac_dat_dst_data61 = sc2mac_dat_data61_d2;
  assign sc2mac_dat_dst_data62 = sc2mac_dat_data62_d2;
  assign sc2mac_dat_dst_data63 = sc2mac_dat_data63_d2;
  assign sc2mac_dat_dst_data64 = sc2mac_dat_data64_d2;
  assign sc2mac_dat_dst_data65 = sc2mac_dat_data65_d2;
  assign sc2mac_dat_dst_data66 = sc2mac_dat_data66_d2;
  assign sc2mac_dat_dst_data67 = sc2mac_dat_data67_d2;
  assign sc2mac_dat_dst_data68 = sc2mac_dat_data68_d2;
  assign sc2mac_dat_dst_data69 = sc2mac_dat_data69_d2;
  assign sc2mac_dat_dst_data7 = sc2mac_dat_data7_d2;
  assign sc2mac_dat_dst_data70 = sc2mac_dat_data70_d2;
  assign sc2mac_dat_dst_data71 = sc2mac_dat_data71_d2;
  assign sc2mac_dat_dst_data72 = sc2mac_dat_data72_d2;
  assign sc2mac_dat_dst_data73 = sc2mac_dat_data73_d2;
  assign sc2mac_dat_dst_data74 = sc2mac_dat_data74_d2;
  assign sc2mac_dat_dst_data75 = sc2mac_dat_data75_d2;
  assign sc2mac_dat_dst_data76 = sc2mac_dat_data76_d2;
  assign sc2mac_dat_dst_data77 = sc2mac_dat_data77_d2;
  assign sc2mac_dat_dst_data78 = sc2mac_dat_data78_d2;
  assign sc2mac_dat_dst_data79 = sc2mac_dat_data79_d2;
  assign sc2mac_dat_dst_data8 = sc2mac_dat_data8_d2;
  assign sc2mac_dat_dst_data80 = sc2mac_dat_data80_d2;
  assign sc2mac_dat_dst_data81 = sc2mac_dat_data81_d2;
  assign sc2mac_dat_dst_data82 = sc2mac_dat_data82_d2;
  assign sc2mac_dat_dst_data83 = sc2mac_dat_data83_d2;
  assign sc2mac_dat_dst_data84 = sc2mac_dat_data84_d2;
  assign sc2mac_dat_dst_data85 = sc2mac_dat_data85_d2;
  assign sc2mac_dat_dst_data86 = sc2mac_dat_data86_d2;
  assign sc2mac_dat_dst_data87 = sc2mac_dat_data87_d2;
  assign sc2mac_dat_dst_data88 = sc2mac_dat_data88_d2;
  assign sc2mac_dat_dst_data89 = sc2mac_dat_data89_d2;
  assign sc2mac_dat_dst_data9 = sc2mac_dat_data9_d2;
  assign sc2mac_dat_dst_data90 = sc2mac_dat_data90_d2;
  assign sc2mac_dat_dst_data91 = sc2mac_dat_data91_d2;
  assign sc2mac_dat_dst_data92 = sc2mac_dat_data92_d2;
  assign sc2mac_dat_dst_data93 = sc2mac_dat_data93_d2;
  assign sc2mac_dat_dst_data94 = sc2mac_dat_data94_d2;
  assign sc2mac_dat_dst_data95 = sc2mac_dat_data95_d2;
  assign sc2mac_dat_dst_data96 = sc2mac_dat_data96_d2;
  assign sc2mac_dat_dst_data97 = sc2mac_dat_data97_d2;
  assign sc2mac_dat_dst_data98 = sc2mac_dat_data98_d2;
  assign sc2mac_dat_dst_data99 = sc2mac_dat_data99_d2;
  assign sc2mac_dat_dst_mask = sc2mac_dat_mask_d2;
  assign sc2mac_dat_dst_pd = sc2mac_dat_pd_d2;
  assign sc2mac_dat_dst_pvld = sc2mac_dat_pvld_d2;
  assign sc2mac_dat_mask_d0 = sc2mac_dat_src_mask;
  assign sc2mac_dat_pd_d0 = sc2mac_dat_src_pd;
  assign sc2mac_dat_pvld_d0 = sc2mac_dat_src_pvld;
  assign sc2mac_wt_data0_d0 = sc2mac_wt_src_data0;
  assign sc2mac_wt_data100_d0 = sc2mac_wt_src_data100;
  assign sc2mac_wt_data101_d0 = sc2mac_wt_src_data101;
  assign sc2mac_wt_data102_d0 = sc2mac_wt_src_data102;
  assign sc2mac_wt_data103_d0 = sc2mac_wt_src_data103;
  assign sc2mac_wt_data104_d0 = sc2mac_wt_src_data104;
  assign sc2mac_wt_data105_d0 = sc2mac_wt_src_data105;
  assign sc2mac_wt_data106_d0 = sc2mac_wt_src_data106;
  assign sc2mac_wt_data107_d0 = sc2mac_wt_src_data107;
  assign sc2mac_wt_data108_d0 = sc2mac_wt_src_data108;
  assign sc2mac_wt_data109_d0 = sc2mac_wt_src_data109;
  assign sc2mac_wt_data10_d0 = sc2mac_wt_src_data10;
  assign sc2mac_wt_data110_d0 = sc2mac_wt_src_data110;
  assign sc2mac_wt_data111_d0 = sc2mac_wt_src_data111;
  assign sc2mac_wt_data112_d0 = sc2mac_wt_src_data112;
  assign sc2mac_wt_data113_d0 = sc2mac_wt_src_data113;
  assign sc2mac_wt_data114_d0 = sc2mac_wt_src_data114;
  assign sc2mac_wt_data115_d0 = sc2mac_wt_src_data115;
  assign sc2mac_wt_data116_d0 = sc2mac_wt_src_data116;
  assign sc2mac_wt_data117_d0 = sc2mac_wt_src_data117;
  assign sc2mac_wt_data118_d0 = sc2mac_wt_src_data118;
  assign sc2mac_wt_data119_d0 = sc2mac_wt_src_data119;
  assign sc2mac_wt_data11_d0 = sc2mac_wt_src_data11;
  assign sc2mac_wt_data120_d0 = sc2mac_wt_src_data120;
  assign sc2mac_wt_data121_d0 = sc2mac_wt_src_data121;
  assign sc2mac_wt_data122_d0 = sc2mac_wt_src_data122;
  assign sc2mac_wt_data123_d0 = sc2mac_wt_src_data123;
  assign sc2mac_wt_data124_d0 = sc2mac_wt_src_data124;
  assign sc2mac_wt_data125_d0 = sc2mac_wt_src_data125;
  assign sc2mac_wt_data126_d0 = sc2mac_wt_src_data126;
  assign sc2mac_wt_data127_d0 = sc2mac_wt_src_data127;
  assign sc2mac_wt_data12_d0 = sc2mac_wt_src_data12;
  assign sc2mac_wt_data13_d0 = sc2mac_wt_src_data13;
  assign sc2mac_wt_data14_d0 = sc2mac_wt_src_data14;
  assign sc2mac_wt_data15_d0 = sc2mac_wt_src_data15;
  assign sc2mac_wt_data16_d0 = sc2mac_wt_src_data16;
  assign sc2mac_wt_data17_d0 = sc2mac_wt_src_data17;
  assign sc2mac_wt_data18_d0 = sc2mac_wt_src_data18;
  assign sc2mac_wt_data19_d0 = sc2mac_wt_src_data19;
  assign sc2mac_wt_data1_d0 = sc2mac_wt_src_data1;
  assign sc2mac_wt_data20_d0 = sc2mac_wt_src_data20;
  assign sc2mac_wt_data21_d0 = sc2mac_wt_src_data21;
  assign sc2mac_wt_data22_d0 = sc2mac_wt_src_data22;
  assign sc2mac_wt_data23_d0 = sc2mac_wt_src_data23;
  assign sc2mac_wt_data24_d0 = sc2mac_wt_src_data24;
  assign sc2mac_wt_data25_d0 = sc2mac_wt_src_data25;
  assign sc2mac_wt_data26_d0 = sc2mac_wt_src_data26;
  assign sc2mac_wt_data27_d0 = sc2mac_wt_src_data27;
  assign sc2mac_wt_data28_d0 = sc2mac_wt_src_data28;
  assign sc2mac_wt_data29_d0 = sc2mac_wt_src_data29;
  assign sc2mac_wt_data2_d0 = sc2mac_wt_src_data2;
  assign sc2mac_wt_data30_d0 = sc2mac_wt_src_data30;
  assign sc2mac_wt_data31_d0 = sc2mac_wt_src_data31;
  assign sc2mac_wt_data32_d0 = sc2mac_wt_src_data32;
  assign sc2mac_wt_data33_d0 = sc2mac_wt_src_data33;
  assign sc2mac_wt_data34_d0 = sc2mac_wt_src_data34;
  assign sc2mac_wt_data35_d0 = sc2mac_wt_src_data35;
  assign sc2mac_wt_data36_d0 = sc2mac_wt_src_data36;
  assign sc2mac_wt_data37_d0 = sc2mac_wt_src_data37;
  assign sc2mac_wt_data38_d0 = sc2mac_wt_src_data38;
  assign sc2mac_wt_data39_d0 = sc2mac_wt_src_data39;
  assign sc2mac_wt_data3_d0 = sc2mac_wt_src_data3;
  assign sc2mac_wt_data40_d0 = sc2mac_wt_src_data40;
  assign sc2mac_wt_data41_d0 = sc2mac_wt_src_data41;
  assign sc2mac_wt_data42_d0 = sc2mac_wt_src_data42;
  assign sc2mac_wt_data43_d0 = sc2mac_wt_src_data43;
  assign sc2mac_wt_data44_d0 = sc2mac_wt_src_data44;
  assign sc2mac_wt_data45_d0 = sc2mac_wt_src_data45;
  assign sc2mac_wt_data46_d0 = sc2mac_wt_src_data46;
  assign sc2mac_wt_data47_d0 = sc2mac_wt_src_data47;
  assign sc2mac_wt_data48_d0 = sc2mac_wt_src_data48;
  assign sc2mac_wt_data49_d0 = sc2mac_wt_src_data49;
  assign sc2mac_wt_data4_d0 = sc2mac_wt_src_data4;
  assign sc2mac_wt_data50_d0 = sc2mac_wt_src_data50;
  assign sc2mac_wt_data51_d0 = sc2mac_wt_src_data51;
  assign sc2mac_wt_data52_d0 = sc2mac_wt_src_data52;
  assign sc2mac_wt_data53_d0 = sc2mac_wt_src_data53;
  assign sc2mac_wt_data54_d0 = sc2mac_wt_src_data54;
  assign sc2mac_wt_data55_d0 = sc2mac_wt_src_data55;
  assign sc2mac_wt_data56_d0 = sc2mac_wt_src_data56;
  assign sc2mac_wt_data57_d0 = sc2mac_wt_src_data57;
  assign sc2mac_wt_data58_d0 = sc2mac_wt_src_data58;
  assign sc2mac_wt_data59_d0 = sc2mac_wt_src_data59;
  assign sc2mac_wt_data5_d0 = sc2mac_wt_src_data5;
  assign sc2mac_wt_data60_d0 = sc2mac_wt_src_data60;
  assign sc2mac_wt_data61_d0 = sc2mac_wt_src_data61;
  assign sc2mac_wt_data62_d0 = sc2mac_wt_src_data62;
  assign sc2mac_wt_data63_d0 = sc2mac_wt_src_data63;
  assign sc2mac_wt_data64_d0 = sc2mac_wt_src_data64;
  assign sc2mac_wt_data65_d0 = sc2mac_wt_src_data65;
  assign sc2mac_wt_data66_d0 = sc2mac_wt_src_data66;
  assign sc2mac_wt_data67_d0 = sc2mac_wt_src_data67;
  assign sc2mac_wt_data68_d0 = sc2mac_wt_src_data68;
  assign sc2mac_wt_data69_d0 = sc2mac_wt_src_data69;
  assign sc2mac_wt_data6_d0 = sc2mac_wt_src_data6;
  assign sc2mac_wt_data70_d0 = sc2mac_wt_src_data70;
  assign sc2mac_wt_data71_d0 = sc2mac_wt_src_data71;
  assign sc2mac_wt_data72_d0 = sc2mac_wt_src_data72;
  assign sc2mac_wt_data73_d0 = sc2mac_wt_src_data73;
  assign sc2mac_wt_data74_d0 = sc2mac_wt_src_data74;
  assign sc2mac_wt_data75_d0 = sc2mac_wt_src_data75;
  assign sc2mac_wt_data76_d0 = sc2mac_wt_src_data76;
  assign sc2mac_wt_data77_d0 = sc2mac_wt_src_data77;
  assign sc2mac_wt_data78_d0 = sc2mac_wt_src_data78;
  assign sc2mac_wt_data79_d0 = sc2mac_wt_src_data79;
  assign sc2mac_wt_data7_d0 = sc2mac_wt_src_data7;
  assign sc2mac_wt_data80_d0 = sc2mac_wt_src_data80;
  assign sc2mac_wt_data81_d0 = sc2mac_wt_src_data81;
  assign sc2mac_wt_data82_d0 = sc2mac_wt_src_data82;
  assign sc2mac_wt_data83_d0 = sc2mac_wt_src_data83;
  assign sc2mac_wt_data84_d0 = sc2mac_wt_src_data84;
  assign sc2mac_wt_data85_d0 = sc2mac_wt_src_data85;
  assign sc2mac_wt_data86_d0 = sc2mac_wt_src_data86;
  assign sc2mac_wt_data87_d0 = sc2mac_wt_src_data87;
  assign sc2mac_wt_data88_d0 = sc2mac_wt_src_data88;
  assign sc2mac_wt_data89_d0 = sc2mac_wt_src_data89;
  assign sc2mac_wt_data8_d0 = sc2mac_wt_src_data8;
  assign sc2mac_wt_data90_d0 = sc2mac_wt_src_data90;
  assign sc2mac_wt_data91_d0 = sc2mac_wt_src_data91;
  assign sc2mac_wt_data92_d0 = sc2mac_wt_src_data92;
  assign sc2mac_wt_data93_d0 = sc2mac_wt_src_data93;
  assign sc2mac_wt_data94_d0 = sc2mac_wt_src_data94;
  assign sc2mac_wt_data95_d0 = sc2mac_wt_src_data95;
  assign sc2mac_wt_data96_d0 = sc2mac_wt_src_data96;
  assign sc2mac_wt_data97_d0 = sc2mac_wt_src_data97;
  assign sc2mac_wt_data98_d0 = sc2mac_wt_src_data98;
  assign sc2mac_wt_data99_d0 = sc2mac_wt_src_data99;
  assign sc2mac_wt_data9_d0 = sc2mac_wt_src_data9;
  assign sc2mac_wt_dst_data0 = sc2mac_wt_data0_d2;
  assign sc2mac_wt_dst_data1 = sc2mac_wt_data1_d2;
  assign sc2mac_wt_dst_data10 = sc2mac_wt_data10_d2;
  assign sc2mac_wt_dst_data100 = sc2mac_wt_data100_d2;
  assign sc2mac_wt_dst_data101 = sc2mac_wt_data101_d2;
  assign sc2mac_wt_dst_data102 = sc2mac_wt_data102_d2;
  assign sc2mac_wt_dst_data103 = sc2mac_wt_data103_d2;
  assign sc2mac_wt_dst_data104 = sc2mac_wt_data104_d2;
  assign sc2mac_wt_dst_data105 = sc2mac_wt_data105_d2;
  assign sc2mac_wt_dst_data106 = sc2mac_wt_data106_d2;
  assign sc2mac_wt_dst_data107 = sc2mac_wt_data107_d2;
  assign sc2mac_wt_dst_data108 = sc2mac_wt_data108_d2;
  assign sc2mac_wt_dst_data109 = sc2mac_wt_data109_d2;
  assign sc2mac_wt_dst_data11 = sc2mac_wt_data11_d2;
  assign sc2mac_wt_dst_data110 = sc2mac_wt_data110_d2;
  assign sc2mac_wt_dst_data111 = sc2mac_wt_data111_d2;
  assign sc2mac_wt_dst_data112 = sc2mac_wt_data112_d2;
  assign sc2mac_wt_dst_data113 = sc2mac_wt_data113_d2;
  assign sc2mac_wt_dst_data114 = sc2mac_wt_data114_d2;
  assign sc2mac_wt_dst_data115 = sc2mac_wt_data115_d2;
  assign sc2mac_wt_dst_data116 = sc2mac_wt_data116_d2;
  assign sc2mac_wt_dst_data117 = sc2mac_wt_data117_d2;
  assign sc2mac_wt_dst_data118 = sc2mac_wt_data118_d2;
  assign sc2mac_wt_dst_data119 = sc2mac_wt_data119_d2;
  assign sc2mac_wt_dst_data12 = sc2mac_wt_data12_d2;
  assign sc2mac_wt_dst_data120 = sc2mac_wt_data120_d2;
  assign sc2mac_wt_dst_data121 = sc2mac_wt_data121_d2;
  assign sc2mac_wt_dst_data122 = sc2mac_wt_data122_d2;
  assign sc2mac_wt_dst_data123 = sc2mac_wt_data123_d2;
  assign sc2mac_wt_dst_data124 = sc2mac_wt_data124_d2;
  assign sc2mac_wt_dst_data125 = sc2mac_wt_data125_d2;
  assign sc2mac_wt_dst_data126 = sc2mac_wt_data126_d2;
  assign sc2mac_wt_dst_data127 = sc2mac_wt_data127_d2;
  assign sc2mac_wt_dst_data13 = sc2mac_wt_data13_d2;
  assign sc2mac_wt_dst_data14 = sc2mac_wt_data14_d2;
  assign sc2mac_wt_dst_data15 = sc2mac_wt_data15_d2;
  assign sc2mac_wt_dst_data16 = sc2mac_wt_data16_d2;
  assign sc2mac_wt_dst_data17 = sc2mac_wt_data17_d2;
  assign sc2mac_wt_dst_data18 = sc2mac_wt_data18_d2;
  assign sc2mac_wt_dst_data19 = sc2mac_wt_data19_d2;
  assign sc2mac_wt_dst_data2 = sc2mac_wt_data2_d2;
  assign sc2mac_wt_dst_data20 = sc2mac_wt_data20_d2;
  assign sc2mac_wt_dst_data21 = sc2mac_wt_data21_d2;
  assign sc2mac_wt_dst_data22 = sc2mac_wt_data22_d2;
  assign sc2mac_wt_dst_data23 = sc2mac_wt_data23_d2;
  assign sc2mac_wt_dst_data24 = sc2mac_wt_data24_d2;
  assign sc2mac_wt_dst_data25 = sc2mac_wt_data25_d2;
  assign sc2mac_wt_dst_data26 = sc2mac_wt_data26_d2;
  assign sc2mac_wt_dst_data27 = sc2mac_wt_data27_d2;
  assign sc2mac_wt_dst_data28 = sc2mac_wt_data28_d2;
  assign sc2mac_wt_dst_data29 = sc2mac_wt_data29_d2;
  assign sc2mac_wt_dst_data3 = sc2mac_wt_data3_d2;
  assign sc2mac_wt_dst_data30 = sc2mac_wt_data30_d2;
  assign sc2mac_wt_dst_data31 = sc2mac_wt_data31_d2;
  assign sc2mac_wt_dst_data32 = sc2mac_wt_data32_d2;
  assign sc2mac_wt_dst_data33 = sc2mac_wt_data33_d2;
  assign sc2mac_wt_dst_data34 = sc2mac_wt_data34_d2;
  assign sc2mac_wt_dst_data35 = sc2mac_wt_data35_d2;
  assign sc2mac_wt_dst_data36 = sc2mac_wt_data36_d2;
  assign sc2mac_wt_dst_data37 = sc2mac_wt_data37_d2;
  assign sc2mac_wt_dst_data38 = sc2mac_wt_data38_d2;
  assign sc2mac_wt_dst_data39 = sc2mac_wt_data39_d2;
  assign sc2mac_wt_dst_data4 = sc2mac_wt_data4_d2;
  assign sc2mac_wt_dst_data40 = sc2mac_wt_data40_d2;
  assign sc2mac_wt_dst_data41 = sc2mac_wt_data41_d2;
  assign sc2mac_wt_dst_data42 = sc2mac_wt_data42_d2;
  assign sc2mac_wt_dst_data43 = sc2mac_wt_data43_d2;
  assign sc2mac_wt_dst_data44 = sc2mac_wt_data44_d2;
  assign sc2mac_wt_dst_data45 = sc2mac_wt_data45_d2;
  assign sc2mac_wt_dst_data46 = sc2mac_wt_data46_d2;
  assign sc2mac_wt_dst_data47 = sc2mac_wt_data47_d2;
  assign sc2mac_wt_dst_data48 = sc2mac_wt_data48_d2;
  assign sc2mac_wt_dst_data49 = sc2mac_wt_data49_d2;
  assign sc2mac_wt_dst_data5 = sc2mac_wt_data5_d2;
  assign sc2mac_wt_dst_data50 = sc2mac_wt_data50_d2;
  assign sc2mac_wt_dst_data51 = sc2mac_wt_data51_d2;
  assign sc2mac_wt_dst_data52 = sc2mac_wt_data52_d2;
  assign sc2mac_wt_dst_data53 = sc2mac_wt_data53_d2;
  assign sc2mac_wt_dst_data54 = sc2mac_wt_data54_d2;
  assign sc2mac_wt_dst_data55 = sc2mac_wt_data55_d2;
  assign sc2mac_wt_dst_data56 = sc2mac_wt_data56_d2;
  assign sc2mac_wt_dst_data57 = sc2mac_wt_data57_d2;
  assign sc2mac_wt_dst_data58 = sc2mac_wt_data58_d2;
  assign sc2mac_wt_dst_data59 = sc2mac_wt_data59_d2;
  assign sc2mac_wt_dst_data6 = sc2mac_wt_data6_d2;
  assign sc2mac_wt_dst_data60 = sc2mac_wt_data60_d2;
  assign sc2mac_wt_dst_data61 = sc2mac_wt_data61_d2;
  assign sc2mac_wt_dst_data62 = sc2mac_wt_data62_d2;
  assign sc2mac_wt_dst_data63 = sc2mac_wt_data63_d2;
  assign sc2mac_wt_dst_data64 = sc2mac_wt_data64_d2;
  assign sc2mac_wt_dst_data65 = sc2mac_wt_data65_d2;
  assign sc2mac_wt_dst_data66 = sc2mac_wt_data66_d2;
  assign sc2mac_wt_dst_data67 = sc2mac_wt_data67_d2;
  assign sc2mac_wt_dst_data68 = sc2mac_wt_data68_d2;
  assign sc2mac_wt_dst_data69 = sc2mac_wt_data69_d2;
  assign sc2mac_wt_dst_data7 = sc2mac_wt_data7_d2;
  assign sc2mac_wt_dst_data70 = sc2mac_wt_data70_d2;
  assign sc2mac_wt_dst_data71 = sc2mac_wt_data71_d2;
  assign sc2mac_wt_dst_data72 = sc2mac_wt_data72_d2;
  assign sc2mac_wt_dst_data73 = sc2mac_wt_data73_d2;
  assign sc2mac_wt_dst_data74 = sc2mac_wt_data74_d2;
  assign sc2mac_wt_dst_data75 = sc2mac_wt_data75_d2;
  assign sc2mac_wt_dst_data76 = sc2mac_wt_data76_d2;
  assign sc2mac_wt_dst_data77 = sc2mac_wt_data77_d2;
  assign sc2mac_wt_dst_data78 = sc2mac_wt_data78_d2;
  assign sc2mac_wt_dst_data79 = sc2mac_wt_data79_d2;
  assign sc2mac_wt_dst_data8 = sc2mac_wt_data8_d2;
  assign sc2mac_wt_dst_data80 = sc2mac_wt_data80_d2;
  assign sc2mac_wt_dst_data81 = sc2mac_wt_data81_d2;
  assign sc2mac_wt_dst_data82 = sc2mac_wt_data82_d2;
  assign sc2mac_wt_dst_data83 = sc2mac_wt_data83_d2;
  assign sc2mac_wt_dst_data84 = sc2mac_wt_data84_d2;
  assign sc2mac_wt_dst_data85 = sc2mac_wt_data85_d2;
  assign sc2mac_wt_dst_data86 = sc2mac_wt_data86_d2;
  assign sc2mac_wt_dst_data87 = sc2mac_wt_data87_d2;
  assign sc2mac_wt_dst_data88 = sc2mac_wt_data88_d2;
  assign sc2mac_wt_dst_data89 = sc2mac_wt_data89_d2;
  assign sc2mac_wt_dst_data9 = sc2mac_wt_data9_d2;
  assign sc2mac_wt_dst_data90 = sc2mac_wt_data90_d2;
  assign sc2mac_wt_dst_data91 = sc2mac_wt_data91_d2;
  assign sc2mac_wt_dst_data92 = sc2mac_wt_data92_d2;
  assign sc2mac_wt_dst_data93 = sc2mac_wt_data93_d2;
  assign sc2mac_wt_dst_data94 = sc2mac_wt_data94_d2;
  assign sc2mac_wt_dst_data95 = sc2mac_wt_data95_d2;
  assign sc2mac_wt_dst_data96 = sc2mac_wt_data96_d2;
  assign sc2mac_wt_dst_data97 = sc2mac_wt_data97_d2;
  assign sc2mac_wt_dst_data98 = sc2mac_wt_data98_d2;
  assign sc2mac_wt_dst_data99 = sc2mac_wt_data99_d2;
  assign sc2mac_wt_dst_mask = sc2mac_wt_mask_d2;
  assign sc2mac_wt_dst_pvld = sc2mac_wt_pvld_d2;
  assign sc2mac_wt_dst_sel = sc2mac_wt_sel_d2;
  assign sc2mac_wt_mask_d0 = sc2mac_wt_src_mask;
  assign sc2mac_wt_pvld_d0 = sc2mac_wt_src_pvld;
  assign sc2mac_wt_sel_d0 = sc2mac_wt_src_sel;
endmodule
