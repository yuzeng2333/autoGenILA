module FP17_MUL_chn_a_rsci_unreg(in_0, outsig);
  (* src = "./vmod/vlibs/HLS_fp17_mul.v:96" *)
  input in_0;
  (* src = "./vmod/vlibs/HLS_fp17_mul.v:97" *)
  output outsig;
  assign outsig = in_0;
endmodule
